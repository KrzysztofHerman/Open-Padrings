magic
tech ihp-sg13g2
magscale 1 2
timestamp 1757428966
<< metal1 >>
rect 71616 151976 152352 152000
rect 71616 151936 75392 151976
rect 75432 151936 75474 151976
rect 75514 151936 75556 151976
rect 75596 151936 75638 151976
rect 75678 151936 75720 151976
rect 75760 151936 90512 151976
rect 90552 151936 90594 151976
rect 90634 151936 90676 151976
rect 90716 151936 90758 151976
rect 90798 151936 90840 151976
rect 90880 151936 105632 151976
rect 105672 151936 105714 151976
rect 105754 151936 105796 151976
rect 105836 151936 105878 151976
rect 105918 151936 105960 151976
rect 106000 151936 120752 151976
rect 120792 151936 120834 151976
rect 120874 151936 120916 151976
rect 120956 151936 120998 151976
rect 121038 151936 121080 151976
rect 121120 151936 135872 151976
rect 135912 151936 135954 151976
rect 135994 151936 136036 151976
rect 136076 151936 136118 151976
rect 136158 151936 136200 151976
rect 136240 151936 150992 151976
rect 151032 151936 151074 151976
rect 151114 151936 151156 151976
rect 151196 151936 151238 151976
rect 151278 151936 151320 151976
rect 151360 151936 152352 151976
rect 71616 151912 152352 151936
rect 71616 151220 152352 151244
rect 71616 151180 74152 151220
rect 74192 151180 74234 151220
rect 74274 151180 74316 151220
rect 74356 151180 74398 151220
rect 74438 151180 74480 151220
rect 74520 151180 89272 151220
rect 89312 151180 89354 151220
rect 89394 151180 89436 151220
rect 89476 151180 89518 151220
rect 89558 151180 89600 151220
rect 89640 151180 104392 151220
rect 104432 151180 104474 151220
rect 104514 151180 104556 151220
rect 104596 151180 104638 151220
rect 104678 151180 104720 151220
rect 104760 151180 119512 151220
rect 119552 151180 119594 151220
rect 119634 151180 119676 151220
rect 119716 151180 119758 151220
rect 119798 151180 119840 151220
rect 119880 151180 134632 151220
rect 134672 151180 134714 151220
rect 134754 151180 134796 151220
rect 134836 151180 134878 151220
rect 134918 151180 134960 151220
rect 135000 151180 149752 151220
rect 149792 151180 149834 151220
rect 149874 151180 149916 151220
rect 149956 151180 149998 151220
rect 150038 151180 150080 151220
rect 150120 151180 152352 151220
rect 71616 151156 152352 151180
rect 71616 150464 152352 150488
rect 71616 150424 75392 150464
rect 75432 150424 75474 150464
rect 75514 150424 75556 150464
rect 75596 150424 75638 150464
rect 75678 150424 75720 150464
rect 75760 150424 90512 150464
rect 90552 150424 90594 150464
rect 90634 150424 90676 150464
rect 90716 150424 90758 150464
rect 90798 150424 90840 150464
rect 90880 150424 105632 150464
rect 105672 150424 105714 150464
rect 105754 150424 105796 150464
rect 105836 150424 105878 150464
rect 105918 150424 105960 150464
rect 106000 150424 120752 150464
rect 120792 150424 120834 150464
rect 120874 150424 120916 150464
rect 120956 150424 120998 150464
rect 121038 150424 121080 150464
rect 121120 150424 135872 150464
rect 135912 150424 135954 150464
rect 135994 150424 136036 150464
rect 136076 150424 136118 150464
rect 136158 150424 136200 150464
rect 136240 150424 150992 150464
rect 151032 150424 151074 150464
rect 151114 150424 151156 150464
rect 151196 150424 151238 150464
rect 151278 150424 151320 150464
rect 151360 150424 152352 150464
rect 71616 150400 152352 150424
rect 71616 149708 152352 149732
rect 71616 149668 74152 149708
rect 74192 149668 74234 149708
rect 74274 149668 74316 149708
rect 74356 149668 74398 149708
rect 74438 149668 74480 149708
rect 74520 149668 89272 149708
rect 89312 149668 89354 149708
rect 89394 149668 89436 149708
rect 89476 149668 89518 149708
rect 89558 149668 89600 149708
rect 89640 149668 104392 149708
rect 104432 149668 104474 149708
rect 104514 149668 104556 149708
rect 104596 149668 104638 149708
rect 104678 149668 104720 149708
rect 104760 149668 119512 149708
rect 119552 149668 119594 149708
rect 119634 149668 119676 149708
rect 119716 149668 119758 149708
rect 119798 149668 119840 149708
rect 119880 149668 134632 149708
rect 134672 149668 134714 149708
rect 134754 149668 134796 149708
rect 134836 149668 134878 149708
rect 134918 149668 134960 149708
rect 135000 149668 149752 149708
rect 149792 149668 149834 149708
rect 149874 149668 149916 149708
rect 149956 149668 149998 149708
rect 150038 149668 150080 149708
rect 150120 149668 152352 149708
rect 71616 149644 152352 149668
rect 71616 148952 152352 148976
rect 71616 148912 75392 148952
rect 75432 148912 75474 148952
rect 75514 148912 75556 148952
rect 75596 148912 75638 148952
rect 75678 148912 75720 148952
rect 75760 148912 90512 148952
rect 90552 148912 90594 148952
rect 90634 148912 90676 148952
rect 90716 148912 90758 148952
rect 90798 148912 90840 148952
rect 90880 148912 105632 148952
rect 105672 148912 105714 148952
rect 105754 148912 105796 148952
rect 105836 148912 105878 148952
rect 105918 148912 105960 148952
rect 106000 148912 120752 148952
rect 120792 148912 120834 148952
rect 120874 148912 120916 148952
rect 120956 148912 120998 148952
rect 121038 148912 121080 148952
rect 121120 148912 135872 148952
rect 135912 148912 135954 148952
rect 135994 148912 136036 148952
rect 136076 148912 136118 148952
rect 136158 148912 136200 148952
rect 136240 148912 150992 148952
rect 151032 148912 151074 148952
rect 151114 148912 151156 148952
rect 151196 148912 151238 148952
rect 151278 148912 151320 148952
rect 151360 148912 152352 148952
rect 71616 148888 152352 148912
rect 71616 148196 152352 148220
rect 71616 148156 74152 148196
rect 74192 148156 74234 148196
rect 74274 148156 74316 148196
rect 74356 148156 74398 148196
rect 74438 148156 74480 148196
rect 74520 148156 89272 148196
rect 89312 148156 89354 148196
rect 89394 148156 89436 148196
rect 89476 148156 89518 148196
rect 89558 148156 89600 148196
rect 89640 148156 104392 148196
rect 104432 148156 104474 148196
rect 104514 148156 104556 148196
rect 104596 148156 104638 148196
rect 104678 148156 104720 148196
rect 104760 148156 119512 148196
rect 119552 148156 119594 148196
rect 119634 148156 119676 148196
rect 119716 148156 119758 148196
rect 119798 148156 119840 148196
rect 119880 148156 134632 148196
rect 134672 148156 134714 148196
rect 134754 148156 134796 148196
rect 134836 148156 134878 148196
rect 134918 148156 134960 148196
rect 135000 148156 149752 148196
rect 149792 148156 149834 148196
rect 149874 148156 149916 148196
rect 149956 148156 149998 148196
rect 150038 148156 150080 148196
rect 150120 148156 152352 148196
rect 71616 148132 152352 148156
rect 71616 147440 152352 147464
rect 71616 147400 75392 147440
rect 75432 147400 75474 147440
rect 75514 147400 75556 147440
rect 75596 147400 75638 147440
rect 75678 147400 75720 147440
rect 75760 147400 90512 147440
rect 90552 147400 90594 147440
rect 90634 147400 90676 147440
rect 90716 147400 90758 147440
rect 90798 147400 90840 147440
rect 90880 147400 105632 147440
rect 105672 147400 105714 147440
rect 105754 147400 105796 147440
rect 105836 147400 105878 147440
rect 105918 147400 105960 147440
rect 106000 147400 120752 147440
rect 120792 147400 120834 147440
rect 120874 147400 120916 147440
rect 120956 147400 120998 147440
rect 121038 147400 121080 147440
rect 121120 147400 135872 147440
rect 135912 147400 135954 147440
rect 135994 147400 136036 147440
rect 136076 147400 136118 147440
rect 136158 147400 136200 147440
rect 136240 147400 150992 147440
rect 151032 147400 151074 147440
rect 151114 147400 151156 147440
rect 151196 147400 151238 147440
rect 151278 147400 151320 147440
rect 151360 147400 152352 147440
rect 71616 147376 152352 147400
rect 71616 146684 152352 146708
rect 71616 146644 74152 146684
rect 74192 146644 74234 146684
rect 74274 146644 74316 146684
rect 74356 146644 74398 146684
rect 74438 146644 74480 146684
rect 74520 146644 89272 146684
rect 89312 146644 89354 146684
rect 89394 146644 89436 146684
rect 89476 146644 89518 146684
rect 89558 146644 89600 146684
rect 89640 146644 104392 146684
rect 104432 146644 104474 146684
rect 104514 146644 104556 146684
rect 104596 146644 104638 146684
rect 104678 146644 104720 146684
rect 104760 146644 119512 146684
rect 119552 146644 119594 146684
rect 119634 146644 119676 146684
rect 119716 146644 119758 146684
rect 119798 146644 119840 146684
rect 119880 146644 134632 146684
rect 134672 146644 134714 146684
rect 134754 146644 134796 146684
rect 134836 146644 134878 146684
rect 134918 146644 134960 146684
rect 135000 146644 149752 146684
rect 149792 146644 149834 146684
rect 149874 146644 149916 146684
rect 149956 146644 149998 146684
rect 150038 146644 150080 146684
rect 150120 146644 152352 146684
rect 71616 146620 152352 146644
rect 71616 145928 152352 145952
rect 71616 145888 75392 145928
rect 75432 145888 75474 145928
rect 75514 145888 75556 145928
rect 75596 145888 75638 145928
rect 75678 145888 75720 145928
rect 75760 145888 90512 145928
rect 90552 145888 90594 145928
rect 90634 145888 90676 145928
rect 90716 145888 90758 145928
rect 90798 145888 90840 145928
rect 90880 145888 105632 145928
rect 105672 145888 105714 145928
rect 105754 145888 105796 145928
rect 105836 145888 105878 145928
rect 105918 145888 105960 145928
rect 106000 145888 120752 145928
rect 120792 145888 120834 145928
rect 120874 145888 120916 145928
rect 120956 145888 120998 145928
rect 121038 145888 121080 145928
rect 121120 145888 135872 145928
rect 135912 145888 135954 145928
rect 135994 145888 136036 145928
rect 136076 145888 136118 145928
rect 136158 145888 136200 145928
rect 136240 145888 150992 145928
rect 151032 145888 151074 145928
rect 151114 145888 151156 145928
rect 151196 145888 151238 145928
rect 151278 145888 151320 145928
rect 151360 145888 152352 145928
rect 71616 145864 152352 145888
rect 71616 145172 152352 145196
rect 71616 145132 74152 145172
rect 74192 145132 74234 145172
rect 74274 145132 74316 145172
rect 74356 145132 74398 145172
rect 74438 145132 74480 145172
rect 74520 145132 89272 145172
rect 89312 145132 89354 145172
rect 89394 145132 89436 145172
rect 89476 145132 89518 145172
rect 89558 145132 89600 145172
rect 89640 145132 104392 145172
rect 104432 145132 104474 145172
rect 104514 145132 104556 145172
rect 104596 145132 104638 145172
rect 104678 145132 104720 145172
rect 104760 145132 119512 145172
rect 119552 145132 119594 145172
rect 119634 145132 119676 145172
rect 119716 145132 119758 145172
rect 119798 145132 119840 145172
rect 119880 145132 134632 145172
rect 134672 145132 134714 145172
rect 134754 145132 134796 145172
rect 134836 145132 134878 145172
rect 134918 145132 134960 145172
rect 135000 145132 149752 145172
rect 149792 145132 149834 145172
rect 149874 145132 149916 145172
rect 149956 145132 149998 145172
rect 150038 145132 150080 145172
rect 150120 145132 152352 145172
rect 71616 145108 152352 145132
rect 71616 144416 152352 144440
rect 71616 144376 75392 144416
rect 75432 144376 75474 144416
rect 75514 144376 75556 144416
rect 75596 144376 75638 144416
rect 75678 144376 75720 144416
rect 75760 144376 90512 144416
rect 90552 144376 90594 144416
rect 90634 144376 90676 144416
rect 90716 144376 90758 144416
rect 90798 144376 90840 144416
rect 90880 144376 105632 144416
rect 105672 144376 105714 144416
rect 105754 144376 105796 144416
rect 105836 144376 105878 144416
rect 105918 144376 105960 144416
rect 106000 144376 120752 144416
rect 120792 144376 120834 144416
rect 120874 144376 120916 144416
rect 120956 144376 120998 144416
rect 121038 144376 121080 144416
rect 121120 144376 135872 144416
rect 135912 144376 135954 144416
rect 135994 144376 136036 144416
rect 136076 144376 136118 144416
rect 136158 144376 136200 144416
rect 136240 144376 150992 144416
rect 151032 144376 151074 144416
rect 151114 144376 151156 144416
rect 151196 144376 151238 144416
rect 151278 144376 151320 144416
rect 151360 144376 152352 144416
rect 71616 144352 152352 144376
rect 71616 143660 152352 143684
rect 71616 143620 74152 143660
rect 74192 143620 74234 143660
rect 74274 143620 74316 143660
rect 74356 143620 74398 143660
rect 74438 143620 74480 143660
rect 74520 143620 89272 143660
rect 89312 143620 89354 143660
rect 89394 143620 89436 143660
rect 89476 143620 89518 143660
rect 89558 143620 89600 143660
rect 89640 143620 104392 143660
rect 104432 143620 104474 143660
rect 104514 143620 104556 143660
rect 104596 143620 104638 143660
rect 104678 143620 104720 143660
rect 104760 143620 119512 143660
rect 119552 143620 119594 143660
rect 119634 143620 119676 143660
rect 119716 143620 119758 143660
rect 119798 143620 119840 143660
rect 119880 143620 134632 143660
rect 134672 143620 134714 143660
rect 134754 143620 134796 143660
rect 134836 143620 134878 143660
rect 134918 143620 134960 143660
rect 135000 143620 149752 143660
rect 149792 143620 149834 143660
rect 149874 143620 149916 143660
rect 149956 143620 149998 143660
rect 150038 143620 150080 143660
rect 150120 143620 152352 143660
rect 71616 143596 152352 143620
rect 71616 142904 152352 142928
rect 71616 142864 75392 142904
rect 75432 142864 75474 142904
rect 75514 142864 75556 142904
rect 75596 142864 75638 142904
rect 75678 142864 75720 142904
rect 75760 142864 90512 142904
rect 90552 142864 90594 142904
rect 90634 142864 90676 142904
rect 90716 142864 90758 142904
rect 90798 142864 90840 142904
rect 90880 142864 105632 142904
rect 105672 142864 105714 142904
rect 105754 142864 105796 142904
rect 105836 142864 105878 142904
rect 105918 142864 105960 142904
rect 106000 142864 120752 142904
rect 120792 142864 120834 142904
rect 120874 142864 120916 142904
rect 120956 142864 120998 142904
rect 121038 142864 121080 142904
rect 121120 142864 135872 142904
rect 135912 142864 135954 142904
rect 135994 142864 136036 142904
rect 136076 142864 136118 142904
rect 136158 142864 136200 142904
rect 136240 142864 150992 142904
rect 151032 142864 151074 142904
rect 151114 142864 151156 142904
rect 151196 142864 151238 142904
rect 151278 142864 151320 142904
rect 151360 142864 152352 142904
rect 71616 142840 152352 142864
rect 71616 142148 152352 142172
rect 71616 142108 74152 142148
rect 74192 142108 74234 142148
rect 74274 142108 74316 142148
rect 74356 142108 74398 142148
rect 74438 142108 74480 142148
rect 74520 142108 89272 142148
rect 89312 142108 89354 142148
rect 89394 142108 89436 142148
rect 89476 142108 89518 142148
rect 89558 142108 89600 142148
rect 89640 142108 104392 142148
rect 104432 142108 104474 142148
rect 104514 142108 104556 142148
rect 104596 142108 104638 142148
rect 104678 142108 104720 142148
rect 104760 142108 119512 142148
rect 119552 142108 119594 142148
rect 119634 142108 119676 142148
rect 119716 142108 119758 142148
rect 119798 142108 119840 142148
rect 119880 142108 134632 142148
rect 134672 142108 134714 142148
rect 134754 142108 134796 142148
rect 134836 142108 134878 142148
rect 134918 142108 134960 142148
rect 135000 142108 149752 142148
rect 149792 142108 149834 142148
rect 149874 142108 149916 142148
rect 149956 142108 149998 142148
rect 150038 142108 150080 142148
rect 150120 142108 152352 142148
rect 71616 142084 152352 142108
rect 71616 141392 152352 141416
rect 71616 141352 75392 141392
rect 75432 141352 75474 141392
rect 75514 141352 75556 141392
rect 75596 141352 75638 141392
rect 75678 141352 75720 141392
rect 75760 141352 90512 141392
rect 90552 141352 90594 141392
rect 90634 141352 90676 141392
rect 90716 141352 90758 141392
rect 90798 141352 90840 141392
rect 90880 141352 105632 141392
rect 105672 141352 105714 141392
rect 105754 141352 105796 141392
rect 105836 141352 105878 141392
rect 105918 141352 105960 141392
rect 106000 141352 120752 141392
rect 120792 141352 120834 141392
rect 120874 141352 120916 141392
rect 120956 141352 120998 141392
rect 121038 141352 121080 141392
rect 121120 141352 135872 141392
rect 135912 141352 135954 141392
rect 135994 141352 136036 141392
rect 136076 141352 136118 141392
rect 136158 141352 136200 141392
rect 136240 141352 150992 141392
rect 151032 141352 151074 141392
rect 151114 141352 151156 141392
rect 151196 141352 151238 141392
rect 151278 141352 151320 141392
rect 151360 141352 152352 141392
rect 71616 141328 152352 141352
rect 71616 140636 152352 140660
rect 71616 140596 74152 140636
rect 74192 140596 74234 140636
rect 74274 140596 74316 140636
rect 74356 140596 74398 140636
rect 74438 140596 74480 140636
rect 74520 140596 89272 140636
rect 89312 140596 89354 140636
rect 89394 140596 89436 140636
rect 89476 140596 89518 140636
rect 89558 140596 89600 140636
rect 89640 140596 104392 140636
rect 104432 140596 104474 140636
rect 104514 140596 104556 140636
rect 104596 140596 104638 140636
rect 104678 140596 104720 140636
rect 104760 140596 119512 140636
rect 119552 140596 119594 140636
rect 119634 140596 119676 140636
rect 119716 140596 119758 140636
rect 119798 140596 119840 140636
rect 119880 140596 134632 140636
rect 134672 140596 134714 140636
rect 134754 140596 134796 140636
rect 134836 140596 134878 140636
rect 134918 140596 134960 140636
rect 135000 140596 149752 140636
rect 149792 140596 149834 140636
rect 149874 140596 149916 140636
rect 149956 140596 149998 140636
rect 150038 140596 150080 140636
rect 150120 140596 152352 140636
rect 71616 140572 152352 140596
rect 71616 139880 152352 139904
rect 71616 139840 75392 139880
rect 75432 139840 75474 139880
rect 75514 139840 75556 139880
rect 75596 139840 75638 139880
rect 75678 139840 75720 139880
rect 75760 139840 90512 139880
rect 90552 139840 90594 139880
rect 90634 139840 90676 139880
rect 90716 139840 90758 139880
rect 90798 139840 90840 139880
rect 90880 139840 105632 139880
rect 105672 139840 105714 139880
rect 105754 139840 105796 139880
rect 105836 139840 105878 139880
rect 105918 139840 105960 139880
rect 106000 139840 120752 139880
rect 120792 139840 120834 139880
rect 120874 139840 120916 139880
rect 120956 139840 120998 139880
rect 121038 139840 121080 139880
rect 121120 139840 135872 139880
rect 135912 139840 135954 139880
rect 135994 139840 136036 139880
rect 136076 139840 136118 139880
rect 136158 139840 136200 139880
rect 136240 139840 150992 139880
rect 151032 139840 151074 139880
rect 151114 139840 151156 139880
rect 151196 139840 151238 139880
rect 151278 139840 151320 139880
rect 151360 139840 152352 139880
rect 71616 139816 152352 139840
rect 71616 139124 152352 139148
rect 71616 139084 74152 139124
rect 74192 139084 74234 139124
rect 74274 139084 74316 139124
rect 74356 139084 74398 139124
rect 74438 139084 74480 139124
rect 74520 139084 89272 139124
rect 89312 139084 89354 139124
rect 89394 139084 89436 139124
rect 89476 139084 89518 139124
rect 89558 139084 89600 139124
rect 89640 139084 104392 139124
rect 104432 139084 104474 139124
rect 104514 139084 104556 139124
rect 104596 139084 104638 139124
rect 104678 139084 104720 139124
rect 104760 139084 119512 139124
rect 119552 139084 119594 139124
rect 119634 139084 119676 139124
rect 119716 139084 119758 139124
rect 119798 139084 119840 139124
rect 119880 139084 134632 139124
rect 134672 139084 134714 139124
rect 134754 139084 134796 139124
rect 134836 139084 134878 139124
rect 134918 139084 134960 139124
rect 135000 139084 149752 139124
rect 149792 139084 149834 139124
rect 149874 139084 149916 139124
rect 149956 139084 149998 139124
rect 150038 139084 150080 139124
rect 150120 139084 152352 139124
rect 71616 139060 152352 139084
rect 71616 138368 152352 138392
rect 71616 138328 75392 138368
rect 75432 138328 75474 138368
rect 75514 138328 75556 138368
rect 75596 138328 75638 138368
rect 75678 138328 75720 138368
rect 75760 138328 90512 138368
rect 90552 138328 90594 138368
rect 90634 138328 90676 138368
rect 90716 138328 90758 138368
rect 90798 138328 90840 138368
rect 90880 138328 105632 138368
rect 105672 138328 105714 138368
rect 105754 138328 105796 138368
rect 105836 138328 105878 138368
rect 105918 138328 105960 138368
rect 106000 138328 120752 138368
rect 120792 138328 120834 138368
rect 120874 138328 120916 138368
rect 120956 138328 120998 138368
rect 121038 138328 121080 138368
rect 121120 138328 135872 138368
rect 135912 138328 135954 138368
rect 135994 138328 136036 138368
rect 136076 138328 136118 138368
rect 136158 138328 136200 138368
rect 136240 138328 150992 138368
rect 151032 138328 151074 138368
rect 151114 138328 151156 138368
rect 151196 138328 151238 138368
rect 151278 138328 151320 138368
rect 151360 138328 152352 138368
rect 71616 138304 152352 138328
rect 71616 137612 152352 137636
rect 71616 137572 74152 137612
rect 74192 137572 74234 137612
rect 74274 137572 74316 137612
rect 74356 137572 74398 137612
rect 74438 137572 74480 137612
rect 74520 137572 89272 137612
rect 89312 137572 89354 137612
rect 89394 137572 89436 137612
rect 89476 137572 89518 137612
rect 89558 137572 89600 137612
rect 89640 137572 104392 137612
rect 104432 137572 104474 137612
rect 104514 137572 104556 137612
rect 104596 137572 104638 137612
rect 104678 137572 104720 137612
rect 104760 137572 119512 137612
rect 119552 137572 119594 137612
rect 119634 137572 119676 137612
rect 119716 137572 119758 137612
rect 119798 137572 119840 137612
rect 119880 137572 134632 137612
rect 134672 137572 134714 137612
rect 134754 137572 134796 137612
rect 134836 137572 134878 137612
rect 134918 137572 134960 137612
rect 135000 137572 149752 137612
rect 149792 137572 149834 137612
rect 149874 137572 149916 137612
rect 149956 137572 149998 137612
rect 150038 137572 150080 137612
rect 150120 137572 152352 137612
rect 71616 137548 152352 137572
rect 71616 136856 152352 136880
rect 71616 136816 75392 136856
rect 75432 136816 75474 136856
rect 75514 136816 75556 136856
rect 75596 136816 75638 136856
rect 75678 136816 75720 136856
rect 75760 136816 90512 136856
rect 90552 136816 90594 136856
rect 90634 136816 90676 136856
rect 90716 136816 90758 136856
rect 90798 136816 90840 136856
rect 90880 136816 105632 136856
rect 105672 136816 105714 136856
rect 105754 136816 105796 136856
rect 105836 136816 105878 136856
rect 105918 136816 105960 136856
rect 106000 136816 120752 136856
rect 120792 136816 120834 136856
rect 120874 136816 120916 136856
rect 120956 136816 120998 136856
rect 121038 136816 121080 136856
rect 121120 136816 135872 136856
rect 135912 136816 135954 136856
rect 135994 136816 136036 136856
rect 136076 136816 136118 136856
rect 136158 136816 136200 136856
rect 136240 136816 150992 136856
rect 151032 136816 151074 136856
rect 151114 136816 151156 136856
rect 151196 136816 151238 136856
rect 151278 136816 151320 136856
rect 151360 136816 152352 136856
rect 71616 136792 152352 136816
rect 71616 136100 152352 136124
rect 71616 136060 74152 136100
rect 74192 136060 74234 136100
rect 74274 136060 74316 136100
rect 74356 136060 74398 136100
rect 74438 136060 74480 136100
rect 74520 136060 89272 136100
rect 89312 136060 89354 136100
rect 89394 136060 89436 136100
rect 89476 136060 89518 136100
rect 89558 136060 89600 136100
rect 89640 136060 104392 136100
rect 104432 136060 104474 136100
rect 104514 136060 104556 136100
rect 104596 136060 104638 136100
rect 104678 136060 104720 136100
rect 104760 136060 119512 136100
rect 119552 136060 119594 136100
rect 119634 136060 119676 136100
rect 119716 136060 119758 136100
rect 119798 136060 119840 136100
rect 119880 136060 134632 136100
rect 134672 136060 134714 136100
rect 134754 136060 134796 136100
rect 134836 136060 134878 136100
rect 134918 136060 134960 136100
rect 135000 136060 149752 136100
rect 149792 136060 149834 136100
rect 149874 136060 149916 136100
rect 149956 136060 149998 136100
rect 150038 136060 150080 136100
rect 150120 136060 152352 136100
rect 71616 136036 152352 136060
rect 71616 135344 152352 135368
rect 71616 135304 75392 135344
rect 75432 135304 75474 135344
rect 75514 135304 75556 135344
rect 75596 135304 75638 135344
rect 75678 135304 75720 135344
rect 75760 135304 90512 135344
rect 90552 135304 90594 135344
rect 90634 135304 90676 135344
rect 90716 135304 90758 135344
rect 90798 135304 90840 135344
rect 90880 135304 105632 135344
rect 105672 135304 105714 135344
rect 105754 135304 105796 135344
rect 105836 135304 105878 135344
rect 105918 135304 105960 135344
rect 106000 135304 120752 135344
rect 120792 135304 120834 135344
rect 120874 135304 120916 135344
rect 120956 135304 120998 135344
rect 121038 135304 121080 135344
rect 121120 135304 135872 135344
rect 135912 135304 135954 135344
rect 135994 135304 136036 135344
rect 136076 135304 136118 135344
rect 136158 135304 136200 135344
rect 136240 135304 150992 135344
rect 151032 135304 151074 135344
rect 151114 135304 151156 135344
rect 151196 135304 151238 135344
rect 151278 135304 151320 135344
rect 151360 135304 152352 135344
rect 71616 135280 152352 135304
rect 71616 134588 152352 134612
rect 71616 134548 74152 134588
rect 74192 134548 74234 134588
rect 74274 134548 74316 134588
rect 74356 134548 74398 134588
rect 74438 134548 74480 134588
rect 74520 134548 89272 134588
rect 89312 134548 89354 134588
rect 89394 134548 89436 134588
rect 89476 134548 89518 134588
rect 89558 134548 89600 134588
rect 89640 134548 104392 134588
rect 104432 134548 104474 134588
rect 104514 134548 104556 134588
rect 104596 134548 104638 134588
rect 104678 134548 104720 134588
rect 104760 134548 119512 134588
rect 119552 134548 119594 134588
rect 119634 134548 119676 134588
rect 119716 134548 119758 134588
rect 119798 134548 119840 134588
rect 119880 134548 134632 134588
rect 134672 134548 134714 134588
rect 134754 134548 134796 134588
rect 134836 134548 134878 134588
rect 134918 134548 134960 134588
rect 135000 134548 149752 134588
rect 149792 134548 149834 134588
rect 149874 134548 149916 134588
rect 149956 134548 149998 134588
rect 150038 134548 150080 134588
rect 150120 134548 152352 134588
rect 71616 134524 152352 134548
rect 71616 133832 152352 133856
rect 71616 133792 75392 133832
rect 75432 133792 75474 133832
rect 75514 133792 75556 133832
rect 75596 133792 75638 133832
rect 75678 133792 75720 133832
rect 75760 133792 90512 133832
rect 90552 133792 90594 133832
rect 90634 133792 90676 133832
rect 90716 133792 90758 133832
rect 90798 133792 90840 133832
rect 90880 133792 105632 133832
rect 105672 133792 105714 133832
rect 105754 133792 105796 133832
rect 105836 133792 105878 133832
rect 105918 133792 105960 133832
rect 106000 133792 120752 133832
rect 120792 133792 120834 133832
rect 120874 133792 120916 133832
rect 120956 133792 120998 133832
rect 121038 133792 121080 133832
rect 121120 133792 135872 133832
rect 135912 133792 135954 133832
rect 135994 133792 136036 133832
rect 136076 133792 136118 133832
rect 136158 133792 136200 133832
rect 136240 133792 150992 133832
rect 151032 133792 151074 133832
rect 151114 133792 151156 133832
rect 151196 133792 151238 133832
rect 151278 133792 151320 133832
rect 151360 133792 152352 133832
rect 71616 133768 152352 133792
rect 71616 133076 152352 133100
rect 71616 133036 74152 133076
rect 74192 133036 74234 133076
rect 74274 133036 74316 133076
rect 74356 133036 74398 133076
rect 74438 133036 74480 133076
rect 74520 133036 89272 133076
rect 89312 133036 89354 133076
rect 89394 133036 89436 133076
rect 89476 133036 89518 133076
rect 89558 133036 89600 133076
rect 89640 133036 104392 133076
rect 104432 133036 104474 133076
rect 104514 133036 104556 133076
rect 104596 133036 104638 133076
rect 104678 133036 104720 133076
rect 104760 133036 119512 133076
rect 119552 133036 119594 133076
rect 119634 133036 119676 133076
rect 119716 133036 119758 133076
rect 119798 133036 119840 133076
rect 119880 133036 134632 133076
rect 134672 133036 134714 133076
rect 134754 133036 134796 133076
rect 134836 133036 134878 133076
rect 134918 133036 134960 133076
rect 135000 133036 149752 133076
rect 149792 133036 149834 133076
rect 149874 133036 149916 133076
rect 149956 133036 149998 133076
rect 150038 133036 150080 133076
rect 150120 133036 152352 133076
rect 71616 133012 152352 133036
rect 71616 132320 152352 132344
rect 71616 132280 75392 132320
rect 75432 132280 75474 132320
rect 75514 132280 75556 132320
rect 75596 132280 75638 132320
rect 75678 132280 75720 132320
rect 75760 132280 90512 132320
rect 90552 132280 90594 132320
rect 90634 132280 90676 132320
rect 90716 132280 90758 132320
rect 90798 132280 90840 132320
rect 90880 132280 105632 132320
rect 105672 132280 105714 132320
rect 105754 132280 105796 132320
rect 105836 132280 105878 132320
rect 105918 132280 105960 132320
rect 106000 132280 120752 132320
rect 120792 132280 120834 132320
rect 120874 132280 120916 132320
rect 120956 132280 120998 132320
rect 121038 132280 121080 132320
rect 121120 132280 135872 132320
rect 135912 132280 135954 132320
rect 135994 132280 136036 132320
rect 136076 132280 136118 132320
rect 136158 132280 136200 132320
rect 136240 132280 150992 132320
rect 151032 132280 151074 132320
rect 151114 132280 151156 132320
rect 151196 132280 151238 132320
rect 151278 132280 151320 132320
rect 151360 132280 152352 132320
rect 71616 132256 152352 132280
rect 71616 131564 152352 131588
rect 71616 131524 74152 131564
rect 74192 131524 74234 131564
rect 74274 131524 74316 131564
rect 74356 131524 74398 131564
rect 74438 131524 74480 131564
rect 74520 131524 89272 131564
rect 89312 131524 89354 131564
rect 89394 131524 89436 131564
rect 89476 131524 89518 131564
rect 89558 131524 89600 131564
rect 89640 131524 104392 131564
rect 104432 131524 104474 131564
rect 104514 131524 104556 131564
rect 104596 131524 104638 131564
rect 104678 131524 104720 131564
rect 104760 131524 119512 131564
rect 119552 131524 119594 131564
rect 119634 131524 119676 131564
rect 119716 131524 119758 131564
rect 119798 131524 119840 131564
rect 119880 131524 134632 131564
rect 134672 131524 134714 131564
rect 134754 131524 134796 131564
rect 134836 131524 134878 131564
rect 134918 131524 134960 131564
rect 135000 131524 149752 131564
rect 149792 131524 149834 131564
rect 149874 131524 149916 131564
rect 149956 131524 149998 131564
rect 150038 131524 150080 131564
rect 150120 131524 152352 131564
rect 71616 131500 152352 131524
rect 71616 130808 152352 130832
rect 71616 130768 75392 130808
rect 75432 130768 75474 130808
rect 75514 130768 75556 130808
rect 75596 130768 75638 130808
rect 75678 130768 75720 130808
rect 75760 130768 90512 130808
rect 90552 130768 90594 130808
rect 90634 130768 90676 130808
rect 90716 130768 90758 130808
rect 90798 130768 90840 130808
rect 90880 130768 105632 130808
rect 105672 130768 105714 130808
rect 105754 130768 105796 130808
rect 105836 130768 105878 130808
rect 105918 130768 105960 130808
rect 106000 130768 120752 130808
rect 120792 130768 120834 130808
rect 120874 130768 120916 130808
rect 120956 130768 120998 130808
rect 121038 130768 121080 130808
rect 121120 130768 135872 130808
rect 135912 130768 135954 130808
rect 135994 130768 136036 130808
rect 136076 130768 136118 130808
rect 136158 130768 136200 130808
rect 136240 130768 150992 130808
rect 151032 130768 151074 130808
rect 151114 130768 151156 130808
rect 151196 130768 151238 130808
rect 151278 130768 151320 130808
rect 151360 130768 152352 130808
rect 71616 130744 152352 130768
rect 71616 130052 152352 130076
rect 71616 130012 74152 130052
rect 74192 130012 74234 130052
rect 74274 130012 74316 130052
rect 74356 130012 74398 130052
rect 74438 130012 74480 130052
rect 74520 130012 89272 130052
rect 89312 130012 89354 130052
rect 89394 130012 89436 130052
rect 89476 130012 89518 130052
rect 89558 130012 89600 130052
rect 89640 130012 104392 130052
rect 104432 130012 104474 130052
rect 104514 130012 104556 130052
rect 104596 130012 104638 130052
rect 104678 130012 104720 130052
rect 104760 130012 119512 130052
rect 119552 130012 119594 130052
rect 119634 130012 119676 130052
rect 119716 130012 119758 130052
rect 119798 130012 119840 130052
rect 119880 130012 134632 130052
rect 134672 130012 134714 130052
rect 134754 130012 134796 130052
rect 134836 130012 134878 130052
rect 134918 130012 134960 130052
rect 135000 130012 149752 130052
rect 149792 130012 149834 130052
rect 149874 130012 149916 130052
rect 149956 130012 149998 130052
rect 150038 130012 150080 130052
rect 150120 130012 152352 130052
rect 71616 129988 152352 130012
rect 71616 129296 152352 129320
rect 71616 129256 75392 129296
rect 75432 129256 75474 129296
rect 75514 129256 75556 129296
rect 75596 129256 75638 129296
rect 75678 129256 75720 129296
rect 75760 129256 90512 129296
rect 90552 129256 90594 129296
rect 90634 129256 90676 129296
rect 90716 129256 90758 129296
rect 90798 129256 90840 129296
rect 90880 129256 105632 129296
rect 105672 129256 105714 129296
rect 105754 129256 105796 129296
rect 105836 129256 105878 129296
rect 105918 129256 105960 129296
rect 106000 129256 120752 129296
rect 120792 129256 120834 129296
rect 120874 129256 120916 129296
rect 120956 129256 120998 129296
rect 121038 129256 121080 129296
rect 121120 129256 135872 129296
rect 135912 129256 135954 129296
rect 135994 129256 136036 129296
rect 136076 129256 136118 129296
rect 136158 129256 136200 129296
rect 136240 129256 150992 129296
rect 151032 129256 151074 129296
rect 151114 129256 151156 129296
rect 151196 129256 151238 129296
rect 151278 129256 151320 129296
rect 151360 129256 152352 129296
rect 71616 129232 152352 129256
rect 71616 128540 152352 128564
rect 71616 128500 74152 128540
rect 74192 128500 74234 128540
rect 74274 128500 74316 128540
rect 74356 128500 74398 128540
rect 74438 128500 74480 128540
rect 74520 128500 89272 128540
rect 89312 128500 89354 128540
rect 89394 128500 89436 128540
rect 89476 128500 89518 128540
rect 89558 128500 89600 128540
rect 89640 128500 104392 128540
rect 104432 128500 104474 128540
rect 104514 128500 104556 128540
rect 104596 128500 104638 128540
rect 104678 128500 104720 128540
rect 104760 128500 119512 128540
rect 119552 128500 119594 128540
rect 119634 128500 119676 128540
rect 119716 128500 119758 128540
rect 119798 128500 119840 128540
rect 119880 128500 134632 128540
rect 134672 128500 134714 128540
rect 134754 128500 134796 128540
rect 134836 128500 134878 128540
rect 134918 128500 134960 128540
rect 135000 128500 149752 128540
rect 149792 128500 149834 128540
rect 149874 128500 149916 128540
rect 149956 128500 149998 128540
rect 150038 128500 150080 128540
rect 150120 128500 152352 128540
rect 71616 128476 152352 128500
rect 71616 127784 152352 127808
rect 71616 127744 75392 127784
rect 75432 127744 75474 127784
rect 75514 127744 75556 127784
rect 75596 127744 75638 127784
rect 75678 127744 75720 127784
rect 75760 127744 90512 127784
rect 90552 127744 90594 127784
rect 90634 127744 90676 127784
rect 90716 127744 90758 127784
rect 90798 127744 90840 127784
rect 90880 127744 105632 127784
rect 105672 127744 105714 127784
rect 105754 127744 105796 127784
rect 105836 127744 105878 127784
rect 105918 127744 105960 127784
rect 106000 127744 120752 127784
rect 120792 127744 120834 127784
rect 120874 127744 120916 127784
rect 120956 127744 120998 127784
rect 121038 127744 121080 127784
rect 121120 127744 135872 127784
rect 135912 127744 135954 127784
rect 135994 127744 136036 127784
rect 136076 127744 136118 127784
rect 136158 127744 136200 127784
rect 136240 127744 150992 127784
rect 151032 127744 151074 127784
rect 151114 127744 151156 127784
rect 151196 127744 151238 127784
rect 151278 127744 151320 127784
rect 151360 127744 152352 127784
rect 71616 127720 152352 127744
rect 71616 127028 152352 127052
rect 71616 126988 74152 127028
rect 74192 126988 74234 127028
rect 74274 126988 74316 127028
rect 74356 126988 74398 127028
rect 74438 126988 74480 127028
rect 74520 126988 89272 127028
rect 89312 126988 89354 127028
rect 89394 126988 89436 127028
rect 89476 126988 89518 127028
rect 89558 126988 89600 127028
rect 89640 126988 104392 127028
rect 104432 126988 104474 127028
rect 104514 126988 104556 127028
rect 104596 126988 104638 127028
rect 104678 126988 104720 127028
rect 104760 126988 119512 127028
rect 119552 126988 119594 127028
rect 119634 126988 119676 127028
rect 119716 126988 119758 127028
rect 119798 126988 119840 127028
rect 119880 126988 134632 127028
rect 134672 126988 134714 127028
rect 134754 126988 134796 127028
rect 134836 126988 134878 127028
rect 134918 126988 134960 127028
rect 135000 126988 149752 127028
rect 149792 126988 149834 127028
rect 149874 126988 149916 127028
rect 149956 126988 149998 127028
rect 150038 126988 150080 127028
rect 150120 126988 152352 127028
rect 71616 126964 152352 126988
rect 71616 126272 152352 126296
rect 71616 126232 75392 126272
rect 75432 126232 75474 126272
rect 75514 126232 75556 126272
rect 75596 126232 75638 126272
rect 75678 126232 75720 126272
rect 75760 126232 90512 126272
rect 90552 126232 90594 126272
rect 90634 126232 90676 126272
rect 90716 126232 90758 126272
rect 90798 126232 90840 126272
rect 90880 126232 105632 126272
rect 105672 126232 105714 126272
rect 105754 126232 105796 126272
rect 105836 126232 105878 126272
rect 105918 126232 105960 126272
rect 106000 126232 120752 126272
rect 120792 126232 120834 126272
rect 120874 126232 120916 126272
rect 120956 126232 120998 126272
rect 121038 126232 121080 126272
rect 121120 126232 135872 126272
rect 135912 126232 135954 126272
rect 135994 126232 136036 126272
rect 136076 126232 136118 126272
rect 136158 126232 136200 126272
rect 136240 126232 150992 126272
rect 151032 126232 151074 126272
rect 151114 126232 151156 126272
rect 151196 126232 151238 126272
rect 151278 126232 151320 126272
rect 151360 126232 152352 126272
rect 71616 126208 152352 126232
rect 71616 125516 152352 125540
rect 71616 125476 74152 125516
rect 74192 125476 74234 125516
rect 74274 125476 74316 125516
rect 74356 125476 74398 125516
rect 74438 125476 74480 125516
rect 74520 125476 89272 125516
rect 89312 125476 89354 125516
rect 89394 125476 89436 125516
rect 89476 125476 89518 125516
rect 89558 125476 89600 125516
rect 89640 125476 104392 125516
rect 104432 125476 104474 125516
rect 104514 125476 104556 125516
rect 104596 125476 104638 125516
rect 104678 125476 104720 125516
rect 104760 125476 119512 125516
rect 119552 125476 119594 125516
rect 119634 125476 119676 125516
rect 119716 125476 119758 125516
rect 119798 125476 119840 125516
rect 119880 125476 134632 125516
rect 134672 125476 134714 125516
rect 134754 125476 134796 125516
rect 134836 125476 134878 125516
rect 134918 125476 134960 125516
rect 135000 125476 149752 125516
rect 149792 125476 149834 125516
rect 149874 125476 149916 125516
rect 149956 125476 149998 125516
rect 150038 125476 150080 125516
rect 150120 125476 152352 125516
rect 71616 125452 152352 125476
rect 71616 124760 152352 124784
rect 71616 124720 75392 124760
rect 75432 124720 75474 124760
rect 75514 124720 75556 124760
rect 75596 124720 75638 124760
rect 75678 124720 75720 124760
rect 75760 124720 90512 124760
rect 90552 124720 90594 124760
rect 90634 124720 90676 124760
rect 90716 124720 90758 124760
rect 90798 124720 90840 124760
rect 90880 124720 105632 124760
rect 105672 124720 105714 124760
rect 105754 124720 105796 124760
rect 105836 124720 105878 124760
rect 105918 124720 105960 124760
rect 106000 124720 120752 124760
rect 120792 124720 120834 124760
rect 120874 124720 120916 124760
rect 120956 124720 120998 124760
rect 121038 124720 121080 124760
rect 121120 124720 135872 124760
rect 135912 124720 135954 124760
rect 135994 124720 136036 124760
rect 136076 124720 136118 124760
rect 136158 124720 136200 124760
rect 136240 124720 150992 124760
rect 151032 124720 151074 124760
rect 151114 124720 151156 124760
rect 151196 124720 151238 124760
rect 151278 124720 151320 124760
rect 151360 124720 152352 124760
rect 71616 124696 152352 124720
rect 71616 124004 152352 124028
rect 71616 123964 74152 124004
rect 74192 123964 74234 124004
rect 74274 123964 74316 124004
rect 74356 123964 74398 124004
rect 74438 123964 74480 124004
rect 74520 123964 89272 124004
rect 89312 123964 89354 124004
rect 89394 123964 89436 124004
rect 89476 123964 89518 124004
rect 89558 123964 89600 124004
rect 89640 123964 104392 124004
rect 104432 123964 104474 124004
rect 104514 123964 104556 124004
rect 104596 123964 104638 124004
rect 104678 123964 104720 124004
rect 104760 123964 119512 124004
rect 119552 123964 119594 124004
rect 119634 123964 119676 124004
rect 119716 123964 119758 124004
rect 119798 123964 119840 124004
rect 119880 123964 134632 124004
rect 134672 123964 134714 124004
rect 134754 123964 134796 124004
rect 134836 123964 134878 124004
rect 134918 123964 134960 124004
rect 135000 123964 149752 124004
rect 149792 123964 149834 124004
rect 149874 123964 149916 124004
rect 149956 123964 149998 124004
rect 150038 123964 150080 124004
rect 150120 123964 152352 124004
rect 71616 123940 152352 123964
rect 71616 123248 152352 123272
rect 71616 123208 75392 123248
rect 75432 123208 75474 123248
rect 75514 123208 75556 123248
rect 75596 123208 75638 123248
rect 75678 123208 75720 123248
rect 75760 123208 90512 123248
rect 90552 123208 90594 123248
rect 90634 123208 90676 123248
rect 90716 123208 90758 123248
rect 90798 123208 90840 123248
rect 90880 123208 105632 123248
rect 105672 123208 105714 123248
rect 105754 123208 105796 123248
rect 105836 123208 105878 123248
rect 105918 123208 105960 123248
rect 106000 123208 120752 123248
rect 120792 123208 120834 123248
rect 120874 123208 120916 123248
rect 120956 123208 120998 123248
rect 121038 123208 121080 123248
rect 121120 123208 135872 123248
rect 135912 123208 135954 123248
rect 135994 123208 136036 123248
rect 136076 123208 136118 123248
rect 136158 123208 136200 123248
rect 136240 123208 150992 123248
rect 151032 123208 151074 123248
rect 151114 123208 151156 123248
rect 151196 123208 151238 123248
rect 151278 123208 151320 123248
rect 151360 123208 152352 123248
rect 71616 123184 152352 123208
rect 71616 122492 152352 122516
rect 71616 122452 74152 122492
rect 74192 122452 74234 122492
rect 74274 122452 74316 122492
rect 74356 122452 74398 122492
rect 74438 122452 74480 122492
rect 74520 122452 89272 122492
rect 89312 122452 89354 122492
rect 89394 122452 89436 122492
rect 89476 122452 89518 122492
rect 89558 122452 89600 122492
rect 89640 122452 104392 122492
rect 104432 122452 104474 122492
rect 104514 122452 104556 122492
rect 104596 122452 104638 122492
rect 104678 122452 104720 122492
rect 104760 122452 119512 122492
rect 119552 122452 119594 122492
rect 119634 122452 119676 122492
rect 119716 122452 119758 122492
rect 119798 122452 119840 122492
rect 119880 122452 134632 122492
rect 134672 122452 134714 122492
rect 134754 122452 134796 122492
rect 134836 122452 134878 122492
rect 134918 122452 134960 122492
rect 135000 122452 149752 122492
rect 149792 122452 149834 122492
rect 149874 122452 149916 122492
rect 149956 122452 149998 122492
rect 150038 122452 150080 122492
rect 150120 122452 152352 122492
rect 71616 122428 152352 122452
rect 71616 121736 152352 121760
rect 71616 121696 75392 121736
rect 75432 121696 75474 121736
rect 75514 121696 75556 121736
rect 75596 121696 75638 121736
rect 75678 121696 75720 121736
rect 75760 121696 90512 121736
rect 90552 121696 90594 121736
rect 90634 121696 90676 121736
rect 90716 121696 90758 121736
rect 90798 121696 90840 121736
rect 90880 121696 105632 121736
rect 105672 121696 105714 121736
rect 105754 121696 105796 121736
rect 105836 121696 105878 121736
rect 105918 121696 105960 121736
rect 106000 121696 120752 121736
rect 120792 121696 120834 121736
rect 120874 121696 120916 121736
rect 120956 121696 120998 121736
rect 121038 121696 121080 121736
rect 121120 121696 135872 121736
rect 135912 121696 135954 121736
rect 135994 121696 136036 121736
rect 136076 121696 136118 121736
rect 136158 121696 136200 121736
rect 136240 121696 150992 121736
rect 151032 121696 151074 121736
rect 151114 121696 151156 121736
rect 151196 121696 151238 121736
rect 151278 121696 151320 121736
rect 151360 121696 152352 121736
rect 71616 121672 152352 121696
rect 71616 120980 152352 121004
rect 71616 120940 74152 120980
rect 74192 120940 74234 120980
rect 74274 120940 74316 120980
rect 74356 120940 74398 120980
rect 74438 120940 74480 120980
rect 74520 120940 89272 120980
rect 89312 120940 89354 120980
rect 89394 120940 89436 120980
rect 89476 120940 89518 120980
rect 89558 120940 89600 120980
rect 89640 120940 104392 120980
rect 104432 120940 104474 120980
rect 104514 120940 104556 120980
rect 104596 120940 104638 120980
rect 104678 120940 104720 120980
rect 104760 120940 119512 120980
rect 119552 120940 119594 120980
rect 119634 120940 119676 120980
rect 119716 120940 119758 120980
rect 119798 120940 119840 120980
rect 119880 120940 134632 120980
rect 134672 120940 134714 120980
rect 134754 120940 134796 120980
rect 134836 120940 134878 120980
rect 134918 120940 134960 120980
rect 135000 120940 149752 120980
rect 149792 120940 149834 120980
rect 149874 120940 149916 120980
rect 149956 120940 149998 120980
rect 150038 120940 150080 120980
rect 150120 120940 152352 120980
rect 71616 120916 152352 120940
rect 71616 120224 152352 120248
rect 71616 120184 75392 120224
rect 75432 120184 75474 120224
rect 75514 120184 75556 120224
rect 75596 120184 75638 120224
rect 75678 120184 75720 120224
rect 75760 120184 90512 120224
rect 90552 120184 90594 120224
rect 90634 120184 90676 120224
rect 90716 120184 90758 120224
rect 90798 120184 90840 120224
rect 90880 120184 105632 120224
rect 105672 120184 105714 120224
rect 105754 120184 105796 120224
rect 105836 120184 105878 120224
rect 105918 120184 105960 120224
rect 106000 120184 120752 120224
rect 120792 120184 120834 120224
rect 120874 120184 120916 120224
rect 120956 120184 120998 120224
rect 121038 120184 121080 120224
rect 121120 120184 135872 120224
rect 135912 120184 135954 120224
rect 135994 120184 136036 120224
rect 136076 120184 136118 120224
rect 136158 120184 136200 120224
rect 136240 120184 150992 120224
rect 151032 120184 151074 120224
rect 151114 120184 151156 120224
rect 151196 120184 151238 120224
rect 151278 120184 151320 120224
rect 151360 120184 152352 120224
rect 71616 120160 152352 120184
rect 71616 119468 152352 119492
rect 71616 119428 74152 119468
rect 74192 119428 74234 119468
rect 74274 119428 74316 119468
rect 74356 119428 74398 119468
rect 74438 119428 74480 119468
rect 74520 119428 89272 119468
rect 89312 119428 89354 119468
rect 89394 119428 89436 119468
rect 89476 119428 89518 119468
rect 89558 119428 89600 119468
rect 89640 119428 104392 119468
rect 104432 119428 104474 119468
rect 104514 119428 104556 119468
rect 104596 119428 104638 119468
rect 104678 119428 104720 119468
rect 104760 119428 119512 119468
rect 119552 119428 119594 119468
rect 119634 119428 119676 119468
rect 119716 119428 119758 119468
rect 119798 119428 119840 119468
rect 119880 119428 134632 119468
rect 134672 119428 134714 119468
rect 134754 119428 134796 119468
rect 134836 119428 134878 119468
rect 134918 119428 134960 119468
rect 135000 119428 149752 119468
rect 149792 119428 149834 119468
rect 149874 119428 149916 119468
rect 149956 119428 149998 119468
rect 150038 119428 150080 119468
rect 150120 119428 152352 119468
rect 71616 119404 152352 119428
rect 71616 118712 152352 118736
rect 71616 118672 75392 118712
rect 75432 118672 75474 118712
rect 75514 118672 75556 118712
rect 75596 118672 75638 118712
rect 75678 118672 75720 118712
rect 75760 118672 90512 118712
rect 90552 118672 90594 118712
rect 90634 118672 90676 118712
rect 90716 118672 90758 118712
rect 90798 118672 90840 118712
rect 90880 118672 105632 118712
rect 105672 118672 105714 118712
rect 105754 118672 105796 118712
rect 105836 118672 105878 118712
rect 105918 118672 105960 118712
rect 106000 118672 120752 118712
rect 120792 118672 120834 118712
rect 120874 118672 120916 118712
rect 120956 118672 120998 118712
rect 121038 118672 121080 118712
rect 121120 118672 135872 118712
rect 135912 118672 135954 118712
rect 135994 118672 136036 118712
rect 136076 118672 136118 118712
rect 136158 118672 136200 118712
rect 136240 118672 150992 118712
rect 151032 118672 151074 118712
rect 151114 118672 151156 118712
rect 151196 118672 151238 118712
rect 151278 118672 151320 118712
rect 151360 118672 152352 118712
rect 71616 118648 152352 118672
rect 71616 117956 152352 117980
rect 71616 117916 74152 117956
rect 74192 117916 74234 117956
rect 74274 117916 74316 117956
rect 74356 117916 74398 117956
rect 74438 117916 74480 117956
rect 74520 117916 89272 117956
rect 89312 117916 89354 117956
rect 89394 117916 89436 117956
rect 89476 117916 89518 117956
rect 89558 117916 89600 117956
rect 89640 117916 104392 117956
rect 104432 117916 104474 117956
rect 104514 117916 104556 117956
rect 104596 117916 104638 117956
rect 104678 117916 104720 117956
rect 104760 117916 119512 117956
rect 119552 117916 119594 117956
rect 119634 117916 119676 117956
rect 119716 117916 119758 117956
rect 119798 117916 119840 117956
rect 119880 117916 134632 117956
rect 134672 117916 134714 117956
rect 134754 117916 134796 117956
rect 134836 117916 134878 117956
rect 134918 117916 134960 117956
rect 135000 117916 149752 117956
rect 149792 117916 149834 117956
rect 149874 117916 149916 117956
rect 149956 117916 149998 117956
rect 150038 117916 150080 117956
rect 150120 117916 152352 117956
rect 71616 117892 152352 117916
rect 71616 117200 152352 117224
rect 71616 117160 75392 117200
rect 75432 117160 75474 117200
rect 75514 117160 75556 117200
rect 75596 117160 75638 117200
rect 75678 117160 75720 117200
rect 75760 117160 90512 117200
rect 90552 117160 90594 117200
rect 90634 117160 90676 117200
rect 90716 117160 90758 117200
rect 90798 117160 90840 117200
rect 90880 117160 105632 117200
rect 105672 117160 105714 117200
rect 105754 117160 105796 117200
rect 105836 117160 105878 117200
rect 105918 117160 105960 117200
rect 106000 117160 120752 117200
rect 120792 117160 120834 117200
rect 120874 117160 120916 117200
rect 120956 117160 120998 117200
rect 121038 117160 121080 117200
rect 121120 117160 135872 117200
rect 135912 117160 135954 117200
rect 135994 117160 136036 117200
rect 136076 117160 136118 117200
rect 136158 117160 136200 117200
rect 136240 117160 150992 117200
rect 151032 117160 151074 117200
rect 151114 117160 151156 117200
rect 151196 117160 151238 117200
rect 151278 117160 151320 117200
rect 151360 117160 152352 117200
rect 71616 117136 152352 117160
rect 71616 116444 152352 116468
rect 71616 116404 74152 116444
rect 74192 116404 74234 116444
rect 74274 116404 74316 116444
rect 74356 116404 74398 116444
rect 74438 116404 74480 116444
rect 74520 116404 89272 116444
rect 89312 116404 89354 116444
rect 89394 116404 89436 116444
rect 89476 116404 89518 116444
rect 89558 116404 89600 116444
rect 89640 116404 104392 116444
rect 104432 116404 104474 116444
rect 104514 116404 104556 116444
rect 104596 116404 104638 116444
rect 104678 116404 104720 116444
rect 104760 116404 119512 116444
rect 119552 116404 119594 116444
rect 119634 116404 119676 116444
rect 119716 116404 119758 116444
rect 119798 116404 119840 116444
rect 119880 116404 134632 116444
rect 134672 116404 134714 116444
rect 134754 116404 134796 116444
rect 134836 116404 134878 116444
rect 134918 116404 134960 116444
rect 135000 116404 149752 116444
rect 149792 116404 149834 116444
rect 149874 116404 149916 116444
rect 149956 116404 149998 116444
rect 150038 116404 150080 116444
rect 150120 116404 152352 116444
rect 71616 116380 152352 116404
rect 71616 115688 152352 115712
rect 71616 115648 75392 115688
rect 75432 115648 75474 115688
rect 75514 115648 75556 115688
rect 75596 115648 75638 115688
rect 75678 115648 75720 115688
rect 75760 115648 90512 115688
rect 90552 115648 90594 115688
rect 90634 115648 90676 115688
rect 90716 115648 90758 115688
rect 90798 115648 90840 115688
rect 90880 115648 105632 115688
rect 105672 115648 105714 115688
rect 105754 115648 105796 115688
rect 105836 115648 105878 115688
rect 105918 115648 105960 115688
rect 106000 115648 120752 115688
rect 120792 115648 120834 115688
rect 120874 115648 120916 115688
rect 120956 115648 120998 115688
rect 121038 115648 121080 115688
rect 121120 115648 135872 115688
rect 135912 115648 135954 115688
rect 135994 115648 136036 115688
rect 136076 115648 136118 115688
rect 136158 115648 136200 115688
rect 136240 115648 150992 115688
rect 151032 115648 151074 115688
rect 151114 115648 151156 115688
rect 151196 115648 151238 115688
rect 151278 115648 151320 115688
rect 151360 115648 152352 115688
rect 71616 115624 152352 115648
rect 71616 114932 152352 114956
rect 71616 114892 74152 114932
rect 74192 114892 74234 114932
rect 74274 114892 74316 114932
rect 74356 114892 74398 114932
rect 74438 114892 74480 114932
rect 74520 114892 89272 114932
rect 89312 114892 89354 114932
rect 89394 114892 89436 114932
rect 89476 114892 89518 114932
rect 89558 114892 89600 114932
rect 89640 114892 104392 114932
rect 104432 114892 104474 114932
rect 104514 114892 104556 114932
rect 104596 114892 104638 114932
rect 104678 114892 104720 114932
rect 104760 114892 119512 114932
rect 119552 114892 119594 114932
rect 119634 114892 119676 114932
rect 119716 114892 119758 114932
rect 119798 114892 119840 114932
rect 119880 114892 134632 114932
rect 134672 114892 134714 114932
rect 134754 114892 134796 114932
rect 134836 114892 134878 114932
rect 134918 114892 134960 114932
rect 135000 114892 149752 114932
rect 149792 114892 149834 114932
rect 149874 114892 149916 114932
rect 149956 114892 149998 114932
rect 150038 114892 150080 114932
rect 150120 114892 152352 114932
rect 71616 114868 152352 114892
rect 71616 114176 152352 114200
rect 71616 114136 75392 114176
rect 75432 114136 75474 114176
rect 75514 114136 75556 114176
rect 75596 114136 75638 114176
rect 75678 114136 75720 114176
rect 75760 114136 90512 114176
rect 90552 114136 90594 114176
rect 90634 114136 90676 114176
rect 90716 114136 90758 114176
rect 90798 114136 90840 114176
rect 90880 114136 105632 114176
rect 105672 114136 105714 114176
rect 105754 114136 105796 114176
rect 105836 114136 105878 114176
rect 105918 114136 105960 114176
rect 106000 114136 120752 114176
rect 120792 114136 120834 114176
rect 120874 114136 120916 114176
rect 120956 114136 120998 114176
rect 121038 114136 121080 114176
rect 121120 114136 135872 114176
rect 135912 114136 135954 114176
rect 135994 114136 136036 114176
rect 136076 114136 136118 114176
rect 136158 114136 136200 114176
rect 136240 114136 150992 114176
rect 151032 114136 151074 114176
rect 151114 114136 151156 114176
rect 151196 114136 151238 114176
rect 151278 114136 151320 114176
rect 151360 114136 152352 114176
rect 71616 114112 152352 114136
rect 71616 113420 152352 113444
rect 71616 113380 74152 113420
rect 74192 113380 74234 113420
rect 74274 113380 74316 113420
rect 74356 113380 74398 113420
rect 74438 113380 74480 113420
rect 74520 113380 89272 113420
rect 89312 113380 89354 113420
rect 89394 113380 89436 113420
rect 89476 113380 89518 113420
rect 89558 113380 89600 113420
rect 89640 113380 104392 113420
rect 104432 113380 104474 113420
rect 104514 113380 104556 113420
rect 104596 113380 104638 113420
rect 104678 113380 104720 113420
rect 104760 113380 119512 113420
rect 119552 113380 119594 113420
rect 119634 113380 119676 113420
rect 119716 113380 119758 113420
rect 119798 113380 119840 113420
rect 119880 113380 134632 113420
rect 134672 113380 134714 113420
rect 134754 113380 134796 113420
rect 134836 113380 134878 113420
rect 134918 113380 134960 113420
rect 135000 113380 149752 113420
rect 149792 113380 149834 113420
rect 149874 113380 149916 113420
rect 149956 113380 149998 113420
rect 150038 113380 150080 113420
rect 150120 113380 152352 113420
rect 71616 113356 152352 113380
rect 71616 112664 152352 112688
rect 71616 112624 75392 112664
rect 75432 112624 75474 112664
rect 75514 112624 75556 112664
rect 75596 112624 75638 112664
rect 75678 112624 75720 112664
rect 75760 112624 90512 112664
rect 90552 112624 90594 112664
rect 90634 112624 90676 112664
rect 90716 112624 90758 112664
rect 90798 112624 90840 112664
rect 90880 112624 105632 112664
rect 105672 112624 105714 112664
rect 105754 112624 105796 112664
rect 105836 112624 105878 112664
rect 105918 112624 105960 112664
rect 106000 112624 120752 112664
rect 120792 112624 120834 112664
rect 120874 112624 120916 112664
rect 120956 112624 120998 112664
rect 121038 112624 121080 112664
rect 121120 112624 135872 112664
rect 135912 112624 135954 112664
rect 135994 112624 136036 112664
rect 136076 112624 136118 112664
rect 136158 112624 136200 112664
rect 136240 112624 150992 112664
rect 151032 112624 151074 112664
rect 151114 112624 151156 112664
rect 151196 112624 151238 112664
rect 151278 112624 151320 112664
rect 151360 112624 152352 112664
rect 71616 112600 152352 112624
rect 71616 111908 152352 111932
rect 71616 111868 74152 111908
rect 74192 111868 74234 111908
rect 74274 111868 74316 111908
rect 74356 111868 74398 111908
rect 74438 111868 74480 111908
rect 74520 111868 89272 111908
rect 89312 111868 89354 111908
rect 89394 111868 89436 111908
rect 89476 111868 89518 111908
rect 89558 111868 89600 111908
rect 89640 111868 104392 111908
rect 104432 111868 104474 111908
rect 104514 111868 104556 111908
rect 104596 111868 104638 111908
rect 104678 111868 104720 111908
rect 104760 111868 119512 111908
rect 119552 111868 119594 111908
rect 119634 111868 119676 111908
rect 119716 111868 119758 111908
rect 119798 111868 119840 111908
rect 119880 111868 134632 111908
rect 134672 111868 134714 111908
rect 134754 111868 134796 111908
rect 134836 111868 134878 111908
rect 134918 111868 134960 111908
rect 135000 111868 149752 111908
rect 149792 111868 149834 111908
rect 149874 111868 149916 111908
rect 149956 111868 149998 111908
rect 150038 111868 150080 111908
rect 150120 111868 152352 111908
rect 71616 111844 152352 111868
rect 71616 111152 152352 111176
rect 71616 111112 75392 111152
rect 75432 111112 75474 111152
rect 75514 111112 75556 111152
rect 75596 111112 75638 111152
rect 75678 111112 75720 111152
rect 75760 111112 90512 111152
rect 90552 111112 90594 111152
rect 90634 111112 90676 111152
rect 90716 111112 90758 111152
rect 90798 111112 90840 111152
rect 90880 111112 105632 111152
rect 105672 111112 105714 111152
rect 105754 111112 105796 111152
rect 105836 111112 105878 111152
rect 105918 111112 105960 111152
rect 106000 111112 120752 111152
rect 120792 111112 120834 111152
rect 120874 111112 120916 111152
rect 120956 111112 120998 111152
rect 121038 111112 121080 111152
rect 121120 111112 135872 111152
rect 135912 111112 135954 111152
rect 135994 111112 136036 111152
rect 136076 111112 136118 111152
rect 136158 111112 136200 111152
rect 136240 111112 150992 111152
rect 151032 111112 151074 111152
rect 151114 111112 151156 111152
rect 151196 111112 151238 111152
rect 151278 111112 151320 111152
rect 151360 111112 152352 111152
rect 71616 111088 152352 111112
rect 71616 110396 152352 110420
rect 71616 110356 74152 110396
rect 74192 110356 74234 110396
rect 74274 110356 74316 110396
rect 74356 110356 74398 110396
rect 74438 110356 74480 110396
rect 74520 110356 89272 110396
rect 89312 110356 89354 110396
rect 89394 110356 89436 110396
rect 89476 110356 89518 110396
rect 89558 110356 89600 110396
rect 89640 110356 104392 110396
rect 104432 110356 104474 110396
rect 104514 110356 104556 110396
rect 104596 110356 104638 110396
rect 104678 110356 104720 110396
rect 104760 110356 119512 110396
rect 119552 110356 119594 110396
rect 119634 110356 119676 110396
rect 119716 110356 119758 110396
rect 119798 110356 119840 110396
rect 119880 110356 134632 110396
rect 134672 110356 134714 110396
rect 134754 110356 134796 110396
rect 134836 110356 134878 110396
rect 134918 110356 134960 110396
rect 135000 110356 149752 110396
rect 149792 110356 149834 110396
rect 149874 110356 149916 110396
rect 149956 110356 149998 110396
rect 150038 110356 150080 110396
rect 150120 110356 152352 110396
rect 71616 110332 152352 110356
rect 71616 109640 152352 109664
rect 71616 109600 75392 109640
rect 75432 109600 75474 109640
rect 75514 109600 75556 109640
rect 75596 109600 75638 109640
rect 75678 109600 75720 109640
rect 75760 109600 90512 109640
rect 90552 109600 90594 109640
rect 90634 109600 90676 109640
rect 90716 109600 90758 109640
rect 90798 109600 90840 109640
rect 90880 109600 105632 109640
rect 105672 109600 105714 109640
rect 105754 109600 105796 109640
rect 105836 109600 105878 109640
rect 105918 109600 105960 109640
rect 106000 109600 120752 109640
rect 120792 109600 120834 109640
rect 120874 109600 120916 109640
rect 120956 109600 120998 109640
rect 121038 109600 121080 109640
rect 121120 109600 135872 109640
rect 135912 109600 135954 109640
rect 135994 109600 136036 109640
rect 136076 109600 136118 109640
rect 136158 109600 136200 109640
rect 136240 109600 150992 109640
rect 151032 109600 151074 109640
rect 151114 109600 151156 109640
rect 151196 109600 151238 109640
rect 151278 109600 151320 109640
rect 151360 109600 152352 109640
rect 71616 109576 152352 109600
rect 71616 108884 152352 108908
rect 71616 108844 74152 108884
rect 74192 108844 74234 108884
rect 74274 108844 74316 108884
rect 74356 108844 74398 108884
rect 74438 108844 74480 108884
rect 74520 108844 89272 108884
rect 89312 108844 89354 108884
rect 89394 108844 89436 108884
rect 89476 108844 89518 108884
rect 89558 108844 89600 108884
rect 89640 108844 104392 108884
rect 104432 108844 104474 108884
rect 104514 108844 104556 108884
rect 104596 108844 104638 108884
rect 104678 108844 104720 108884
rect 104760 108844 119512 108884
rect 119552 108844 119594 108884
rect 119634 108844 119676 108884
rect 119716 108844 119758 108884
rect 119798 108844 119840 108884
rect 119880 108844 134632 108884
rect 134672 108844 134714 108884
rect 134754 108844 134796 108884
rect 134836 108844 134878 108884
rect 134918 108844 134960 108884
rect 135000 108844 149752 108884
rect 149792 108844 149834 108884
rect 149874 108844 149916 108884
rect 149956 108844 149998 108884
rect 150038 108844 150080 108884
rect 150120 108844 152352 108884
rect 71616 108820 152352 108844
rect 71616 108128 152352 108152
rect 71616 108088 75392 108128
rect 75432 108088 75474 108128
rect 75514 108088 75556 108128
rect 75596 108088 75638 108128
rect 75678 108088 75720 108128
rect 75760 108088 90512 108128
rect 90552 108088 90594 108128
rect 90634 108088 90676 108128
rect 90716 108088 90758 108128
rect 90798 108088 90840 108128
rect 90880 108088 105632 108128
rect 105672 108088 105714 108128
rect 105754 108088 105796 108128
rect 105836 108088 105878 108128
rect 105918 108088 105960 108128
rect 106000 108088 120752 108128
rect 120792 108088 120834 108128
rect 120874 108088 120916 108128
rect 120956 108088 120998 108128
rect 121038 108088 121080 108128
rect 121120 108088 135872 108128
rect 135912 108088 135954 108128
rect 135994 108088 136036 108128
rect 136076 108088 136118 108128
rect 136158 108088 136200 108128
rect 136240 108088 150992 108128
rect 151032 108088 151074 108128
rect 151114 108088 151156 108128
rect 151196 108088 151238 108128
rect 151278 108088 151320 108128
rect 151360 108088 152352 108128
rect 71616 108064 152352 108088
rect 71616 107372 152352 107396
rect 71616 107332 74152 107372
rect 74192 107332 74234 107372
rect 74274 107332 74316 107372
rect 74356 107332 74398 107372
rect 74438 107332 74480 107372
rect 74520 107332 89272 107372
rect 89312 107332 89354 107372
rect 89394 107332 89436 107372
rect 89476 107332 89518 107372
rect 89558 107332 89600 107372
rect 89640 107332 104392 107372
rect 104432 107332 104474 107372
rect 104514 107332 104556 107372
rect 104596 107332 104638 107372
rect 104678 107332 104720 107372
rect 104760 107332 119512 107372
rect 119552 107332 119594 107372
rect 119634 107332 119676 107372
rect 119716 107332 119758 107372
rect 119798 107332 119840 107372
rect 119880 107332 134632 107372
rect 134672 107332 134714 107372
rect 134754 107332 134796 107372
rect 134836 107332 134878 107372
rect 134918 107332 134960 107372
rect 135000 107332 149752 107372
rect 149792 107332 149834 107372
rect 149874 107332 149916 107372
rect 149956 107332 149998 107372
rect 150038 107332 150080 107372
rect 150120 107332 152352 107372
rect 71616 107308 152352 107332
rect 71616 106616 152352 106640
rect 71616 106576 75392 106616
rect 75432 106576 75474 106616
rect 75514 106576 75556 106616
rect 75596 106576 75638 106616
rect 75678 106576 75720 106616
rect 75760 106576 90512 106616
rect 90552 106576 90594 106616
rect 90634 106576 90676 106616
rect 90716 106576 90758 106616
rect 90798 106576 90840 106616
rect 90880 106576 105632 106616
rect 105672 106576 105714 106616
rect 105754 106576 105796 106616
rect 105836 106576 105878 106616
rect 105918 106576 105960 106616
rect 106000 106576 120752 106616
rect 120792 106576 120834 106616
rect 120874 106576 120916 106616
rect 120956 106576 120998 106616
rect 121038 106576 121080 106616
rect 121120 106576 135872 106616
rect 135912 106576 135954 106616
rect 135994 106576 136036 106616
rect 136076 106576 136118 106616
rect 136158 106576 136200 106616
rect 136240 106576 150992 106616
rect 151032 106576 151074 106616
rect 151114 106576 151156 106616
rect 151196 106576 151238 106616
rect 151278 106576 151320 106616
rect 151360 106576 152352 106616
rect 71616 106552 152352 106576
rect 71616 105860 152352 105884
rect 71616 105820 74152 105860
rect 74192 105820 74234 105860
rect 74274 105820 74316 105860
rect 74356 105820 74398 105860
rect 74438 105820 74480 105860
rect 74520 105820 89272 105860
rect 89312 105820 89354 105860
rect 89394 105820 89436 105860
rect 89476 105820 89518 105860
rect 89558 105820 89600 105860
rect 89640 105820 104392 105860
rect 104432 105820 104474 105860
rect 104514 105820 104556 105860
rect 104596 105820 104638 105860
rect 104678 105820 104720 105860
rect 104760 105820 119512 105860
rect 119552 105820 119594 105860
rect 119634 105820 119676 105860
rect 119716 105820 119758 105860
rect 119798 105820 119840 105860
rect 119880 105820 134632 105860
rect 134672 105820 134714 105860
rect 134754 105820 134796 105860
rect 134836 105820 134878 105860
rect 134918 105820 134960 105860
rect 135000 105820 149752 105860
rect 149792 105820 149834 105860
rect 149874 105820 149916 105860
rect 149956 105820 149998 105860
rect 150038 105820 150080 105860
rect 150120 105820 152352 105860
rect 71616 105796 152352 105820
rect 71616 105104 152352 105128
rect 71616 105064 75392 105104
rect 75432 105064 75474 105104
rect 75514 105064 75556 105104
rect 75596 105064 75638 105104
rect 75678 105064 75720 105104
rect 75760 105064 90512 105104
rect 90552 105064 90594 105104
rect 90634 105064 90676 105104
rect 90716 105064 90758 105104
rect 90798 105064 90840 105104
rect 90880 105064 105632 105104
rect 105672 105064 105714 105104
rect 105754 105064 105796 105104
rect 105836 105064 105878 105104
rect 105918 105064 105960 105104
rect 106000 105064 120752 105104
rect 120792 105064 120834 105104
rect 120874 105064 120916 105104
rect 120956 105064 120998 105104
rect 121038 105064 121080 105104
rect 121120 105064 135872 105104
rect 135912 105064 135954 105104
rect 135994 105064 136036 105104
rect 136076 105064 136118 105104
rect 136158 105064 136200 105104
rect 136240 105064 150992 105104
rect 151032 105064 151074 105104
rect 151114 105064 151156 105104
rect 151196 105064 151238 105104
rect 151278 105064 151320 105104
rect 151360 105064 152352 105104
rect 71616 105040 152352 105064
rect 71616 104348 152352 104372
rect 71616 104308 74152 104348
rect 74192 104308 74234 104348
rect 74274 104308 74316 104348
rect 74356 104308 74398 104348
rect 74438 104308 74480 104348
rect 74520 104308 89272 104348
rect 89312 104308 89354 104348
rect 89394 104308 89436 104348
rect 89476 104308 89518 104348
rect 89558 104308 89600 104348
rect 89640 104308 104392 104348
rect 104432 104308 104474 104348
rect 104514 104308 104556 104348
rect 104596 104308 104638 104348
rect 104678 104308 104720 104348
rect 104760 104308 119512 104348
rect 119552 104308 119594 104348
rect 119634 104308 119676 104348
rect 119716 104308 119758 104348
rect 119798 104308 119840 104348
rect 119880 104308 134632 104348
rect 134672 104308 134714 104348
rect 134754 104308 134796 104348
rect 134836 104308 134878 104348
rect 134918 104308 134960 104348
rect 135000 104308 149752 104348
rect 149792 104308 149834 104348
rect 149874 104308 149916 104348
rect 149956 104308 149998 104348
rect 150038 104308 150080 104348
rect 150120 104308 152352 104348
rect 71616 104284 152352 104308
rect 71616 103592 152352 103616
rect 71616 103552 75392 103592
rect 75432 103552 75474 103592
rect 75514 103552 75556 103592
rect 75596 103552 75638 103592
rect 75678 103552 75720 103592
rect 75760 103552 90512 103592
rect 90552 103552 90594 103592
rect 90634 103552 90676 103592
rect 90716 103552 90758 103592
rect 90798 103552 90840 103592
rect 90880 103552 105632 103592
rect 105672 103552 105714 103592
rect 105754 103552 105796 103592
rect 105836 103552 105878 103592
rect 105918 103552 105960 103592
rect 106000 103552 120752 103592
rect 120792 103552 120834 103592
rect 120874 103552 120916 103592
rect 120956 103552 120998 103592
rect 121038 103552 121080 103592
rect 121120 103552 135872 103592
rect 135912 103552 135954 103592
rect 135994 103552 136036 103592
rect 136076 103552 136118 103592
rect 136158 103552 136200 103592
rect 136240 103552 150992 103592
rect 151032 103552 151074 103592
rect 151114 103552 151156 103592
rect 151196 103552 151238 103592
rect 151278 103552 151320 103592
rect 151360 103552 152352 103592
rect 71616 103528 152352 103552
rect 71616 102836 152352 102860
rect 71616 102796 74152 102836
rect 74192 102796 74234 102836
rect 74274 102796 74316 102836
rect 74356 102796 74398 102836
rect 74438 102796 74480 102836
rect 74520 102796 89272 102836
rect 89312 102796 89354 102836
rect 89394 102796 89436 102836
rect 89476 102796 89518 102836
rect 89558 102796 89600 102836
rect 89640 102796 104392 102836
rect 104432 102796 104474 102836
rect 104514 102796 104556 102836
rect 104596 102796 104638 102836
rect 104678 102796 104720 102836
rect 104760 102796 119512 102836
rect 119552 102796 119594 102836
rect 119634 102796 119676 102836
rect 119716 102796 119758 102836
rect 119798 102796 119840 102836
rect 119880 102796 134632 102836
rect 134672 102796 134714 102836
rect 134754 102796 134796 102836
rect 134836 102796 134878 102836
rect 134918 102796 134960 102836
rect 135000 102796 149752 102836
rect 149792 102796 149834 102836
rect 149874 102796 149916 102836
rect 149956 102796 149998 102836
rect 150038 102796 150080 102836
rect 150120 102796 152352 102836
rect 71616 102772 152352 102796
rect 71616 102080 152352 102104
rect 71616 102040 75392 102080
rect 75432 102040 75474 102080
rect 75514 102040 75556 102080
rect 75596 102040 75638 102080
rect 75678 102040 75720 102080
rect 75760 102040 90512 102080
rect 90552 102040 90594 102080
rect 90634 102040 90676 102080
rect 90716 102040 90758 102080
rect 90798 102040 90840 102080
rect 90880 102040 105632 102080
rect 105672 102040 105714 102080
rect 105754 102040 105796 102080
rect 105836 102040 105878 102080
rect 105918 102040 105960 102080
rect 106000 102040 120752 102080
rect 120792 102040 120834 102080
rect 120874 102040 120916 102080
rect 120956 102040 120998 102080
rect 121038 102040 121080 102080
rect 121120 102040 135872 102080
rect 135912 102040 135954 102080
rect 135994 102040 136036 102080
rect 136076 102040 136118 102080
rect 136158 102040 136200 102080
rect 136240 102040 150992 102080
rect 151032 102040 151074 102080
rect 151114 102040 151156 102080
rect 151196 102040 151238 102080
rect 151278 102040 151320 102080
rect 151360 102040 152352 102080
rect 71616 102016 152352 102040
rect 71616 101324 152352 101348
rect 71616 101284 74152 101324
rect 74192 101284 74234 101324
rect 74274 101284 74316 101324
rect 74356 101284 74398 101324
rect 74438 101284 74480 101324
rect 74520 101284 89272 101324
rect 89312 101284 89354 101324
rect 89394 101284 89436 101324
rect 89476 101284 89518 101324
rect 89558 101284 89600 101324
rect 89640 101284 104392 101324
rect 104432 101284 104474 101324
rect 104514 101284 104556 101324
rect 104596 101284 104638 101324
rect 104678 101284 104720 101324
rect 104760 101284 119512 101324
rect 119552 101284 119594 101324
rect 119634 101284 119676 101324
rect 119716 101284 119758 101324
rect 119798 101284 119840 101324
rect 119880 101284 134632 101324
rect 134672 101284 134714 101324
rect 134754 101284 134796 101324
rect 134836 101284 134878 101324
rect 134918 101284 134960 101324
rect 135000 101284 149752 101324
rect 149792 101284 149834 101324
rect 149874 101284 149916 101324
rect 149956 101284 149998 101324
rect 150038 101284 150080 101324
rect 150120 101284 152352 101324
rect 71616 101260 152352 101284
rect 71616 100568 152352 100592
rect 71616 100528 75392 100568
rect 75432 100528 75474 100568
rect 75514 100528 75556 100568
rect 75596 100528 75638 100568
rect 75678 100528 75720 100568
rect 75760 100528 90512 100568
rect 90552 100528 90594 100568
rect 90634 100528 90676 100568
rect 90716 100528 90758 100568
rect 90798 100528 90840 100568
rect 90880 100528 105632 100568
rect 105672 100528 105714 100568
rect 105754 100528 105796 100568
rect 105836 100528 105878 100568
rect 105918 100528 105960 100568
rect 106000 100528 120752 100568
rect 120792 100528 120834 100568
rect 120874 100528 120916 100568
rect 120956 100528 120998 100568
rect 121038 100528 121080 100568
rect 121120 100528 135872 100568
rect 135912 100528 135954 100568
rect 135994 100528 136036 100568
rect 136076 100528 136118 100568
rect 136158 100528 136200 100568
rect 136240 100528 150992 100568
rect 151032 100528 151074 100568
rect 151114 100528 151156 100568
rect 151196 100528 151238 100568
rect 151278 100528 151320 100568
rect 151360 100528 152352 100568
rect 71616 100504 152352 100528
rect 71616 99812 152352 99836
rect 71616 99772 74152 99812
rect 74192 99772 74234 99812
rect 74274 99772 74316 99812
rect 74356 99772 74398 99812
rect 74438 99772 74480 99812
rect 74520 99772 89272 99812
rect 89312 99772 89354 99812
rect 89394 99772 89436 99812
rect 89476 99772 89518 99812
rect 89558 99772 89600 99812
rect 89640 99772 104392 99812
rect 104432 99772 104474 99812
rect 104514 99772 104556 99812
rect 104596 99772 104638 99812
rect 104678 99772 104720 99812
rect 104760 99772 119512 99812
rect 119552 99772 119594 99812
rect 119634 99772 119676 99812
rect 119716 99772 119758 99812
rect 119798 99772 119840 99812
rect 119880 99772 134632 99812
rect 134672 99772 134714 99812
rect 134754 99772 134796 99812
rect 134836 99772 134878 99812
rect 134918 99772 134960 99812
rect 135000 99772 149752 99812
rect 149792 99772 149834 99812
rect 149874 99772 149916 99812
rect 149956 99772 149998 99812
rect 150038 99772 150080 99812
rect 150120 99772 152352 99812
rect 71616 99748 152352 99772
rect 71616 99056 152352 99080
rect 71616 99016 75392 99056
rect 75432 99016 75474 99056
rect 75514 99016 75556 99056
rect 75596 99016 75638 99056
rect 75678 99016 75720 99056
rect 75760 99016 90512 99056
rect 90552 99016 90594 99056
rect 90634 99016 90676 99056
rect 90716 99016 90758 99056
rect 90798 99016 90840 99056
rect 90880 99016 105632 99056
rect 105672 99016 105714 99056
rect 105754 99016 105796 99056
rect 105836 99016 105878 99056
rect 105918 99016 105960 99056
rect 106000 99016 120752 99056
rect 120792 99016 120834 99056
rect 120874 99016 120916 99056
rect 120956 99016 120998 99056
rect 121038 99016 121080 99056
rect 121120 99016 135872 99056
rect 135912 99016 135954 99056
rect 135994 99016 136036 99056
rect 136076 99016 136118 99056
rect 136158 99016 136200 99056
rect 136240 99016 150992 99056
rect 151032 99016 151074 99056
rect 151114 99016 151156 99056
rect 151196 99016 151238 99056
rect 151278 99016 151320 99056
rect 151360 99016 152352 99056
rect 71616 98992 152352 99016
rect 71616 98300 152352 98324
rect 71616 98260 74152 98300
rect 74192 98260 74234 98300
rect 74274 98260 74316 98300
rect 74356 98260 74398 98300
rect 74438 98260 74480 98300
rect 74520 98260 89272 98300
rect 89312 98260 89354 98300
rect 89394 98260 89436 98300
rect 89476 98260 89518 98300
rect 89558 98260 89600 98300
rect 89640 98260 104392 98300
rect 104432 98260 104474 98300
rect 104514 98260 104556 98300
rect 104596 98260 104638 98300
rect 104678 98260 104720 98300
rect 104760 98260 119512 98300
rect 119552 98260 119594 98300
rect 119634 98260 119676 98300
rect 119716 98260 119758 98300
rect 119798 98260 119840 98300
rect 119880 98260 134632 98300
rect 134672 98260 134714 98300
rect 134754 98260 134796 98300
rect 134836 98260 134878 98300
rect 134918 98260 134960 98300
rect 135000 98260 149752 98300
rect 149792 98260 149834 98300
rect 149874 98260 149916 98300
rect 149956 98260 149998 98300
rect 150038 98260 150080 98300
rect 150120 98260 152352 98300
rect 71616 98236 152352 98260
rect 71616 97544 152352 97568
rect 71616 97504 75392 97544
rect 75432 97504 75474 97544
rect 75514 97504 75556 97544
rect 75596 97504 75638 97544
rect 75678 97504 75720 97544
rect 75760 97504 90512 97544
rect 90552 97504 90594 97544
rect 90634 97504 90676 97544
rect 90716 97504 90758 97544
rect 90798 97504 90840 97544
rect 90880 97504 105632 97544
rect 105672 97504 105714 97544
rect 105754 97504 105796 97544
rect 105836 97504 105878 97544
rect 105918 97504 105960 97544
rect 106000 97504 120752 97544
rect 120792 97504 120834 97544
rect 120874 97504 120916 97544
rect 120956 97504 120998 97544
rect 121038 97504 121080 97544
rect 121120 97504 135872 97544
rect 135912 97504 135954 97544
rect 135994 97504 136036 97544
rect 136076 97504 136118 97544
rect 136158 97504 136200 97544
rect 136240 97504 150992 97544
rect 151032 97504 151074 97544
rect 151114 97504 151156 97544
rect 151196 97504 151238 97544
rect 151278 97504 151320 97544
rect 151360 97504 152352 97544
rect 71616 97480 152352 97504
rect 71616 96788 152352 96812
rect 71616 96748 74152 96788
rect 74192 96748 74234 96788
rect 74274 96748 74316 96788
rect 74356 96748 74398 96788
rect 74438 96748 74480 96788
rect 74520 96748 89272 96788
rect 89312 96748 89354 96788
rect 89394 96748 89436 96788
rect 89476 96748 89518 96788
rect 89558 96748 89600 96788
rect 89640 96748 104392 96788
rect 104432 96748 104474 96788
rect 104514 96748 104556 96788
rect 104596 96748 104638 96788
rect 104678 96748 104720 96788
rect 104760 96748 119512 96788
rect 119552 96748 119594 96788
rect 119634 96748 119676 96788
rect 119716 96748 119758 96788
rect 119798 96748 119840 96788
rect 119880 96748 134632 96788
rect 134672 96748 134714 96788
rect 134754 96748 134796 96788
rect 134836 96748 134878 96788
rect 134918 96748 134960 96788
rect 135000 96748 149752 96788
rect 149792 96748 149834 96788
rect 149874 96748 149916 96788
rect 149956 96748 149998 96788
rect 150038 96748 150080 96788
rect 150120 96748 152352 96788
rect 71616 96724 152352 96748
rect 71616 96032 152352 96056
rect 71616 95992 75392 96032
rect 75432 95992 75474 96032
rect 75514 95992 75556 96032
rect 75596 95992 75638 96032
rect 75678 95992 75720 96032
rect 75760 95992 90512 96032
rect 90552 95992 90594 96032
rect 90634 95992 90676 96032
rect 90716 95992 90758 96032
rect 90798 95992 90840 96032
rect 90880 95992 105632 96032
rect 105672 95992 105714 96032
rect 105754 95992 105796 96032
rect 105836 95992 105878 96032
rect 105918 95992 105960 96032
rect 106000 95992 120752 96032
rect 120792 95992 120834 96032
rect 120874 95992 120916 96032
rect 120956 95992 120998 96032
rect 121038 95992 121080 96032
rect 121120 95992 135872 96032
rect 135912 95992 135954 96032
rect 135994 95992 136036 96032
rect 136076 95992 136118 96032
rect 136158 95992 136200 96032
rect 136240 95992 150992 96032
rect 151032 95992 151074 96032
rect 151114 95992 151156 96032
rect 151196 95992 151238 96032
rect 151278 95992 151320 96032
rect 151360 95992 152352 96032
rect 71616 95968 152352 95992
rect 71616 95276 152352 95300
rect 71616 95236 74152 95276
rect 74192 95236 74234 95276
rect 74274 95236 74316 95276
rect 74356 95236 74398 95276
rect 74438 95236 74480 95276
rect 74520 95236 89272 95276
rect 89312 95236 89354 95276
rect 89394 95236 89436 95276
rect 89476 95236 89518 95276
rect 89558 95236 89600 95276
rect 89640 95236 104392 95276
rect 104432 95236 104474 95276
rect 104514 95236 104556 95276
rect 104596 95236 104638 95276
rect 104678 95236 104720 95276
rect 104760 95236 119512 95276
rect 119552 95236 119594 95276
rect 119634 95236 119676 95276
rect 119716 95236 119758 95276
rect 119798 95236 119840 95276
rect 119880 95236 134632 95276
rect 134672 95236 134714 95276
rect 134754 95236 134796 95276
rect 134836 95236 134878 95276
rect 134918 95236 134960 95276
rect 135000 95236 149752 95276
rect 149792 95236 149834 95276
rect 149874 95236 149916 95276
rect 149956 95236 149998 95276
rect 150038 95236 150080 95276
rect 150120 95236 152352 95276
rect 71616 95212 152352 95236
rect 71616 94520 152352 94544
rect 71616 94480 75392 94520
rect 75432 94480 75474 94520
rect 75514 94480 75556 94520
rect 75596 94480 75638 94520
rect 75678 94480 75720 94520
rect 75760 94480 90512 94520
rect 90552 94480 90594 94520
rect 90634 94480 90676 94520
rect 90716 94480 90758 94520
rect 90798 94480 90840 94520
rect 90880 94480 105632 94520
rect 105672 94480 105714 94520
rect 105754 94480 105796 94520
rect 105836 94480 105878 94520
rect 105918 94480 105960 94520
rect 106000 94480 120752 94520
rect 120792 94480 120834 94520
rect 120874 94480 120916 94520
rect 120956 94480 120998 94520
rect 121038 94480 121080 94520
rect 121120 94480 135872 94520
rect 135912 94480 135954 94520
rect 135994 94480 136036 94520
rect 136076 94480 136118 94520
rect 136158 94480 136200 94520
rect 136240 94480 150992 94520
rect 151032 94480 151074 94520
rect 151114 94480 151156 94520
rect 151196 94480 151238 94520
rect 151278 94480 151320 94520
rect 151360 94480 152352 94520
rect 71616 94456 152352 94480
rect 71616 93764 152352 93788
rect 71616 93724 74152 93764
rect 74192 93724 74234 93764
rect 74274 93724 74316 93764
rect 74356 93724 74398 93764
rect 74438 93724 74480 93764
rect 74520 93724 89272 93764
rect 89312 93724 89354 93764
rect 89394 93724 89436 93764
rect 89476 93724 89518 93764
rect 89558 93724 89600 93764
rect 89640 93724 104392 93764
rect 104432 93724 104474 93764
rect 104514 93724 104556 93764
rect 104596 93724 104638 93764
rect 104678 93724 104720 93764
rect 104760 93724 119512 93764
rect 119552 93724 119594 93764
rect 119634 93724 119676 93764
rect 119716 93724 119758 93764
rect 119798 93724 119840 93764
rect 119880 93724 134632 93764
rect 134672 93724 134714 93764
rect 134754 93724 134796 93764
rect 134836 93724 134878 93764
rect 134918 93724 134960 93764
rect 135000 93724 149752 93764
rect 149792 93724 149834 93764
rect 149874 93724 149916 93764
rect 149956 93724 149998 93764
rect 150038 93724 150080 93764
rect 150120 93724 152352 93764
rect 71616 93700 152352 93724
rect 71616 93008 152352 93032
rect 71616 92968 75392 93008
rect 75432 92968 75474 93008
rect 75514 92968 75556 93008
rect 75596 92968 75638 93008
rect 75678 92968 75720 93008
rect 75760 92968 90512 93008
rect 90552 92968 90594 93008
rect 90634 92968 90676 93008
rect 90716 92968 90758 93008
rect 90798 92968 90840 93008
rect 90880 92968 105632 93008
rect 105672 92968 105714 93008
rect 105754 92968 105796 93008
rect 105836 92968 105878 93008
rect 105918 92968 105960 93008
rect 106000 92968 120752 93008
rect 120792 92968 120834 93008
rect 120874 92968 120916 93008
rect 120956 92968 120998 93008
rect 121038 92968 121080 93008
rect 121120 92968 135872 93008
rect 135912 92968 135954 93008
rect 135994 92968 136036 93008
rect 136076 92968 136118 93008
rect 136158 92968 136200 93008
rect 136240 92968 150992 93008
rect 151032 92968 151074 93008
rect 151114 92968 151156 93008
rect 151196 92968 151238 93008
rect 151278 92968 151320 93008
rect 151360 92968 152352 93008
rect 71616 92944 152352 92968
rect 71616 92252 152352 92276
rect 71616 92212 74152 92252
rect 74192 92212 74234 92252
rect 74274 92212 74316 92252
rect 74356 92212 74398 92252
rect 74438 92212 74480 92252
rect 74520 92212 89272 92252
rect 89312 92212 89354 92252
rect 89394 92212 89436 92252
rect 89476 92212 89518 92252
rect 89558 92212 89600 92252
rect 89640 92212 104392 92252
rect 104432 92212 104474 92252
rect 104514 92212 104556 92252
rect 104596 92212 104638 92252
rect 104678 92212 104720 92252
rect 104760 92212 119512 92252
rect 119552 92212 119594 92252
rect 119634 92212 119676 92252
rect 119716 92212 119758 92252
rect 119798 92212 119840 92252
rect 119880 92212 134632 92252
rect 134672 92212 134714 92252
rect 134754 92212 134796 92252
rect 134836 92212 134878 92252
rect 134918 92212 134960 92252
rect 135000 92212 149752 92252
rect 149792 92212 149834 92252
rect 149874 92212 149916 92252
rect 149956 92212 149998 92252
rect 150038 92212 150080 92252
rect 150120 92212 152352 92252
rect 71616 92188 152352 92212
rect 71616 91496 152352 91520
rect 71616 91456 75392 91496
rect 75432 91456 75474 91496
rect 75514 91456 75556 91496
rect 75596 91456 75638 91496
rect 75678 91456 75720 91496
rect 75760 91456 90512 91496
rect 90552 91456 90594 91496
rect 90634 91456 90676 91496
rect 90716 91456 90758 91496
rect 90798 91456 90840 91496
rect 90880 91456 105632 91496
rect 105672 91456 105714 91496
rect 105754 91456 105796 91496
rect 105836 91456 105878 91496
rect 105918 91456 105960 91496
rect 106000 91456 120752 91496
rect 120792 91456 120834 91496
rect 120874 91456 120916 91496
rect 120956 91456 120998 91496
rect 121038 91456 121080 91496
rect 121120 91456 135872 91496
rect 135912 91456 135954 91496
rect 135994 91456 136036 91496
rect 136076 91456 136118 91496
rect 136158 91456 136200 91496
rect 136240 91456 150992 91496
rect 151032 91456 151074 91496
rect 151114 91456 151156 91496
rect 151196 91456 151238 91496
rect 151278 91456 151320 91496
rect 151360 91456 152352 91496
rect 71616 91432 152352 91456
rect 71616 90740 152352 90764
rect 71616 90700 74152 90740
rect 74192 90700 74234 90740
rect 74274 90700 74316 90740
rect 74356 90700 74398 90740
rect 74438 90700 74480 90740
rect 74520 90700 89272 90740
rect 89312 90700 89354 90740
rect 89394 90700 89436 90740
rect 89476 90700 89518 90740
rect 89558 90700 89600 90740
rect 89640 90700 104392 90740
rect 104432 90700 104474 90740
rect 104514 90700 104556 90740
rect 104596 90700 104638 90740
rect 104678 90700 104720 90740
rect 104760 90700 119512 90740
rect 119552 90700 119594 90740
rect 119634 90700 119676 90740
rect 119716 90700 119758 90740
rect 119798 90700 119840 90740
rect 119880 90700 134632 90740
rect 134672 90700 134714 90740
rect 134754 90700 134796 90740
rect 134836 90700 134878 90740
rect 134918 90700 134960 90740
rect 135000 90700 149752 90740
rect 149792 90700 149834 90740
rect 149874 90700 149916 90740
rect 149956 90700 149998 90740
rect 150038 90700 150080 90740
rect 150120 90700 152352 90740
rect 71616 90676 152352 90700
rect 71616 89984 152352 90008
rect 71616 89944 75392 89984
rect 75432 89944 75474 89984
rect 75514 89944 75556 89984
rect 75596 89944 75638 89984
rect 75678 89944 75720 89984
rect 75760 89944 90512 89984
rect 90552 89944 90594 89984
rect 90634 89944 90676 89984
rect 90716 89944 90758 89984
rect 90798 89944 90840 89984
rect 90880 89944 105632 89984
rect 105672 89944 105714 89984
rect 105754 89944 105796 89984
rect 105836 89944 105878 89984
rect 105918 89944 105960 89984
rect 106000 89944 120752 89984
rect 120792 89944 120834 89984
rect 120874 89944 120916 89984
rect 120956 89944 120998 89984
rect 121038 89944 121080 89984
rect 121120 89944 135872 89984
rect 135912 89944 135954 89984
rect 135994 89944 136036 89984
rect 136076 89944 136118 89984
rect 136158 89944 136200 89984
rect 136240 89944 150992 89984
rect 151032 89944 151074 89984
rect 151114 89944 151156 89984
rect 151196 89944 151238 89984
rect 151278 89944 151320 89984
rect 151360 89944 152352 89984
rect 71616 89920 152352 89944
rect 71616 89228 152352 89252
rect 71616 89188 74152 89228
rect 74192 89188 74234 89228
rect 74274 89188 74316 89228
rect 74356 89188 74398 89228
rect 74438 89188 74480 89228
rect 74520 89188 89272 89228
rect 89312 89188 89354 89228
rect 89394 89188 89436 89228
rect 89476 89188 89518 89228
rect 89558 89188 89600 89228
rect 89640 89188 104392 89228
rect 104432 89188 104474 89228
rect 104514 89188 104556 89228
rect 104596 89188 104638 89228
rect 104678 89188 104720 89228
rect 104760 89188 119512 89228
rect 119552 89188 119594 89228
rect 119634 89188 119676 89228
rect 119716 89188 119758 89228
rect 119798 89188 119840 89228
rect 119880 89188 134632 89228
rect 134672 89188 134714 89228
rect 134754 89188 134796 89228
rect 134836 89188 134878 89228
rect 134918 89188 134960 89228
rect 135000 89188 149752 89228
rect 149792 89188 149834 89228
rect 149874 89188 149916 89228
rect 149956 89188 149998 89228
rect 150038 89188 150080 89228
rect 150120 89188 152352 89228
rect 71616 89164 152352 89188
rect 71616 88472 152352 88496
rect 71616 88432 75392 88472
rect 75432 88432 75474 88472
rect 75514 88432 75556 88472
rect 75596 88432 75638 88472
rect 75678 88432 75720 88472
rect 75760 88432 90512 88472
rect 90552 88432 90594 88472
rect 90634 88432 90676 88472
rect 90716 88432 90758 88472
rect 90798 88432 90840 88472
rect 90880 88432 105632 88472
rect 105672 88432 105714 88472
rect 105754 88432 105796 88472
rect 105836 88432 105878 88472
rect 105918 88432 105960 88472
rect 106000 88432 120752 88472
rect 120792 88432 120834 88472
rect 120874 88432 120916 88472
rect 120956 88432 120998 88472
rect 121038 88432 121080 88472
rect 121120 88432 135872 88472
rect 135912 88432 135954 88472
rect 135994 88432 136036 88472
rect 136076 88432 136118 88472
rect 136158 88432 136200 88472
rect 136240 88432 150992 88472
rect 151032 88432 151074 88472
rect 151114 88432 151156 88472
rect 151196 88432 151238 88472
rect 151278 88432 151320 88472
rect 151360 88432 152352 88472
rect 71616 88408 152352 88432
rect 71616 87716 152352 87740
rect 71616 87676 74152 87716
rect 74192 87676 74234 87716
rect 74274 87676 74316 87716
rect 74356 87676 74398 87716
rect 74438 87676 74480 87716
rect 74520 87676 89272 87716
rect 89312 87676 89354 87716
rect 89394 87676 89436 87716
rect 89476 87676 89518 87716
rect 89558 87676 89600 87716
rect 89640 87676 104392 87716
rect 104432 87676 104474 87716
rect 104514 87676 104556 87716
rect 104596 87676 104638 87716
rect 104678 87676 104720 87716
rect 104760 87676 119512 87716
rect 119552 87676 119594 87716
rect 119634 87676 119676 87716
rect 119716 87676 119758 87716
rect 119798 87676 119840 87716
rect 119880 87676 134632 87716
rect 134672 87676 134714 87716
rect 134754 87676 134796 87716
rect 134836 87676 134878 87716
rect 134918 87676 134960 87716
rect 135000 87676 149752 87716
rect 149792 87676 149834 87716
rect 149874 87676 149916 87716
rect 149956 87676 149998 87716
rect 150038 87676 150080 87716
rect 150120 87676 152352 87716
rect 71616 87652 152352 87676
rect 71616 86960 152352 86984
rect 71616 86920 75392 86960
rect 75432 86920 75474 86960
rect 75514 86920 75556 86960
rect 75596 86920 75638 86960
rect 75678 86920 75720 86960
rect 75760 86920 90512 86960
rect 90552 86920 90594 86960
rect 90634 86920 90676 86960
rect 90716 86920 90758 86960
rect 90798 86920 90840 86960
rect 90880 86920 105632 86960
rect 105672 86920 105714 86960
rect 105754 86920 105796 86960
rect 105836 86920 105878 86960
rect 105918 86920 105960 86960
rect 106000 86920 120752 86960
rect 120792 86920 120834 86960
rect 120874 86920 120916 86960
rect 120956 86920 120998 86960
rect 121038 86920 121080 86960
rect 121120 86920 135872 86960
rect 135912 86920 135954 86960
rect 135994 86920 136036 86960
rect 136076 86920 136118 86960
rect 136158 86920 136200 86960
rect 136240 86920 150992 86960
rect 151032 86920 151074 86960
rect 151114 86920 151156 86960
rect 151196 86920 151238 86960
rect 151278 86920 151320 86960
rect 151360 86920 152352 86960
rect 71616 86896 152352 86920
rect 71616 86204 152352 86228
rect 71616 86164 74152 86204
rect 74192 86164 74234 86204
rect 74274 86164 74316 86204
rect 74356 86164 74398 86204
rect 74438 86164 74480 86204
rect 74520 86164 89272 86204
rect 89312 86164 89354 86204
rect 89394 86164 89436 86204
rect 89476 86164 89518 86204
rect 89558 86164 89600 86204
rect 89640 86164 104392 86204
rect 104432 86164 104474 86204
rect 104514 86164 104556 86204
rect 104596 86164 104638 86204
rect 104678 86164 104720 86204
rect 104760 86164 119512 86204
rect 119552 86164 119594 86204
rect 119634 86164 119676 86204
rect 119716 86164 119758 86204
rect 119798 86164 119840 86204
rect 119880 86164 134632 86204
rect 134672 86164 134714 86204
rect 134754 86164 134796 86204
rect 134836 86164 134878 86204
rect 134918 86164 134960 86204
rect 135000 86164 149752 86204
rect 149792 86164 149834 86204
rect 149874 86164 149916 86204
rect 149956 86164 149998 86204
rect 150038 86164 150080 86204
rect 150120 86164 152352 86204
rect 71616 86140 152352 86164
rect 71616 85448 152352 85472
rect 71616 85408 75392 85448
rect 75432 85408 75474 85448
rect 75514 85408 75556 85448
rect 75596 85408 75638 85448
rect 75678 85408 75720 85448
rect 75760 85408 90512 85448
rect 90552 85408 90594 85448
rect 90634 85408 90676 85448
rect 90716 85408 90758 85448
rect 90798 85408 90840 85448
rect 90880 85408 105632 85448
rect 105672 85408 105714 85448
rect 105754 85408 105796 85448
rect 105836 85408 105878 85448
rect 105918 85408 105960 85448
rect 106000 85408 120752 85448
rect 120792 85408 120834 85448
rect 120874 85408 120916 85448
rect 120956 85408 120998 85448
rect 121038 85408 121080 85448
rect 121120 85408 135872 85448
rect 135912 85408 135954 85448
rect 135994 85408 136036 85448
rect 136076 85408 136118 85448
rect 136158 85408 136200 85448
rect 136240 85408 150992 85448
rect 151032 85408 151074 85448
rect 151114 85408 151156 85448
rect 151196 85408 151238 85448
rect 151278 85408 151320 85448
rect 151360 85408 152352 85448
rect 71616 85384 152352 85408
rect 71616 84692 152352 84716
rect 71616 84652 74152 84692
rect 74192 84652 74234 84692
rect 74274 84652 74316 84692
rect 74356 84652 74398 84692
rect 74438 84652 74480 84692
rect 74520 84652 89272 84692
rect 89312 84652 89354 84692
rect 89394 84652 89436 84692
rect 89476 84652 89518 84692
rect 89558 84652 89600 84692
rect 89640 84652 104392 84692
rect 104432 84652 104474 84692
rect 104514 84652 104556 84692
rect 104596 84652 104638 84692
rect 104678 84652 104720 84692
rect 104760 84652 119512 84692
rect 119552 84652 119594 84692
rect 119634 84652 119676 84692
rect 119716 84652 119758 84692
rect 119798 84652 119840 84692
rect 119880 84652 134632 84692
rect 134672 84652 134714 84692
rect 134754 84652 134796 84692
rect 134836 84652 134878 84692
rect 134918 84652 134960 84692
rect 135000 84652 149752 84692
rect 149792 84652 149834 84692
rect 149874 84652 149916 84692
rect 149956 84652 149998 84692
rect 150038 84652 150080 84692
rect 150120 84652 152352 84692
rect 71616 84628 152352 84652
rect 71616 83936 152352 83960
rect 71616 83896 75392 83936
rect 75432 83896 75474 83936
rect 75514 83896 75556 83936
rect 75596 83896 75638 83936
rect 75678 83896 75720 83936
rect 75760 83896 90512 83936
rect 90552 83896 90594 83936
rect 90634 83896 90676 83936
rect 90716 83896 90758 83936
rect 90798 83896 90840 83936
rect 90880 83896 105632 83936
rect 105672 83896 105714 83936
rect 105754 83896 105796 83936
rect 105836 83896 105878 83936
rect 105918 83896 105960 83936
rect 106000 83896 120752 83936
rect 120792 83896 120834 83936
rect 120874 83896 120916 83936
rect 120956 83896 120998 83936
rect 121038 83896 121080 83936
rect 121120 83896 135872 83936
rect 135912 83896 135954 83936
rect 135994 83896 136036 83936
rect 136076 83896 136118 83936
rect 136158 83896 136200 83936
rect 136240 83896 150992 83936
rect 151032 83896 151074 83936
rect 151114 83896 151156 83936
rect 151196 83896 151238 83936
rect 151278 83896 151320 83936
rect 151360 83896 152352 83936
rect 71616 83872 152352 83896
rect 71616 83180 152352 83204
rect 71616 83140 74152 83180
rect 74192 83140 74234 83180
rect 74274 83140 74316 83180
rect 74356 83140 74398 83180
rect 74438 83140 74480 83180
rect 74520 83140 89272 83180
rect 89312 83140 89354 83180
rect 89394 83140 89436 83180
rect 89476 83140 89518 83180
rect 89558 83140 89600 83180
rect 89640 83140 104392 83180
rect 104432 83140 104474 83180
rect 104514 83140 104556 83180
rect 104596 83140 104638 83180
rect 104678 83140 104720 83180
rect 104760 83140 119512 83180
rect 119552 83140 119594 83180
rect 119634 83140 119676 83180
rect 119716 83140 119758 83180
rect 119798 83140 119840 83180
rect 119880 83140 134632 83180
rect 134672 83140 134714 83180
rect 134754 83140 134796 83180
rect 134836 83140 134878 83180
rect 134918 83140 134960 83180
rect 135000 83140 149752 83180
rect 149792 83140 149834 83180
rect 149874 83140 149916 83180
rect 149956 83140 149998 83180
rect 150038 83140 150080 83180
rect 150120 83140 152352 83180
rect 71616 83116 152352 83140
rect 71616 82424 152352 82448
rect 71616 82384 75392 82424
rect 75432 82384 75474 82424
rect 75514 82384 75556 82424
rect 75596 82384 75638 82424
rect 75678 82384 75720 82424
rect 75760 82384 90512 82424
rect 90552 82384 90594 82424
rect 90634 82384 90676 82424
rect 90716 82384 90758 82424
rect 90798 82384 90840 82424
rect 90880 82384 105632 82424
rect 105672 82384 105714 82424
rect 105754 82384 105796 82424
rect 105836 82384 105878 82424
rect 105918 82384 105960 82424
rect 106000 82384 120752 82424
rect 120792 82384 120834 82424
rect 120874 82384 120916 82424
rect 120956 82384 120998 82424
rect 121038 82384 121080 82424
rect 121120 82384 135872 82424
rect 135912 82384 135954 82424
rect 135994 82384 136036 82424
rect 136076 82384 136118 82424
rect 136158 82384 136200 82424
rect 136240 82384 150992 82424
rect 151032 82384 151074 82424
rect 151114 82384 151156 82424
rect 151196 82384 151238 82424
rect 151278 82384 151320 82424
rect 151360 82384 152352 82424
rect 71616 82360 152352 82384
rect 71616 81668 152352 81692
rect 71616 81628 74152 81668
rect 74192 81628 74234 81668
rect 74274 81628 74316 81668
rect 74356 81628 74398 81668
rect 74438 81628 74480 81668
rect 74520 81628 89272 81668
rect 89312 81628 89354 81668
rect 89394 81628 89436 81668
rect 89476 81628 89518 81668
rect 89558 81628 89600 81668
rect 89640 81628 104392 81668
rect 104432 81628 104474 81668
rect 104514 81628 104556 81668
rect 104596 81628 104638 81668
rect 104678 81628 104720 81668
rect 104760 81628 119512 81668
rect 119552 81628 119594 81668
rect 119634 81628 119676 81668
rect 119716 81628 119758 81668
rect 119798 81628 119840 81668
rect 119880 81628 134632 81668
rect 134672 81628 134714 81668
rect 134754 81628 134796 81668
rect 134836 81628 134878 81668
rect 134918 81628 134960 81668
rect 135000 81628 149752 81668
rect 149792 81628 149834 81668
rect 149874 81628 149916 81668
rect 149956 81628 149998 81668
rect 150038 81628 150080 81668
rect 150120 81628 152352 81668
rect 71616 81604 152352 81628
rect 71616 80912 152352 80936
rect 71616 80872 75392 80912
rect 75432 80872 75474 80912
rect 75514 80872 75556 80912
rect 75596 80872 75638 80912
rect 75678 80872 75720 80912
rect 75760 80872 90512 80912
rect 90552 80872 90594 80912
rect 90634 80872 90676 80912
rect 90716 80872 90758 80912
rect 90798 80872 90840 80912
rect 90880 80872 105632 80912
rect 105672 80872 105714 80912
rect 105754 80872 105796 80912
rect 105836 80872 105878 80912
rect 105918 80872 105960 80912
rect 106000 80872 120752 80912
rect 120792 80872 120834 80912
rect 120874 80872 120916 80912
rect 120956 80872 120998 80912
rect 121038 80872 121080 80912
rect 121120 80872 135872 80912
rect 135912 80872 135954 80912
rect 135994 80872 136036 80912
rect 136076 80872 136118 80912
rect 136158 80872 136200 80912
rect 136240 80872 150992 80912
rect 151032 80872 151074 80912
rect 151114 80872 151156 80912
rect 151196 80872 151238 80912
rect 151278 80872 151320 80912
rect 151360 80872 152352 80912
rect 71616 80848 152352 80872
rect 71616 80156 152352 80180
rect 71616 80116 74152 80156
rect 74192 80116 74234 80156
rect 74274 80116 74316 80156
rect 74356 80116 74398 80156
rect 74438 80116 74480 80156
rect 74520 80116 89272 80156
rect 89312 80116 89354 80156
rect 89394 80116 89436 80156
rect 89476 80116 89518 80156
rect 89558 80116 89600 80156
rect 89640 80116 104392 80156
rect 104432 80116 104474 80156
rect 104514 80116 104556 80156
rect 104596 80116 104638 80156
rect 104678 80116 104720 80156
rect 104760 80116 119512 80156
rect 119552 80116 119594 80156
rect 119634 80116 119676 80156
rect 119716 80116 119758 80156
rect 119798 80116 119840 80156
rect 119880 80116 134632 80156
rect 134672 80116 134714 80156
rect 134754 80116 134796 80156
rect 134836 80116 134878 80156
rect 134918 80116 134960 80156
rect 135000 80116 149752 80156
rect 149792 80116 149834 80156
rect 149874 80116 149916 80156
rect 149956 80116 149998 80156
rect 150038 80116 150080 80156
rect 150120 80116 152352 80156
rect 71616 80092 152352 80116
rect 71616 79400 152352 79424
rect 71616 79360 75392 79400
rect 75432 79360 75474 79400
rect 75514 79360 75556 79400
rect 75596 79360 75638 79400
rect 75678 79360 75720 79400
rect 75760 79360 90512 79400
rect 90552 79360 90594 79400
rect 90634 79360 90676 79400
rect 90716 79360 90758 79400
rect 90798 79360 90840 79400
rect 90880 79360 105632 79400
rect 105672 79360 105714 79400
rect 105754 79360 105796 79400
rect 105836 79360 105878 79400
rect 105918 79360 105960 79400
rect 106000 79360 120752 79400
rect 120792 79360 120834 79400
rect 120874 79360 120916 79400
rect 120956 79360 120998 79400
rect 121038 79360 121080 79400
rect 121120 79360 135872 79400
rect 135912 79360 135954 79400
rect 135994 79360 136036 79400
rect 136076 79360 136118 79400
rect 136158 79360 136200 79400
rect 136240 79360 150992 79400
rect 151032 79360 151074 79400
rect 151114 79360 151156 79400
rect 151196 79360 151238 79400
rect 151278 79360 151320 79400
rect 151360 79360 152352 79400
rect 71616 79336 152352 79360
rect 71616 78644 152352 78668
rect 71616 78604 74152 78644
rect 74192 78604 74234 78644
rect 74274 78604 74316 78644
rect 74356 78604 74398 78644
rect 74438 78604 74480 78644
rect 74520 78604 89272 78644
rect 89312 78604 89354 78644
rect 89394 78604 89436 78644
rect 89476 78604 89518 78644
rect 89558 78604 89600 78644
rect 89640 78604 104392 78644
rect 104432 78604 104474 78644
rect 104514 78604 104556 78644
rect 104596 78604 104638 78644
rect 104678 78604 104720 78644
rect 104760 78604 119512 78644
rect 119552 78604 119594 78644
rect 119634 78604 119676 78644
rect 119716 78604 119758 78644
rect 119798 78604 119840 78644
rect 119880 78604 134632 78644
rect 134672 78604 134714 78644
rect 134754 78604 134796 78644
rect 134836 78604 134878 78644
rect 134918 78604 134960 78644
rect 135000 78604 149752 78644
rect 149792 78604 149834 78644
rect 149874 78604 149916 78644
rect 149956 78604 149998 78644
rect 150038 78604 150080 78644
rect 150120 78604 152352 78644
rect 71616 78580 152352 78604
rect 71616 77888 152352 77912
rect 71616 77848 75392 77888
rect 75432 77848 75474 77888
rect 75514 77848 75556 77888
rect 75596 77848 75638 77888
rect 75678 77848 75720 77888
rect 75760 77848 90512 77888
rect 90552 77848 90594 77888
rect 90634 77848 90676 77888
rect 90716 77848 90758 77888
rect 90798 77848 90840 77888
rect 90880 77848 105632 77888
rect 105672 77848 105714 77888
rect 105754 77848 105796 77888
rect 105836 77848 105878 77888
rect 105918 77848 105960 77888
rect 106000 77848 120752 77888
rect 120792 77848 120834 77888
rect 120874 77848 120916 77888
rect 120956 77848 120998 77888
rect 121038 77848 121080 77888
rect 121120 77848 135872 77888
rect 135912 77848 135954 77888
rect 135994 77848 136036 77888
rect 136076 77848 136118 77888
rect 136158 77848 136200 77888
rect 136240 77848 150992 77888
rect 151032 77848 151074 77888
rect 151114 77848 151156 77888
rect 151196 77848 151238 77888
rect 151278 77848 151320 77888
rect 151360 77848 152352 77888
rect 71616 77824 152352 77848
rect 71616 77132 152352 77156
rect 71616 77092 74152 77132
rect 74192 77092 74234 77132
rect 74274 77092 74316 77132
rect 74356 77092 74398 77132
rect 74438 77092 74480 77132
rect 74520 77092 89272 77132
rect 89312 77092 89354 77132
rect 89394 77092 89436 77132
rect 89476 77092 89518 77132
rect 89558 77092 89600 77132
rect 89640 77092 104392 77132
rect 104432 77092 104474 77132
rect 104514 77092 104556 77132
rect 104596 77092 104638 77132
rect 104678 77092 104720 77132
rect 104760 77092 119512 77132
rect 119552 77092 119594 77132
rect 119634 77092 119676 77132
rect 119716 77092 119758 77132
rect 119798 77092 119840 77132
rect 119880 77092 134632 77132
rect 134672 77092 134714 77132
rect 134754 77092 134796 77132
rect 134836 77092 134878 77132
rect 134918 77092 134960 77132
rect 135000 77092 149752 77132
rect 149792 77092 149834 77132
rect 149874 77092 149916 77132
rect 149956 77092 149998 77132
rect 150038 77092 150080 77132
rect 150120 77092 152352 77132
rect 71616 77068 152352 77092
rect 71616 76376 152352 76400
rect 71616 76336 75392 76376
rect 75432 76336 75474 76376
rect 75514 76336 75556 76376
rect 75596 76336 75638 76376
rect 75678 76336 75720 76376
rect 75760 76336 90512 76376
rect 90552 76336 90594 76376
rect 90634 76336 90676 76376
rect 90716 76336 90758 76376
rect 90798 76336 90840 76376
rect 90880 76336 105632 76376
rect 105672 76336 105714 76376
rect 105754 76336 105796 76376
rect 105836 76336 105878 76376
rect 105918 76336 105960 76376
rect 106000 76336 120752 76376
rect 120792 76336 120834 76376
rect 120874 76336 120916 76376
rect 120956 76336 120998 76376
rect 121038 76336 121080 76376
rect 121120 76336 135872 76376
rect 135912 76336 135954 76376
rect 135994 76336 136036 76376
rect 136076 76336 136118 76376
rect 136158 76336 136200 76376
rect 136240 76336 150992 76376
rect 151032 76336 151074 76376
rect 151114 76336 151156 76376
rect 151196 76336 151238 76376
rect 151278 76336 151320 76376
rect 151360 76336 152352 76376
rect 71616 76312 152352 76336
rect 71616 75620 152352 75644
rect 71616 75580 74152 75620
rect 74192 75580 74234 75620
rect 74274 75580 74316 75620
rect 74356 75580 74398 75620
rect 74438 75580 74480 75620
rect 74520 75580 89272 75620
rect 89312 75580 89354 75620
rect 89394 75580 89436 75620
rect 89476 75580 89518 75620
rect 89558 75580 89600 75620
rect 89640 75580 104392 75620
rect 104432 75580 104474 75620
rect 104514 75580 104556 75620
rect 104596 75580 104638 75620
rect 104678 75580 104720 75620
rect 104760 75580 119512 75620
rect 119552 75580 119594 75620
rect 119634 75580 119676 75620
rect 119716 75580 119758 75620
rect 119798 75580 119840 75620
rect 119880 75580 134632 75620
rect 134672 75580 134714 75620
rect 134754 75580 134796 75620
rect 134836 75580 134878 75620
rect 134918 75580 134960 75620
rect 135000 75580 149752 75620
rect 149792 75580 149834 75620
rect 149874 75580 149916 75620
rect 149956 75580 149998 75620
rect 150038 75580 150080 75620
rect 150120 75580 152352 75620
rect 71616 75556 152352 75580
rect 71616 74864 152352 74888
rect 71616 74824 75392 74864
rect 75432 74824 75474 74864
rect 75514 74824 75556 74864
rect 75596 74824 75638 74864
rect 75678 74824 75720 74864
rect 75760 74824 90512 74864
rect 90552 74824 90594 74864
rect 90634 74824 90676 74864
rect 90716 74824 90758 74864
rect 90798 74824 90840 74864
rect 90880 74824 105632 74864
rect 105672 74824 105714 74864
rect 105754 74824 105796 74864
rect 105836 74824 105878 74864
rect 105918 74824 105960 74864
rect 106000 74824 120752 74864
rect 120792 74824 120834 74864
rect 120874 74824 120916 74864
rect 120956 74824 120998 74864
rect 121038 74824 121080 74864
rect 121120 74824 135872 74864
rect 135912 74824 135954 74864
rect 135994 74824 136036 74864
rect 136076 74824 136118 74864
rect 136158 74824 136200 74864
rect 136240 74824 150992 74864
rect 151032 74824 151074 74864
rect 151114 74824 151156 74864
rect 151196 74824 151238 74864
rect 151278 74824 151320 74864
rect 151360 74824 152352 74864
rect 71616 74800 152352 74824
rect 71616 74108 152352 74132
rect 71616 74068 74152 74108
rect 74192 74068 74234 74108
rect 74274 74068 74316 74108
rect 74356 74068 74398 74108
rect 74438 74068 74480 74108
rect 74520 74068 89272 74108
rect 89312 74068 89354 74108
rect 89394 74068 89436 74108
rect 89476 74068 89518 74108
rect 89558 74068 89600 74108
rect 89640 74068 104392 74108
rect 104432 74068 104474 74108
rect 104514 74068 104556 74108
rect 104596 74068 104638 74108
rect 104678 74068 104720 74108
rect 104760 74068 119512 74108
rect 119552 74068 119594 74108
rect 119634 74068 119676 74108
rect 119716 74068 119758 74108
rect 119798 74068 119840 74108
rect 119880 74068 134632 74108
rect 134672 74068 134714 74108
rect 134754 74068 134796 74108
rect 134836 74068 134878 74108
rect 134918 74068 134960 74108
rect 135000 74068 149752 74108
rect 149792 74068 149834 74108
rect 149874 74068 149916 74108
rect 149956 74068 149998 74108
rect 150038 74068 150080 74108
rect 150120 74068 152352 74108
rect 71616 74044 152352 74068
rect 71616 73352 152352 73376
rect 71616 73312 75392 73352
rect 75432 73312 75474 73352
rect 75514 73312 75556 73352
rect 75596 73312 75638 73352
rect 75678 73312 75720 73352
rect 75760 73312 90512 73352
rect 90552 73312 90594 73352
rect 90634 73312 90676 73352
rect 90716 73312 90758 73352
rect 90798 73312 90840 73352
rect 90880 73312 105632 73352
rect 105672 73312 105714 73352
rect 105754 73312 105796 73352
rect 105836 73312 105878 73352
rect 105918 73312 105960 73352
rect 106000 73312 120752 73352
rect 120792 73312 120834 73352
rect 120874 73312 120916 73352
rect 120956 73312 120998 73352
rect 121038 73312 121080 73352
rect 121120 73312 135872 73352
rect 135912 73312 135954 73352
rect 135994 73312 136036 73352
rect 136076 73312 136118 73352
rect 136158 73312 136200 73352
rect 136240 73312 150992 73352
rect 151032 73312 151074 73352
rect 151114 73312 151156 73352
rect 151196 73312 151238 73352
rect 151278 73312 151320 73352
rect 151360 73312 152352 73352
rect 71616 73288 152352 73312
rect 71616 72596 152352 72620
rect 71616 72556 74152 72596
rect 74192 72556 74234 72596
rect 74274 72556 74316 72596
rect 74356 72556 74398 72596
rect 74438 72556 74480 72596
rect 74520 72556 89272 72596
rect 89312 72556 89354 72596
rect 89394 72556 89436 72596
rect 89476 72556 89518 72596
rect 89558 72556 89600 72596
rect 89640 72556 104392 72596
rect 104432 72556 104474 72596
rect 104514 72556 104556 72596
rect 104596 72556 104638 72596
rect 104678 72556 104720 72596
rect 104760 72556 119512 72596
rect 119552 72556 119594 72596
rect 119634 72556 119676 72596
rect 119716 72556 119758 72596
rect 119798 72556 119840 72596
rect 119880 72556 134632 72596
rect 134672 72556 134714 72596
rect 134754 72556 134796 72596
rect 134836 72556 134878 72596
rect 134918 72556 134960 72596
rect 135000 72556 149752 72596
rect 149792 72556 149834 72596
rect 149874 72556 149916 72596
rect 149956 72556 149998 72596
rect 150038 72556 150080 72596
rect 150120 72556 152352 72596
rect 71616 72532 152352 72556
rect 71616 71840 152352 71864
rect 71616 71800 75392 71840
rect 75432 71800 75474 71840
rect 75514 71800 75556 71840
rect 75596 71800 75638 71840
rect 75678 71800 75720 71840
rect 75760 71800 90512 71840
rect 90552 71800 90594 71840
rect 90634 71800 90676 71840
rect 90716 71800 90758 71840
rect 90798 71800 90840 71840
rect 90880 71800 105632 71840
rect 105672 71800 105714 71840
rect 105754 71800 105796 71840
rect 105836 71800 105878 71840
rect 105918 71800 105960 71840
rect 106000 71800 120752 71840
rect 120792 71800 120834 71840
rect 120874 71800 120916 71840
rect 120956 71800 120998 71840
rect 121038 71800 121080 71840
rect 121120 71800 135872 71840
rect 135912 71800 135954 71840
rect 135994 71800 136036 71840
rect 136076 71800 136118 71840
rect 136158 71800 136200 71840
rect 136240 71800 150992 71840
rect 151032 71800 151074 71840
rect 151114 71800 151156 71840
rect 151196 71800 151238 71840
rect 151278 71800 151320 71840
rect 151360 71800 152352 71840
rect 71616 71776 152352 71800
<< via1 >>
rect 75392 151936 75432 151976
rect 75474 151936 75514 151976
rect 75556 151936 75596 151976
rect 75638 151936 75678 151976
rect 75720 151936 75760 151976
rect 90512 151936 90552 151976
rect 90594 151936 90634 151976
rect 90676 151936 90716 151976
rect 90758 151936 90798 151976
rect 90840 151936 90880 151976
rect 105632 151936 105672 151976
rect 105714 151936 105754 151976
rect 105796 151936 105836 151976
rect 105878 151936 105918 151976
rect 105960 151936 106000 151976
rect 120752 151936 120792 151976
rect 120834 151936 120874 151976
rect 120916 151936 120956 151976
rect 120998 151936 121038 151976
rect 121080 151936 121120 151976
rect 135872 151936 135912 151976
rect 135954 151936 135994 151976
rect 136036 151936 136076 151976
rect 136118 151936 136158 151976
rect 136200 151936 136240 151976
rect 150992 151936 151032 151976
rect 151074 151936 151114 151976
rect 151156 151936 151196 151976
rect 151238 151936 151278 151976
rect 151320 151936 151360 151976
rect 74152 151180 74192 151220
rect 74234 151180 74274 151220
rect 74316 151180 74356 151220
rect 74398 151180 74438 151220
rect 74480 151180 74520 151220
rect 89272 151180 89312 151220
rect 89354 151180 89394 151220
rect 89436 151180 89476 151220
rect 89518 151180 89558 151220
rect 89600 151180 89640 151220
rect 104392 151180 104432 151220
rect 104474 151180 104514 151220
rect 104556 151180 104596 151220
rect 104638 151180 104678 151220
rect 104720 151180 104760 151220
rect 119512 151180 119552 151220
rect 119594 151180 119634 151220
rect 119676 151180 119716 151220
rect 119758 151180 119798 151220
rect 119840 151180 119880 151220
rect 134632 151180 134672 151220
rect 134714 151180 134754 151220
rect 134796 151180 134836 151220
rect 134878 151180 134918 151220
rect 134960 151180 135000 151220
rect 149752 151180 149792 151220
rect 149834 151180 149874 151220
rect 149916 151180 149956 151220
rect 149998 151180 150038 151220
rect 150080 151180 150120 151220
rect 75392 150424 75432 150464
rect 75474 150424 75514 150464
rect 75556 150424 75596 150464
rect 75638 150424 75678 150464
rect 75720 150424 75760 150464
rect 90512 150424 90552 150464
rect 90594 150424 90634 150464
rect 90676 150424 90716 150464
rect 90758 150424 90798 150464
rect 90840 150424 90880 150464
rect 105632 150424 105672 150464
rect 105714 150424 105754 150464
rect 105796 150424 105836 150464
rect 105878 150424 105918 150464
rect 105960 150424 106000 150464
rect 120752 150424 120792 150464
rect 120834 150424 120874 150464
rect 120916 150424 120956 150464
rect 120998 150424 121038 150464
rect 121080 150424 121120 150464
rect 135872 150424 135912 150464
rect 135954 150424 135994 150464
rect 136036 150424 136076 150464
rect 136118 150424 136158 150464
rect 136200 150424 136240 150464
rect 150992 150424 151032 150464
rect 151074 150424 151114 150464
rect 151156 150424 151196 150464
rect 151238 150424 151278 150464
rect 151320 150424 151360 150464
rect 74152 149668 74192 149708
rect 74234 149668 74274 149708
rect 74316 149668 74356 149708
rect 74398 149668 74438 149708
rect 74480 149668 74520 149708
rect 89272 149668 89312 149708
rect 89354 149668 89394 149708
rect 89436 149668 89476 149708
rect 89518 149668 89558 149708
rect 89600 149668 89640 149708
rect 104392 149668 104432 149708
rect 104474 149668 104514 149708
rect 104556 149668 104596 149708
rect 104638 149668 104678 149708
rect 104720 149668 104760 149708
rect 119512 149668 119552 149708
rect 119594 149668 119634 149708
rect 119676 149668 119716 149708
rect 119758 149668 119798 149708
rect 119840 149668 119880 149708
rect 134632 149668 134672 149708
rect 134714 149668 134754 149708
rect 134796 149668 134836 149708
rect 134878 149668 134918 149708
rect 134960 149668 135000 149708
rect 149752 149668 149792 149708
rect 149834 149668 149874 149708
rect 149916 149668 149956 149708
rect 149998 149668 150038 149708
rect 150080 149668 150120 149708
rect 75392 148912 75432 148952
rect 75474 148912 75514 148952
rect 75556 148912 75596 148952
rect 75638 148912 75678 148952
rect 75720 148912 75760 148952
rect 90512 148912 90552 148952
rect 90594 148912 90634 148952
rect 90676 148912 90716 148952
rect 90758 148912 90798 148952
rect 90840 148912 90880 148952
rect 105632 148912 105672 148952
rect 105714 148912 105754 148952
rect 105796 148912 105836 148952
rect 105878 148912 105918 148952
rect 105960 148912 106000 148952
rect 120752 148912 120792 148952
rect 120834 148912 120874 148952
rect 120916 148912 120956 148952
rect 120998 148912 121038 148952
rect 121080 148912 121120 148952
rect 135872 148912 135912 148952
rect 135954 148912 135994 148952
rect 136036 148912 136076 148952
rect 136118 148912 136158 148952
rect 136200 148912 136240 148952
rect 150992 148912 151032 148952
rect 151074 148912 151114 148952
rect 151156 148912 151196 148952
rect 151238 148912 151278 148952
rect 151320 148912 151360 148952
rect 74152 148156 74192 148196
rect 74234 148156 74274 148196
rect 74316 148156 74356 148196
rect 74398 148156 74438 148196
rect 74480 148156 74520 148196
rect 89272 148156 89312 148196
rect 89354 148156 89394 148196
rect 89436 148156 89476 148196
rect 89518 148156 89558 148196
rect 89600 148156 89640 148196
rect 104392 148156 104432 148196
rect 104474 148156 104514 148196
rect 104556 148156 104596 148196
rect 104638 148156 104678 148196
rect 104720 148156 104760 148196
rect 119512 148156 119552 148196
rect 119594 148156 119634 148196
rect 119676 148156 119716 148196
rect 119758 148156 119798 148196
rect 119840 148156 119880 148196
rect 134632 148156 134672 148196
rect 134714 148156 134754 148196
rect 134796 148156 134836 148196
rect 134878 148156 134918 148196
rect 134960 148156 135000 148196
rect 149752 148156 149792 148196
rect 149834 148156 149874 148196
rect 149916 148156 149956 148196
rect 149998 148156 150038 148196
rect 150080 148156 150120 148196
rect 75392 147400 75432 147440
rect 75474 147400 75514 147440
rect 75556 147400 75596 147440
rect 75638 147400 75678 147440
rect 75720 147400 75760 147440
rect 90512 147400 90552 147440
rect 90594 147400 90634 147440
rect 90676 147400 90716 147440
rect 90758 147400 90798 147440
rect 90840 147400 90880 147440
rect 105632 147400 105672 147440
rect 105714 147400 105754 147440
rect 105796 147400 105836 147440
rect 105878 147400 105918 147440
rect 105960 147400 106000 147440
rect 120752 147400 120792 147440
rect 120834 147400 120874 147440
rect 120916 147400 120956 147440
rect 120998 147400 121038 147440
rect 121080 147400 121120 147440
rect 135872 147400 135912 147440
rect 135954 147400 135994 147440
rect 136036 147400 136076 147440
rect 136118 147400 136158 147440
rect 136200 147400 136240 147440
rect 150992 147400 151032 147440
rect 151074 147400 151114 147440
rect 151156 147400 151196 147440
rect 151238 147400 151278 147440
rect 151320 147400 151360 147440
rect 74152 146644 74192 146684
rect 74234 146644 74274 146684
rect 74316 146644 74356 146684
rect 74398 146644 74438 146684
rect 74480 146644 74520 146684
rect 89272 146644 89312 146684
rect 89354 146644 89394 146684
rect 89436 146644 89476 146684
rect 89518 146644 89558 146684
rect 89600 146644 89640 146684
rect 104392 146644 104432 146684
rect 104474 146644 104514 146684
rect 104556 146644 104596 146684
rect 104638 146644 104678 146684
rect 104720 146644 104760 146684
rect 119512 146644 119552 146684
rect 119594 146644 119634 146684
rect 119676 146644 119716 146684
rect 119758 146644 119798 146684
rect 119840 146644 119880 146684
rect 134632 146644 134672 146684
rect 134714 146644 134754 146684
rect 134796 146644 134836 146684
rect 134878 146644 134918 146684
rect 134960 146644 135000 146684
rect 149752 146644 149792 146684
rect 149834 146644 149874 146684
rect 149916 146644 149956 146684
rect 149998 146644 150038 146684
rect 150080 146644 150120 146684
rect 75392 145888 75432 145928
rect 75474 145888 75514 145928
rect 75556 145888 75596 145928
rect 75638 145888 75678 145928
rect 75720 145888 75760 145928
rect 90512 145888 90552 145928
rect 90594 145888 90634 145928
rect 90676 145888 90716 145928
rect 90758 145888 90798 145928
rect 90840 145888 90880 145928
rect 105632 145888 105672 145928
rect 105714 145888 105754 145928
rect 105796 145888 105836 145928
rect 105878 145888 105918 145928
rect 105960 145888 106000 145928
rect 120752 145888 120792 145928
rect 120834 145888 120874 145928
rect 120916 145888 120956 145928
rect 120998 145888 121038 145928
rect 121080 145888 121120 145928
rect 135872 145888 135912 145928
rect 135954 145888 135994 145928
rect 136036 145888 136076 145928
rect 136118 145888 136158 145928
rect 136200 145888 136240 145928
rect 150992 145888 151032 145928
rect 151074 145888 151114 145928
rect 151156 145888 151196 145928
rect 151238 145888 151278 145928
rect 151320 145888 151360 145928
rect 74152 145132 74192 145172
rect 74234 145132 74274 145172
rect 74316 145132 74356 145172
rect 74398 145132 74438 145172
rect 74480 145132 74520 145172
rect 89272 145132 89312 145172
rect 89354 145132 89394 145172
rect 89436 145132 89476 145172
rect 89518 145132 89558 145172
rect 89600 145132 89640 145172
rect 104392 145132 104432 145172
rect 104474 145132 104514 145172
rect 104556 145132 104596 145172
rect 104638 145132 104678 145172
rect 104720 145132 104760 145172
rect 119512 145132 119552 145172
rect 119594 145132 119634 145172
rect 119676 145132 119716 145172
rect 119758 145132 119798 145172
rect 119840 145132 119880 145172
rect 134632 145132 134672 145172
rect 134714 145132 134754 145172
rect 134796 145132 134836 145172
rect 134878 145132 134918 145172
rect 134960 145132 135000 145172
rect 149752 145132 149792 145172
rect 149834 145132 149874 145172
rect 149916 145132 149956 145172
rect 149998 145132 150038 145172
rect 150080 145132 150120 145172
rect 75392 144376 75432 144416
rect 75474 144376 75514 144416
rect 75556 144376 75596 144416
rect 75638 144376 75678 144416
rect 75720 144376 75760 144416
rect 90512 144376 90552 144416
rect 90594 144376 90634 144416
rect 90676 144376 90716 144416
rect 90758 144376 90798 144416
rect 90840 144376 90880 144416
rect 105632 144376 105672 144416
rect 105714 144376 105754 144416
rect 105796 144376 105836 144416
rect 105878 144376 105918 144416
rect 105960 144376 106000 144416
rect 120752 144376 120792 144416
rect 120834 144376 120874 144416
rect 120916 144376 120956 144416
rect 120998 144376 121038 144416
rect 121080 144376 121120 144416
rect 135872 144376 135912 144416
rect 135954 144376 135994 144416
rect 136036 144376 136076 144416
rect 136118 144376 136158 144416
rect 136200 144376 136240 144416
rect 150992 144376 151032 144416
rect 151074 144376 151114 144416
rect 151156 144376 151196 144416
rect 151238 144376 151278 144416
rect 151320 144376 151360 144416
rect 74152 143620 74192 143660
rect 74234 143620 74274 143660
rect 74316 143620 74356 143660
rect 74398 143620 74438 143660
rect 74480 143620 74520 143660
rect 89272 143620 89312 143660
rect 89354 143620 89394 143660
rect 89436 143620 89476 143660
rect 89518 143620 89558 143660
rect 89600 143620 89640 143660
rect 104392 143620 104432 143660
rect 104474 143620 104514 143660
rect 104556 143620 104596 143660
rect 104638 143620 104678 143660
rect 104720 143620 104760 143660
rect 119512 143620 119552 143660
rect 119594 143620 119634 143660
rect 119676 143620 119716 143660
rect 119758 143620 119798 143660
rect 119840 143620 119880 143660
rect 134632 143620 134672 143660
rect 134714 143620 134754 143660
rect 134796 143620 134836 143660
rect 134878 143620 134918 143660
rect 134960 143620 135000 143660
rect 149752 143620 149792 143660
rect 149834 143620 149874 143660
rect 149916 143620 149956 143660
rect 149998 143620 150038 143660
rect 150080 143620 150120 143660
rect 75392 142864 75432 142904
rect 75474 142864 75514 142904
rect 75556 142864 75596 142904
rect 75638 142864 75678 142904
rect 75720 142864 75760 142904
rect 90512 142864 90552 142904
rect 90594 142864 90634 142904
rect 90676 142864 90716 142904
rect 90758 142864 90798 142904
rect 90840 142864 90880 142904
rect 105632 142864 105672 142904
rect 105714 142864 105754 142904
rect 105796 142864 105836 142904
rect 105878 142864 105918 142904
rect 105960 142864 106000 142904
rect 120752 142864 120792 142904
rect 120834 142864 120874 142904
rect 120916 142864 120956 142904
rect 120998 142864 121038 142904
rect 121080 142864 121120 142904
rect 135872 142864 135912 142904
rect 135954 142864 135994 142904
rect 136036 142864 136076 142904
rect 136118 142864 136158 142904
rect 136200 142864 136240 142904
rect 150992 142864 151032 142904
rect 151074 142864 151114 142904
rect 151156 142864 151196 142904
rect 151238 142864 151278 142904
rect 151320 142864 151360 142904
rect 74152 142108 74192 142148
rect 74234 142108 74274 142148
rect 74316 142108 74356 142148
rect 74398 142108 74438 142148
rect 74480 142108 74520 142148
rect 89272 142108 89312 142148
rect 89354 142108 89394 142148
rect 89436 142108 89476 142148
rect 89518 142108 89558 142148
rect 89600 142108 89640 142148
rect 104392 142108 104432 142148
rect 104474 142108 104514 142148
rect 104556 142108 104596 142148
rect 104638 142108 104678 142148
rect 104720 142108 104760 142148
rect 119512 142108 119552 142148
rect 119594 142108 119634 142148
rect 119676 142108 119716 142148
rect 119758 142108 119798 142148
rect 119840 142108 119880 142148
rect 134632 142108 134672 142148
rect 134714 142108 134754 142148
rect 134796 142108 134836 142148
rect 134878 142108 134918 142148
rect 134960 142108 135000 142148
rect 149752 142108 149792 142148
rect 149834 142108 149874 142148
rect 149916 142108 149956 142148
rect 149998 142108 150038 142148
rect 150080 142108 150120 142148
rect 75392 141352 75432 141392
rect 75474 141352 75514 141392
rect 75556 141352 75596 141392
rect 75638 141352 75678 141392
rect 75720 141352 75760 141392
rect 90512 141352 90552 141392
rect 90594 141352 90634 141392
rect 90676 141352 90716 141392
rect 90758 141352 90798 141392
rect 90840 141352 90880 141392
rect 105632 141352 105672 141392
rect 105714 141352 105754 141392
rect 105796 141352 105836 141392
rect 105878 141352 105918 141392
rect 105960 141352 106000 141392
rect 120752 141352 120792 141392
rect 120834 141352 120874 141392
rect 120916 141352 120956 141392
rect 120998 141352 121038 141392
rect 121080 141352 121120 141392
rect 135872 141352 135912 141392
rect 135954 141352 135994 141392
rect 136036 141352 136076 141392
rect 136118 141352 136158 141392
rect 136200 141352 136240 141392
rect 150992 141352 151032 141392
rect 151074 141352 151114 141392
rect 151156 141352 151196 141392
rect 151238 141352 151278 141392
rect 151320 141352 151360 141392
rect 74152 140596 74192 140636
rect 74234 140596 74274 140636
rect 74316 140596 74356 140636
rect 74398 140596 74438 140636
rect 74480 140596 74520 140636
rect 89272 140596 89312 140636
rect 89354 140596 89394 140636
rect 89436 140596 89476 140636
rect 89518 140596 89558 140636
rect 89600 140596 89640 140636
rect 104392 140596 104432 140636
rect 104474 140596 104514 140636
rect 104556 140596 104596 140636
rect 104638 140596 104678 140636
rect 104720 140596 104760 140636
rect 119512 140596 119552 140636
rect 119594 140596 119634 140636
rect 119676 140596 119716 140636
rect 119758 140596 119798 140636
rect 119840 140596 119880 140636
rect 134632 140596 134672 140636
rect 134714 140596 134754 140636
rect 134796 140596 134836 140636
rect 134878 140596 134918 140636
rect 134960 140596 135000 140636
rect 149752 140596 149792 140636
rect 149834 140596 149874 140636
rect 149916 140596 149956 140636
rect 149998 140596 150038 140636
rect 150080 140596 150120 140636
rect 75392 139840 75432 139880
rect 75474 139840 75514 139880
rect 75556 139840 75596 139880
rect 75638 139840 75678 139880
rect 75720 139840 75760 139880
rect 90512 139840 90552 139880
rect 90594 139840 90634 139880
rect 90676 139840 90716 139880
rect 90758 139840 90798 139880
rect 90840 139840 90880 139880
rect 105632 139840 105672 139880
rect 105714 139840 105754 139880
rect 105796 139840 105836 139880
rect 105878 139840 105918 139880
rect 105960 139840 106000 139880
rect 120752 139840 120792 139880
rect 120834 139840 120874 139880
rect 120916 139840 120956 139880
rect 120998 139840 121038 139880
rect 121080 139840 121120 139880
rect 135872 139840 135912 139880
rect 135954 139840 135994 139880
rect 136036 139840 136076 139880
rect 136118 139840 136158 139880
rect 136200 139840 136240 139880
rect 150992 139840 151032 139880
rect 151074 139840 151114 139880
rect 151156 139840 151196 139880
rect 151238 139840 151278 139880
rect 151320 139840 151360 139880
rect 74152 139084 74192 139124
rect 74234 139084 74274 139124
rect 74316 139084 74356 139124
rect 74398 139084 74438 139124
rect 74480 139084 74520 139124
rect 89272 139084 89312 139124
rect 89354 139084 89394 139124
rect 89436 139084 89476 139124
rect 89518 139084 89558 139124
rect 89600 139084 89640 139124
rect 104392 139084 104432 139124
rect 104474 139084 104514 139124
rect 104556 139084 104596 139124
rect 104638 139084 104678 139124
rect 104720 139084 104760 139124
rect 119512 139084 119552 139124
rect 119594 139084 119634 139124
rect 119676 139084 119716 139124
rect 119758 139084 119798 139124
rect 119840 139084 119880 139124
rect 134632 139084 134672 139124
rect 134714 139084 134754 139124
rect 134796 139084 134836 139124
rect 134878 139084 134918 139124
rect 134960 139084 135000 139124
rect 149752 139084 149792 139124
rect 149834 139084 149874 139124
rect 149916 139084 149956 139124
rect 149998 139084 150038 139124
rect 150080 139084 150120 139124
rect 75392 138328 75432 138368
rect 75474 138328 75514 138368
rect 75556 138328 75596 138368
rect 75638 138328 75678 138368
rect 75720 138328 75760 138368
rect 90512 138328 90552 138368
rect 90594 138328 90634 138368
rect 90676 138328 90716 138368
rect 90758 138328 90798 138368
rect 90840 138328 90880 138368
rect 105632 138328 105672 138368
rect 105714 138328 105754 138368
rect 105796 138328 105836 138368
rect 105878 138328 105918 138368
rect 105960 138328 106000 138368
rect 120752 138328 120792 138368
rect 120834 138328 120874 138368
rect 120916 138328 120956 138368
rect 120998 138328 121038 138368
rect 121080 138328 121120 138368
rect 135872 138328 135912 138368
rect 135954 138328 135994 138368
rect 136036 138328 136076 138368
rect 136118 138328 136158 138368
rect 136200 138328 136240 138368
rect 150992 138328 151032 138368
rect 151074 138328 151114 138368
rect 151156 138328 151196 138368
rect 151238 138328 151278 138368
rect 151320 138328 151360 138368
rect 74152 137572 74192 137612
rect 74234 137572 74274 137612
rect 74316 137572 74356 137612
rect 74398 137572 74438 137612
rect 74480 137572 74520 137612
rect 89272 137572 89312 137612
rect 89354 137572 89394 137612
rect 89436 137572 89476 137612
rect 89518 137572 89558 137612
rect 89600 137572 89640 137612
rect 104392 137572 104432 137612
rect 104474 137572 104514 137612
rect 104556 137572 104596 137612
rect 104638 137572 104678 137612
rect 104720 137572 104760 137612
rect 119512 137572 119552 137612
rect 119594 137572 119634 137612
rect 119676 137572 119716 137612
rect 119758 137572 119798 137612
rect 119840 137572 119880 137612
rect 134632 137572 134672 137612
rect 134714 137572 134754 137612
rect 134796 137572 134836 137612
rect 134878 137572 134918 137612
rect 134960 137572 135000 137612
rect 149752 137572 149792 137612
rect 149834 137572 149874 137612
rect 149916 137572 149956 137612
rect 149998 137572 150038 137612
rect 150080 137572 150120 137612
rect 75392 136816 75432 136856
rect 75474 136816 75514 136856
rect 75556 136816 75596 136856
rect 75638 136816 75678 136856
rect 75720 136816 75760 136856
rect 90512 136816 90552 136856
rect 90594 136816 90634 136856
rect 90676 136816 90716 136856
rect 90758 136816 90798 136856
rect 90840 136816 90880 136856
rect 105632 136816 105672 136856
rect 105714 136816 105754 136856
rect 105796 136816 105836 136856
rect 105878 136816 105918 136856
rect 105960 136816 106000 136856
rect 120752 136816 120792 136856
rect 120834 136816 120874 136856
rect 120916 136816 120956 136856
rect 120998 136816 121038 136856
rect 121080 136816 121120 136856
rect 135872 136816 135912 136856
rect 135954 136816 135994 136856
rect 136036 136816 136076 136856
rect 136118 136816 136158 136856
rect 136200 136816 136240 136856
rect 150992 136816 151032 136856
rect 151074 136816 151114 136856
rect 151156 136816 151196 136856
rect 151238 136816 151278 136856
rect 151320 136816 151360 136856
rect 74152 136060 74192 136100
rect 74234 136060 74274 136100
rect 74316 136060 74356 136100
rect 74398 136060 74438 136100
rect 74480 136060 74520 136100
rect 89272 136060 89312 136100
rect 89354 136060 89394 136100
rect 89436 136060 89476 136100
rect 89518 136060 89558 136100
rect 89600 136060 89640 136100
rect 104392 136060 104432 136100
rect 104474 136060 104514 136100
rect 104556 136060 104596 136100
rect 104638 136060 104678 136100
rect 104720 136060 104760 136100
rect 119512 136060 119552 136100
rect 119594 136060 119634 136100
rect 119676 136060 119716 136100
rect 119758 136060 119798 136100
rect 119840 136060 119880 136100
rect 134632 136060 134672 136100
rect 134714 136060 134754 136100
rect 134796 136060 134836 136100
rect 134878 136060 134918 136100
rect 134960 136060 135000 136100
rect 149752 136060 149792 136100
rect 149834 136060 149874 136100
rect 149916 136060 149956 136100
rect 149998 136060 150038 136100
rect 150080 136060 150120 136100
rect 75392 135304 75432 135344
rect 75474 135304 75514 135344
rect 75556 135304 75596 135344
rect 75638 135304 75678 135344
rect 75720 135304 75760 135344
rect 90512 135304 90552 135344
rect 90594 135304 90634 135344
rect 90676 135304 90716 135344
rect 90758 135304 90798 135344
rect 90840 135304 90880 135344
rect 105632 135304 105672 135344
rect 105714 135304 105754 135344
rect 105796 135304 105836 135344
rect 105878 135304 105918 135344
rect 105960 135304 106000 135344
rect 120752 135304 120792 135344
rect 120834 135304 120874 135344
rect 120916 135304 120956 135344
rect 120998 135304 121038 135344
rect 121080 135304 121120 135344
rect 135872 135304 135912 135344
rect 135954 135304 135994 135344
rect 136036 135304 136076 135344
rect 136118 135304 136158 135344
rect 136200 135304 136240 135344
rect 150992 135304 151032 135344
rect 151074 135304 151114 135344
rect 151156 135304 151196 135344
rect 151238 135304 151278 135344
rect 151320 135304 151360 135344
rect 74152 134548 74192 134588
rect 74234 134548 74274 134588
rect 74316 134548 74356 134588
rect 74398 134548 74438 134588
rect 74480 134548 74520 134588
rect 89272 134548 89312 134588
rect 89354 134548 89394 134588
rect 89436 134548 89476 134588
rect 89518 134548 89558 134588
rect 89600 134548 89640 134588
rect 104392 134548 104432 134588
rect 104474 134548 104514 134588
rect 104556 134548 104596 134588
rect 104638 134548 104678 134588
rect 104720 134548 104760 134588
rect 119512 134548 119552 134588
rect 119594 134548 119634 134588
rect 119676 134548 119716 134588
rect 119758 134548 119798 134588
rect 119840 134548 119880 134588
rect 134632 134548 134672 134588
rect 134714 134548 134754 134588
rect 134796 134548 134836 134588
rect 134878 134548 134918 134588
rect 134960 134548 135000 134588
rect 149752 134548 149792 134588
rect 149834 134548 149874 134588
rect 149916 134548 149956 134588
rect 149998 134548 150038 134588
rect 150080 134548 150120 134588
rect 75392 133792 75432 133832
rect 75474 133792 75514 133832
rect 75556 133792 75596 133832
rect 75638 133792 75678 133832
rect 75720 133792 75760 133832
rect 90512 133792 90552 133832
rect 90594 133792 90634 133832
rect 90676 133792 90716 133832
rect 90758 133792 90798 133832
rect 90840 133792 90880 133832
rect 105632 133792 105672 133832
rect 105714 133792 105754 133832
rect 105796 133792 105836 133832
rect 105878 133792 105918 133832
rect 105960 133792 106000 133832
rect 120752 133792 120792 133832
rect 120834 133792 120874 133832
rect 120916 133792 120956 133832
rect 120998 133792 121038 133832
rect 121080 133792 121120 133832
rect 135872 133792 135912 133832
rect 135954 133792 135994 133832
rect 136036 133792 136076 133832
rect 136118 133792 136158 133832
rect 136200 133792 136240 133832
rect 150992 133792 151032 133832
rect 151074 133792 151114 133832
rect 151156 133792 151196 133832
rect 151238 133792 151278 133832
rect 151320 133792 151360 133832
rect 74152 133036 74192 133076
rect 74234 133036 74274 133076
rect 74316 133036 74356 133076
rect 74398 133036 74438 133076
rect 74480 133036 74520 133076
rect 89272 133036 89312 133076
rect 89354 133036 89394 133076
rect 89436 133036 89476 133076
rect 89518 133036 89558 133076
rect 89600 133036 89640 133076
rect 104392 133036 104432 133076
rect 104474 133036 104514 133076
rect 104556 133036 104596 133076
rect 104638 133036 104678 133076
rect 104720 133036 104760 133076
rect 119512 133036 119552 133076
rect 119594 133036 119634 133076
rect 119676 133036 119716 133076
rect 119758 133036 119798 133076
rect 119840 133036 119880 133076
rect 134632 133036 134672 133076
rect 134714 133036 134754 133076
rect 134796 133036 134836 133076
rect 134878 133036 134918 133076
rect 134960 133036 135000 133076
rect 149752 133036 149792 133076
rect 149834 133036 149874 133076
rect 149916 133036 149956 133076
rect 149998 133036 150038 133076
rect 150080 133036 150120 133076
rect 75392 132280 75432 132320
rect 75474 132280 75514 132320
rect 75556 132280 75596 132320
rect 75638 132280 75678 132320
rect 75720 132280 75760 132320
rect 90512 132280 90552 132320
rect 90594 132280 90634 132320
rect 90676 132280 90716 132320
rect 90758 132280 90798 132320
rect 90840 132280 90880 132320
rect 105632 132280 105672 132320
rect 105714 132280 105754 132320
rect 105796 132280 105836 132320
rect 105878 132280 105918 132320
rect 105960 132280 106000 132320
rect 120752 132280 120792 132320
rect 120834 132280 120874 132320
rect 120916 132280 120956 132320
rect 120998 132280 121038 132320
rect 121080 132280 121120 132320
rect 135872 132280 135912 132320
rect 135954 132280 135994 132320
rect 136036 132280 136076 132320
rect 136118 132280 136158 132320
rect 136200 132280 136240 132320
rect 150992 132280 151032 132320
rect 151074 132280 151114 132320
rect 151156 132280 151196 132320
rect 151238 132280 151278 132320
rect 151320 132280 151360 132320
rect 74152 131524 74192 131564
rect 74234 131524 74274 131564
rect 74316 131524 74356 131564
rect 74398 131524 74438 131564
rect 74480 131524 74520 131564
rect 89272 131524 89312 131564
rect 89354 131524 89394 131564
rect 89436 131524 89476 131564
rect 89518 131524 89558 131564
rect 89600 131524 89640 131564
rect 104392 131524 104432 131564
rect 104474 131524 104514 131564
rect 104556 131524 104596 131564
rect 104638 131524 104678 131564
rect 104720 131524 104760 131564
rect 119512 131524 119552 131564
rect 119594 131524 119634 131564
rect 119676 131524 119716 131564
rect 119758 131524 119798 131564
rect 119840 131524 119880 131564
rect 134632 131524 134672 131564
rect 134714 131524 134754 131564
rect 134796 131524 134836 131564
rect 134878 131524 134918 131564
rect 134960 131524 135000 131564
rect 149752 131524 149792 131564
rect 149834 131524 149874 131564
rect 149916 131524 149956 131564
rect 149998 131524 150038 131564
rect 150080 131524 150120 131564
rect 75392 130768 75432 130808
rect 75474 130768 75514 130808
rect 75556 130768 75596 130808
rect 75638 130768 75678 130808
rect 75720 130768 75760 130808
rect 90512 130768 90552 130808
rect 90594 130768 90634 130808
rect 90676 130768 90716 130808
rect 90758 130768 90798 130808
rect 90840 130768 90880 130808
rect 105632 130768 105672 130808
rect 105714 130768 105754 130808
rect 105796 130768 105836 130808
rect 105878 130768 105918 130808
rect 105960 130768 106000 130808
rect 120752 130768 120792 130808
rect 120834 130768 120874 130808
rect 120916 130768 120956 130808
rect 120998 130768 121038 130808
rect 121080 130768 121120 130808
rect 135872 130768 135912 130808
rect 135954 130768 135994 130808
rect 136036 130768 136076 130808
rect 136118 130768 136158 130808
rect 136200 130768 136240 130808
rect 150992 130768 151032 130808
rect 151074 130768 151114 130808
rect 151156 130768 151196 130808
rect 151238 130768 151278 130808
rect 151320 130768 151360 130808
rect 74152 130012 74192 130052
rect 74234 130012 74274 130052
rect 74316 130012 74356 130052
rect 74398 130012 74438 130052
rect 74480 130012 74520 130052
rect 89272 130012 89312 130052
rect 89354 130012 89394 130052
rect 89436 130012 89476 130052
rect 89518 130012 89558 130052
rect 89600 130012 89640 130052
rect 104392 130012 104432 130052
rect 104474 130012 104514 130052
rect 104556 130012 104596 130052
rect 104638 130012 104678 130052
rect 104720 130012 104760 130052
rect 119512 130012 119552 130052
rect 119594 130012 119634 130052
rect 119676 130012 119716 130052
rect 119758 130012 119798 130052
rect 119840 130012 119880 130052
rect 134632 130012 134672 130052
rect 134714 130012 134754 130052
rect 134796 130012 134836 130052
rect 134878 130012 134918 130052
rect 134960 130012 135000 130052
rect 149752 130012 149792 130052
rect 149834 130012 149874 130052
rect 149916 130012 149956 130052
rect 149998 130012 150038 130052
rect 150080 130012 150120 130052
rect 75392 129256 75432 129296
rect 75474 129256 75514 129296
rect 75556 129256 75596 129296
rect 75638 129256 75678 129296
rect 75720 129256 75760 129296
rect 90512 129256 90552 129296
rect 90594 129256 90634 129296
rect 90676 129256 90716 129296
rect 90758 129256 90798 129296
rect 90840 129256 90880 129296
rect 105632 129256 105672 129296
rect 105714 129256 105754 129296
rect 105796 129256 105836 129296
rect 105878 129256 105918 129296
rect 105960 129256 106000 129296
rect 120752 129256 120792 129296
rect 120834 129256 120874 129296
rect 120916 129256 120956 129296
rect 120998 129256 121038 129296
rect 121080 129256 121120 129296
rect 135872 129256 135912 129296
rect 135954 129256 135994 129296
rect 136036 129256 136076 129296
rect 136118 129256 136158 129296
rect 136200 129256 136240 129296
rect 150992 129256 151032 129296
rect 151074 129256 151114 129296
rect 151156 129256 151196 129296
rect 151238 129256 151278 129296
rect 151320 129256 151360 129296
rect 74152 128500 74192 128540
rect 74234 128500 74274 128540
rect 74316 128500 74356 128540
rect 74398 128500 74438 128540
rect 74480 128500 74520 128540
rect 89272 128500 89312 128540
rect 89354 128500 89394 128540
rect 89436 128500 89476 128540
rect 89518 128500 89558 128540
rect 89600 128500 89640 128540
rect 104392 128500 104432 128540
rect 104474 128500 104514 128540
rect 104556 128500 104596 128540
rect 104638 128500 104678 128540
rect 104720 128500 104760 128540
rect 119512 128500 119552 128540
rect 119594 128500 119634 128540
rect 119676 128500 119716 128540
rect 119758 128500 119798 128540
rect 119840 128500 119880 128540
rect 134632 128500 134672 128540
rect 134714 128500 134754 128540
rect 134796 128500 134836 128540
rect 134878 128500 134918 128540
rect 134960 128500 135000 128540
rect 149752 128500 149792 128540
rect 149834 128500 149874 128540
rect 149916 128500 149956 128540
rect 149998 128500 150038 128540
rect 150080 128500 150120 128540
rect 75392 127744 75432 127784
rect 75474 127744 75514 127784
rect 75556 127744 75596 127784
rect 75638 127744 75678 127784
rect 75720 127744 75760 127784
rect 90512 127744 90552 127784
rect 90594 127744 90634 127784
rect 90676 127744 90716 127784
rect 90758 127744 90798 127784
rect 90840 127744 90880 127784
rect 105632 127744 105672 127784
rect 105714 127744 105754 127784
rect 105796 127744 105836 127784
rect 105878 127744 105918 127784
rect 105960 127744 106000 127784
rect 120752 127744 120792 127784
rect 120834 127744 120874 127784
rect 120916 127744 120956 127784
rect 120998 127744 121038 127784
rect 121080 127744 121120 127784
rect 135872 127744 135912 127784
rect 135954 127744 135994 127784
rect 136036 127744 136076 127784
rect 136118 127744 136158 127784
rect 136200 127744 136240 127784
rect 150992 127744 151032 127784
rect 151074 127744 151114 127784
rect 151156 127744 151196 127784
rect 151238 127744 151278 127784
rect 151320 127744 151360 127784
rect 74152 126988 74192 127028
rect 74234 126988 74274 127028
rect 74316 126988 74356 127028
rect 74398 126988 74438 127028
rect 74480 126988 74520 127028
rect 89272 126988 89312 127028
rect 89354 126988 89394 127028
rect 89436 126988 89476 127028
rect 89518 126988 89558 127028
rect 89600 126988 89640 127028
rect 104392 126988 104432 127028
rect 104474 126988 104514 127028
rect 104556 126988 104596 127028
rect 104638 126988 104678 127028
rect 104720 126988 104760 127028
rect 119512 126988 119552 127028
rect 119594 126988 119634 127028
rect 119676 126988 119716 127028
rect 119758 126988 119798 127028
rect 119840 126988 119880 127028
rect 134632 126988 134672 127028
rect 134714 126988 134754 127028
rect 134796 126988 134836 127028
rect 134878 126988 134918 127028
rect 134960 126988 135000 127028
rect 149752 126988 149792 127028
rect 149834 126988 149874 127028
rect 149916 126988 149956 127028
rect 149998 126988 150038 127028
rect 150080 126988 150120 127028
rect 75392 126232 75432 126272
rect 75474 126232 75514 126272
rect 75556 126232 75596 126272
rect 75638 126232 75678 126272
rect 75720 126232 75760 126272
rect 90512 126232 90552 126272
rect 90594 126232 90634 126272
rect 90676 126232 90716 126272
rect 90758 126232 90798 126272
rect 90840 126232 90880 126272
rect 105632 126232 105672 126272
rect 105714 126232 105754 126272
rect 105796 126232 105836 126272
rect 105878 126232 105918 126272
rect 105960 126232 106000 126272
rect 120752 126232 120792 126272
rect 120834 126232 120874 126272
rect 120916 126232 120956 126272
rect 120998 126232 121038 126272
rect 121080 126232 121120 126272
rect 135872 126232 135912 126272
rect 135954 126232 135994 126272
rect 136036 126232 136076 126272
rect 136118 126232 136158 126272
rect 136200 126232 136240 126272
rect 150992 126232 151032 126272
rect 151074 126232 151114 126272
rect 151156 126232 151196 126272
rect 151238 126232 151278 126272
rect 151320 126232 151360 126272
rect 74152 125476 74192 125516
rect 74234 125476 74274 125516
rect 74316 125476 74356 125516
rect 74398 125476 74438 125516
rect 74480 125476 74520 125516
rect 89272 125476 89312 125516
rect 89354 125476 89394 125516
rect 89436 125476 89476 125516
rect 89518 125476 89558 125516
rect 89600 125476 89640 125516
rect 104392 125476 104432 125516
rect 104474 125476 104514 125516
rect 104556 125476 104596 125516
rect 104638 125476 104678 125516
rect 104720 125476 104760 125516
rect 119512 125476 119552 125516
rect 119594 125476 119634 125516
rect 119676 125476 119716 125516
rect 119758 125476 119798 125516
rect 119840 125476 119880 125516
rect 134632 125476 134672 125516
rect 134714 125476 134754 125516
rect 134796 125476 134836 125516
rect 134878 125476 134918 125516
rect 134960 125476 135000 125516
rect 149752 125476 149792 125516
rect 149834 125476 149874 125516
rect 149916 125476 149956 125516
rect 149998 125476 150038 125516
rect 150080 125476 150120 125516
rect 75392 124720 75432 124760
rect 75474 124720 75514 124760
rect 75556 124720 75596 124760
rect 75638 124720 75678 124760
rect 75720 124720 75760 124760
rect 90512 124720 90552 124760
rect 90594 124720 90634 124760
rect 90676 124720 90716 124760
rect 90758 124720 90798 124760
rect 90840 124720 90880 124760
rect 105632 124720 105672 124760
rect 105714 124720 105754 124760
rect 105796 124720 105836 124760
rect 105878 124720 105918 124760
rect 105960 124720 106000 124760
rect 120752 124720 120792 124760
rect 120834 124720 120874 124760
rect 120916 124720 120956 124760
rect 120998 124720 121038 124760
rect 121080 124720 121120 124760
rect 135872 124720 135912 124760
rect 135954 124720 135994 124760
rect 136036 124720 136076 124760
rect 136118 124720 136158 124760
rect 136200 124720 136240 124760
rect 150992 124720 151032 124760
rect 151074 124720 151114 124760
rect 151156 124720 151196 124760
rect 151238 124720 151278 124760
rect 151320 124720 151360 124760
rect 74152 123964 74192 124004
rect 74234 123964 74274 124004
rect 74316 123964 74356 124004
rect 74398 123964 74438 124004
rect 74480 123964 74520 124004
rect 89272 123964 89312 124004
rect 89354 123964 89394 124004
rect 89436 123964 89476 124004
rect 89518 123964 89558 124004
rect 89600 123964 89640 124004
rect 104392 123964 104432 124004
rect 104474 123964 104514 124004
rect 104556 123964 104596 124004
rect 104638 123964 104678 124004
rect 104720 123964 104760 124004
rect 119512 123964 119552 124004
rect 119594 123964 119634 124004
rect 119676 123964 119716 124004
rect 119758 123964 119798 124004
rect 119840 123964 119880 124004
rect 134632 123964 134672 124004
rect 134714 123964 134754 124004
rect 134796 123964 134836 124004
rect 134878 123964 134918 124004
rect 134960 123964 135000 124004
rect 149752 123964 149792 124004
rect 149834 123964 149874 124004
rect 149916 123964 149956 124004
rect 149998 123964 150038 124004
rect 150080 123964 150120 124004
rect 75392 123208 75432 123248
rect 75474 123208 75514 123248
rect 75556 123208 75596 123248
rect 75638 123208 75678 123248
rect 75720 123208 75760 123248
rect 90512 123208 90552 123248
rect 90594 123208 90634 123248
rect 90676 123208 90716 123248
rect 90758 123208 90798 123248
rect 90840 123208 90880 123248
rect 105632 123208 105672 123248
rect 105714 123208 105754 123248
rect 105796 123208 105836 123248
rect 105878 123208 105918 123248
rect 105960 123208 106000 123248
rect 120752 123208 120792 123248
rect 120834 123208 120874 123248
rect 120916 123208 120956 123248
rect 120998 123208 121038 123248
rect 121080 123208 121120 123248
rect 135872 123208 135912 123248
rect 135954 123208 135994 123248
rect 136036 123208 136076 123248
rect 136118 123208 136158 123248
rect 136200 123208 136240 123248
rect 150992 123208 151032 123248
rect 151074 123208 151114 123248
rect 151156 123208 151196 123248
rect 151238 123208 151278 123248
rect 151320 123208 151360 123248
rect 74152 122452 74192 122492
rect 74234 122452 74274 122492
rect 74316 122452 74356 122492
rect 74398 122452 74438 122492
rect 74480 122452 74520 122492
rect 89272 122452 89312 122492
rect 89354 122452 89394 122492
rect 89436 122452 89476 122492
rect 89518 122452 89558 122492
rect 89600 122452 89640 122492
rect 104392 122452 104432 122492
rect 104474 122452 104514 122492
rect 104556 122452 104596 122492
rect 104638 122452 104678 122492
rect 104720 122452 104760 122492
rect 119512 122452 119552 122492
rect 119594 122452 119634 122492
rect 119676 122452 119716 122492
rect 119758 122452 119798 122492
rect 119840 122452 119880 122492
rect 134632 122452 134672 122492
rect 134714 122452 134754 122492
rect 134796 122452 134836 122492
rect 134878 122452 134918 122492
rect 134960 122452 135000 122492
rect 149752 122452 149792 122492
rect 149834 122452 149874 122492
rect 149916 122452 149956 122492
rect 149998 122452 150038 122492
rect 150080 122452 150120 122492
rect 75392 121696 75432 121736
rect 75474 121696 75514 121736
rect 75556 121696 75596 121736
rect 75638 121696 75678 121736
rect 75720 121696 75760 121736
rect 90512 121696 90552 121736
rect 90594 121696 90634 121736
rect 90676 121696 90716 121736
rect 90758 121696 90798 121736
rect 90840 121696 90880 121736
rect 105632 121696 105672 121736
rect 105714 121696 105754 121736
rect 105796 121696 105836 121736
rect 105878 121696 105918 121736
rect 105960 121696 106000 121736
rect 120752 121696 120792 121736
rect 120834 121696 120874 121736
rect 120916 121696 120956 121736
rect 120998 121696 121038 121736
rect 121080 121696 121120 121736
rect 135872 121696 135912 121736
rect 135954 121696 135994 121736
rect 136036 121696 136076 121736
rect 136118 121696 136158 121736
rect 136200 121696 136240 121736
rect 150992 121696 151032 121736
rect 151074 121696 151114 121736
rect 151156 121696 151196 121736
rect 151238 121696 151278 121736
rect 151320 121696 151360 121736
rect 74152 120940 74192 120980
rect 74234 120940 74274 120980
rect 74316 120940 74356 120980
rect 74398 120940 74438 120980
rect 74480 120940 74520 120980
rect 89272 120940 89312 120980
rect 89354 120940 89394 120980
rect 89436 120940 89476 120980
rect 89518 120940 89558 120980
rect 89600 120940 89640 120980
rect 104392 120940 104432 120980
rect 104474 120940 104514 120980
rect 104556 120940 104596 120980
rect 104638 120940 104678 120980
rect 104720 120940 104760 120980
rect 119512 120940 119552 120980
rect 119594 120940 119634 120980
rect 119676 120940 119716 120980
rect 119758 120940 119798 120980
rect 119840 120940 119880 120980
rect 134632 120940 134672 120980
rect 134714 120940 134754 120980
rect 134796 120940 134836 120980
rect 134878 120940 134918 120980
rect 134960 120940 135000 120980
rect 149752 120940 149792 120980
rect 149834 120940 149874 120980
rect 149916 120940 149956 120980
rect 149998 120940 150038 120980
rect 150080 120940 150120 120980
rect 75392 120184 75432 120224
rect 75474 120184 75514 120224
rect 75556 120184 75596 120224
rect 75638 120184 75678 120224
rect 75720 120184 75760 120224
rect 90512 120184 90552 120224
rect 90594 120184 90634 120224
rect 90676 120184 90716 120224
rect 90758 120184 90798 120224
rect 90840 120184 90880 120224
rect 105632 120184 105672 120224
rect 105714 120184 105754 120224
rect 105796 120184 105836 120224
rect 105878 120184 105918 120224
rect 105960 120184 106000 120224
rect 120752 120184 120792 120224
rect 120834 120184 120874 120224
rect 120916 120184 120956 120224
rect 120998 120184 121038 120224
rect 121080 120184 121120 120224
rect 135872 120184 135912 120224
rect 135954 120184 135994 120224
rect 136036 120184 136076 120224
rect 136118 120184 136158 120224
rect 136200 120184 136240 120224
rect 150992 120184 151032 120224
rect 151074 120184 151114 120224
rect 151156 120184 151196 120224
rect 151238 120184 151278 120224
rect 151320 120184 151360 120224
rect 74152 119428 74192 119468
rect 74234 119428 74274 119468
rect 74316 119428 74356 119468
rect 74398 119428 74438 119468
rect 74480 119428 74520 119468
rect 89272 119428 89312 119468
rect 89354 119428 89394 119468
rect 89436 119428 89476 119468
rect 89518 119428 89558 119468
rect 89600 119428 89640 119468
rect 104392 119428 104432 119468
rect 104474 119428 104514 119468
rect 104556 119428 104596 119468
rect 104638 119428 104678 119468
rect 104720 119428 104760 119468
rect 119512 119428 119552 119468
rect 119594 119428 119634 119468
rect 119676 119428 119716 119468
rect 119758 119428 119798 119468
rect 119840 119428 119880 119468
rect 134632 119428 134672 119468
rect 134714 119428 134754 119468
rect 134796 119428 134836 119468
rect 134878 119428 134918 119468
rect 134960 119428 135000 119468
rect 149752 119428 149792 119468
rect 149834 119428 149874 119468
rect 149916 119428 149956 119468
rect 149998 119428 150038 119468
rect 150080 119428 150120 119468
rect 75392 118672 75432 118712
rect 75474 118672 75514 118712
rect 75556 118672 75596 118712
rect 75638 118672 75678 118712
rect 75720 118672 75760 118712
rect 90512 118672 90552 118712
rect 90594 118672 90634 118712
rect 90676 118672 90716 118712
rect 90758 118672 90798 118712
rect 90840 118672 90880 118712
rect 105632 118672 105672 118712
rect 105714 118672 105754 118712
rect 105796 118672 105836 118712
rect 105878 118672 105918 118712
rect 105960 118672 106000 118712
rect 120752 118672 120792 118712
rect 120834 118672 120874 118712
rect 120916 118672 120956 118712
rect 120998 118672 121038 118712
rect 121080 118672 121120 118712
rect 135872 118672 135912 118712
rect 135954 118672 135994 118712
rect 136036 118672 136076 118712
rect 136118 118672 136158 118712
rect 136200 118672 136240 118712
rect 150992 118672 151032 118712
rect 151074 118672 151114 118712
rect 151156 118672 151196 118712
rect 151238 118672 151278 118712
rect 151320 118672 151360 118712
rect 74152 117916 74192 117956
rect 74234 117916 74274 117956
rect 74316 117916 74356 117956
rect 74398 117916 74438 117956
rect 74480 117916 74520 117956
rect 89272 117916 89312 117956
rect 89354 117916 89394 117956
rect 89436 117916 89476 117956
rect 89518 117916 89558 117956
rect 89600 117916 89640 117956
rect 104392 117916 104432 117956
rect 104474 117916 104514 117956
rect 104556 117916 104596 117956
rect 104638 117916 104678 117956
rect 104720 117916 104760 117956
rect 119512 117916 119552 117956
rect 119594 117916 119634 117956
rect 119676 117916 119716 117956
rect 119758 117916 119798 117956
rect 119840 117916 119880 117956
rect 134632 117916 134672 117956
rect 134714 117916 134754 117956
rect 134796 117916 134836 117956
rect 134878 117916 134918 117956
rect 134960 117916 135000 117956
rect 149752 117916 149792 117956
rect 149834 117916 149874 117956
rect 149916 117916 149956 117956
rect 149998 117916 150038 117956
rect 150080 117916 150120 117956
rect 75392 117160 75432 117200
rect 75474 117160 75514 117200
rect 75556 117160 75596 117200
rect 75638 117160 75678 117200
rect 75720 117160 75760 117200
rect 90512 117160 90552 117200
rect 90594 117160 90634 117200
rect 90676 117160 90716 117200
rect 90758 117160 90798 117200
rect 90840 117160 90880 117200
rect 105632 117160 105672 117200
rect 105714 117160 105754 117200
rect 105796 117160 105836 117200
rect 105878 117160 105918 117200
rect 105960 117160 106000 117200
rect 120752 117160 120792 117200
rect 120834 117160 120874 117200
rect 120916 117160 120956 117200
rect 120998 117160 121038 117200
rect 121080 117160 121120 117200
rect 135872 117160 135912 117200
rect 135954 117160 135994 117200
rect 136036 117160 136076 117200
rect 136118 117160 136158 117200
rect 136200 117160 136240 117200
rect 150992 117160 151032 117200
rect 151074 117160 151114 117200
rect 151156 117160 151196 117200
rect 151238 117160 151278 117200
rect 151320 117160 151360 117200
rect 74152 116404 74192 116444
rect 74234 116404 74274 116444
rect 74316 116404 74356 116444
rect 74398 116404 74438 116444
rect 74480 116404 74520 116444
rect 89272 116404 89312 116444
rect 89354 116404 89394 116444
rect 89436 116404 89476 116444
rect 89518 116404 89558 116444
rect 89600 116404 89640 116444
rect 104392 116404 104432 116444
rect 104474 116404 104514 116444
rect 104556 116404 104596 116444
rect 104638 116404 104678 116444
rect 104720 116404 104760 116444
rect 119512 116404 119552 116444
rect 119594 116404 119634 116444
rect 119676 116404 119716 116444
rect 119758 116404 119798 116444
rect 119840 116404 119880 116444
rect 134632 116404 134672 116444
rect 134714 116404 134754 116444
rect 134796 116404 134836 116444
rect 134878 116404 134918 116444
rect 134960 116404 135000 116444
rect 149752 116404 149792 116444
rect 149834 116404 149874 116444
rect 149916 116404 149956 116444
rect 149998 116404 150038 116444
rect 150080 116404 150120 116444
rect 75392 115648 75432 115688
rect 75474 115648 75514 115688
rect 75556 115648 75596 115688
rect 75638 115648 75678 115688
rect 75720 115648 75760 115688
rect 90512 115648 90552 115688
rect 90594 115648 90634 115688
rect 90676 115648 90716 115688
rect 90758 115648 90798 115688
rect 90840 115648 90880 115688
rect 105632 115648 105672 115688
rect 105714 115648 105754 115688
rect 105796 115648 105836 115688
rect 105878 115648 105918 115688
rect 105960 115648 106000 115688
rect 120752 115648 120792 115688
rect 120834 115648 120874 115688
rect 120916 115648 120956 115688
rect 120998 115648 121038 115688
rect 121080 115648 121120 115688
rect 135872 115648 135912 115688
rect 135954 115648 135994 115688
rect 136036 115648 136076 115688
rect 136118 115648 136158 115688
rect 136200 115648 136240 115688
rect 150992 115648 151032 115688
rect 151074 115648 151114 115688
rect 151156 115648 151196 115688
rect 151238 115648 151278 115688
rect 151320 115648 151360 115688
rect 74152 114892 74192 114932
rect 74234 114892 74274 114932
rect 74316 114892 74356 114932
rect 74398 114892 74438 114932
rect 74480 114892 74520 114932
rect 89272 114892 89312 114932
rect 89354 114892 89394 114932
rect 89436 114892 89476 114932
rect 89518 114892 89558 114932
rect 89600 114892 89640 114932
rect 104392 114892 104432 114932
rect 104474 114892 104514 114932
rect 104556 114892 104596 114932
rect 104638 114892 104678 114932
rect 104720 114892 104760 114932
rect 119512 114892 119552 114932
rect 119594 114892 119634 114932
rect 119676 114892 119716 114932
rect 119758 114892 119798 114932
rect 119840 114892 119880 114932
rect 134632 114892 134672 114932
rect 134714 114892 134754 114932
rect 134796 114892 134836 114932
rect 134878 114892 134918 114932
rect 134960 114892 135000 114932
rect 149752 114892 149792 114932
rect 149834 114892 149874 114932
rect 149916 114892 149956 114932
rect 149998 114892 150038 114932
rect 150080 114892 150120 114932
rect 75392 114136 75432 114176
rect 75474 114136 75514 114176
rect 75556 114136 75596 114176
rect 75638 114136 75678 114176
rect 75720 114136 75760 114176
rect 90512 114136 90552 114176
rect 90594 114136 90634 114176
rect 90676 114136 90716 114176
rect 90758 114136 90798 114176
rect 90840 114136 90880 114176
rect 105632 114136 105672 114176
rect 105714 114136 105754 114176
rect 105796 114136 105836 114176
rect 105878 114136 105918 114176
rect 105960 114136 106000 114176
rect 120752 114136 120792 114176
rect 120834 114136 120874 114176
rect 120916 114136 120956 114176
rect 120998 114136 121038 114176
rect 121080 114136 121120 114176
rect 135872 114136 135912 114176
rect 135954 114136 135994 114176
rect 136036 114136 136076 114176
rect 136118 114136 136158 114176
rect 136200 114136 136240 114176
rect 150992 114136 151032 114176
rect 151074 114136 151114 114176
rect 151156 114136 151196 114176
rect 151238 114136 151278 114176
rect 151320 114136 151360 114176
rect 74152 113380 74192 113420
rect 74234 113380 74274 113420
rect 74316 113380 74356 113420
rect 74398 113380 74438 113420
rect 74480 113380 74520 113420
rect 89272 113380 89312 113420
rect 89354 113380 89394 113420
rect 89436 113380 89476 113420
rect 89518 113380 89558 113420
rect 89600 113380 89640 113420
rect 104392 113380 104432 113420
rect 104474 113380 104514 113420
rect 104556 113380 104596 113420
rect 104638 113380 104678 113420
rect 104720 113380 104760 113420
rect 119512 113380 119552 113420
rect 119594 113380 119634 113420
rect 119676 113380 119716 113420
rect 119758 113380 119798 113420
rect 119840 113380 119880 113420
rect 134632 113380 134672 113420
rect 134714 113380 134754 113420
rect 134796 113380 134836 113420
rect 134878 113380 134918 113420
rect 134960 113380 135000 113420
rect 149752 113380 149792 113420
rect 149834 113380 149874 113420
rect 149916 113380 149956 113420
rect 149998 113380 150038 113420
rect 150080 113380 150120 113420
rect 75392 112624 75432 112664
rect 75474 112624 75514 112664
rect 75556 112624 75596 112664
rect 75638 112624 75678 112664
rect 75720 112624 75760 112664
rect 90512 112624 90552 112664
rect 90594 112624 90634 112664
rect 90676 112624 90716 112664
rect 90758 112624 90798 112664
rect 90840 112624 90880 112664
rect 105632 112624 105672 112664
rect 105714 112624 105754 112664
rect 105796 112624 105836 112664
rect 105878 112624 105918 112664
rect 105960 112624 106000 112664
rect 120752 112624 120792 112664
rect 120834 112624 120874 112664
rect 120916 112624 120956 112664
rect 120998 112624 121038 112664
rect 121080 112624 121120 112664
rect 135872 112624 135912 112664
rect 135954 112624 135994 112664
rect 136036 112624 136076 112664
rect 136118 112624 136158 112664
rect 136200 112624 136240 112664
rect 150992 112624 151032 112664
rect 151074 112624 151114 112664
rect 151156 112624 151196 112664
rect 151238 112624 151278 112664
rect 151320 112624 151360 112664
rect 74152 111868 74192 111908
rect 74234 111868 74274 111908
rect 74316 111868 74356 111908
rect 74398 111868 74438 111908
rect 74480 111868 74520 111908
rect 89272 111868 89312 111908
rect 89354 111868 89394 111908
rect 89436 111868 89476 111908
rect 89518 111868 89558 111908
rect 89600 111868 89640 111908
rect 104392 111868 104432 111908
rect 104474 111868 104514 111908
rect 104556 111868 104596 111908
rect 104638 111868 104678 111908
rect 104720 111868 104760 111908
rect 119512 111868 119552 111908
rect 119594 111868 119634 111908
rect 119676 111868 119716 111908
rect 119758 111868 119798 111908
rect 119840 111868 119880 111908
rect 134632 111868 134672 111908
rect 134714 111868 134754 111908
rect 134796 111868 134836 111908
rect 134878 111868 134918 111908
rect 134960 111868 135000 111908
rect 149752 111868 149792 111908
rect 149834 111868 149874 111908
rect 149916 111868 149956 111908
rect 149998 111868 150038 111908
rect 150080 111868 150120 111908
rect 75392 111112 75432 111152
rect 75474 111112 75514 111152
rect 75556 111112 75596 111152
rect 75638 111112 75678 111152
rect 75720 111112 75760 111152
rect 90512 111112 90552 111152
rect 90594 111112 90634 111152
rect 90676 111112 90716 111152
rect 90758 111112 90798 111152
rect 90840 111112 90880 111152
rect 105632 111112 105672 111152
rect 105714 111112 105754 111152
rect 105796 111112 105836 111152
rect 105878 111112 105918 111152
rect 105960 111112 106000 111152
rect 120752 111112 120792 111152
rect 120834 111112 120874 111152
rect 120916 111112 120956 111152
rect 120998 111112 121038 111152
rect 121080 111112 121120 111152
rect 135872 111112 135912 111152
rect 135954 111112 135994 111152
rect 136036 111112 136076 111152
rect 136118 111112 136158 111152
rect 136200 111112 136240 111152
rect 150992 111112 151032 111152
rect 151074 111112 151114 111152
rect 151156 111112 151196 111152
rect 151238 111112 151278 111152
rect 151320 111112 151360 111152
rect 74152 110356 74192 110396
rect 74234 110356 74274 110396
rect 74316 110356 74356 110396
rect 74398 110356 74438 110396
rect 74480 110356 74520 110396
rect 89272 110356 89312 110396
rect 89354 110356 89394 110396
rect 89436 110356 89476 110396
rect 89518 110356 89558 110396
rect 89600 110356 89640 110396
rect 104392 110356 104432 110396
rect 104474 110356 104514 110396
rect 104556 110356 104596 110396
rect 104638 110356 104678 110396
rect 104720 110356 104760 110396
rect 119512 110356 119552 110396
rect 119594 110356 119634 110396
rect 119676 110356 119716 110396
rect 119758 110356 119798 110396
rect 119840 110356 119880 110396
rect 134632 110356 134672 110396
rect 134714 110356 134754 110396
rect 134796 110356 134836 110396
rect 134878 110356 134918 110396
rect 134960 110356 135000 110396
rect 149752 110356 149792 110396
rect 149834 110356 149874 110396
rect 149916 110356 149956 110396
rect 149998 110356 150038 110396
rect 150080 110356 150120 110396
rect 75392 109600 75432 109640
rect 75474 109600 75514 109640
rect 75556 109600 75596 109640
rect 75638 109600 75678 109640
rect 75720 109600 75760 109640
rect 90512 109600 90552 109640
rect 90594 109600 90634 109640
rect 90676 109600 90716 109640
rect 90758 109600 90798 109640
rect 90840 109600 90880 109640
rect 105632 109600 105672 109640
rect 105714 109600 105754 109640
rect 105796 109600 105836 109640
rect 105878 109600 105918 109640
rect 105960 109600 106000 109640
rect 120752 109600 120792 109640
rect 120834 109600 120874 109640
rect 120916 109600 120956 109640
rect 120998 109600 121038 109640
rect 121080 109600 121120 109640
rect 135872 109600 135912 109640
rect 135954 109600 135994 109640
rect 136036 109600 136076 109640
rect 136118 109600 136158 109640
rect 136200 109600 136240 109640
rect 150992 109600 151032 109640
rect 151074 109600 151114 109640
rect 151156 109600 151196 109640
rect 151238 109600 151278 109640
rect 151320 109600 151360 109640
rect 74152 108844 74192 108884
rect 74234 108844 74274 108884
rect 74316 108844 74356 108884
rect 74398 108844 74438 108884
rect 74480 108844 74520 108884
rect 89272 108844 89312 108884
rect 89354 108844 89394 108884
rect 89436 108844 89476 108884
rect 89518 108844 89558 108884
rect 89600 108844 89640 108884
rect 104392 108844 104432 108884
rect 104474 108844 104514 108884
rect 104556 108844 104596 108884
rect 104638 108844 104678 108884
rect 104720 108844 104760 108884
rect 119512 108844 119552 108884
rect 119594 108844 119634 108884
rect 119676 108844 119716 108884
rect 119758 108844 119798 108884
rect 119840 108844 119880 108884
rect 134632 108844 134672 108884
rect 134714 108844 134754 108884
rect 134796 108844 134836 108884
rect 134878 108844 134918 108884
rect 134960 108844 135000 108884
rect 149752 108844 149792 108884
rect 149834 108844 149874 108884
rect 149916 108844 149956 108884
rect 149998 108844 150038 108884
rect 150080 108844 150120 108884
rect 75392 108088 75432 108128
rect 75474 108088 75514 108128
rect 75556 108088 75596 108128
rect 75638 108088 75678 108128
rect 75720 108088 75760 108128
rect 90512 108088 90552 108128
rect 90594 108088 90634 108128
rect 90676 108088 90716 108128
rect 90758 108088 90798 108128
rect 90840 108088 90880 108128
rect 105632 108088 105672 108128
rect 105714 108088 105754 108128
rect 105796 108088 105836 108128
rect 105878 108088 105918 108128
rect 105960 108088 106000 108128
rect 120752 108088 120792 108128
rect 120834 108088 120874 108128
rect 120916 108088 120956 108128
rect 120998 108088 121038 108128
rect 121080 108088 121120 108128
rect 135872 108088 135912 108128
rect 135954 108088 135994 108128
rect 136036 108088 136076 108128
rect 136118 108088 136158 108128
rect 136200 108088 136240 108128
rect 150992 108088 151032 108128
rect 151074 108088 151114 108128
rect 151156 108088 151196 108128
rect 151238 108088 151278 108128
rect 151320 108088 151360 108128
rect 74152 107332 74192 107372
rect 74234 107332 74274 107372
rect 74316 107332 74356 107372
rect 74398 107332 74438 107372
rect 74480 107332 74520 107372
rect 89272 107332 89312 107372
rect 89354 107332 89394 107372
rect 89436 107332 89476 107372
rect 89518 107332 89558 107372
rect 89600 107332 89640 107372
rect 104392 107332 104432 107372
rect 104474 107332 104514 107372
rect 104556 107332 104596 107372
rect 104638 107332 104678 107372
rect 104720 107332 104760 107372
rect 119512 107332 119552 107372
rect 119594 107332 119634 107372
rect 119676 107332 119716 107372
rect 119758 107332 119798 107372
rect 119840 107332 119880 107372
rect 134632 107332 134672 107372
rect 134714 107332 134754 107372
rect 134796 107332 134836 107372
rect 134878 107332 134918 107372
rect 134960 107332 135000 107372
rect 149752 107332 149792 107372
rect 149834 107332 149874 107372
rect 149916 107332 149956 107372
rect 149998 107332 150038 107372
rect 150080 107332 150120 107372
rect 75392 106576 75432 106616
rect 75474 106576 75514 106616
rect 75556 106576 75596 106616
rect 75638 106576 75678 106616
rect 75720 106576 75760 106616
rect 90512 106576 90552 106616
rect 90594 106576 90634 106616
rect 90676 106576 90716 106616
rect 90758 106576 90798 106616
rect 90840 106576 90880 106616
rect 105632 106576 105672 106616
rect 105714 106576 105754 106616
rect 105796 106576 105836 106616
rect 105878 106576 105918 106616
rect 105960 106576 106000 106616
rect 120752 106576 120792 106616
rect 120834 106576 120874 106616
rect 120916 106576 120956 106616
rect 120998 106576 121038 106616
rect 121080 106576 121120 106616
rect 135872 106576 135912 106616
rect 135954 106576 135994 106616
rect 136036 106576 136076 106616
rect 136118 106576 136158 106616
rect 136200 106576 136240 106616
rect 150992 106576 151032 106616
rect 151074 106576 151114 106616
rect 151156 106576 151196 106616
rect 151238 106576 151278 106616
rect 151320 106576 151360 106616
rect 74152 105820 74192 105860
rect 74234 105820 74274 105860
rect 74316 105820 74356 105860
rect 74398 105820 74438 105860
rect 74480 105820 74520 105860
rect 89272 105820 89312 105860
rect 89354 105820 89394 105860
rect 89436 105820 89476 105860
rect 89518 105820 89558 105860
rect 89600 105820 89640 105860
rect 104392 105820 104432 105860
rect 104474 105820 104514 105860
rect 104556 105820 104596 105860
rect 104638 105820 104678 105860
rect 104720 105820 104760 105860
rect 119512 105820 119552 105860
rect 119594 105820 119634 105860
rect 119676 105820 119716 105860
rect 119758 105820 119798 105860
rect 119840 105820 119880 105860
rect 134632 105820 134672 105860
rect 134714 105820 134754 105860
rect 134796 105820 134836 105860
rect 134878 105820 134918 105860
rect 134960 105820 135000 105860
rect 149752 105820 149792 105860
rect 149834 105820 149874 105860
rect 149916 105820 149956 105860
rect 149998 105820 150038 105860
rect 150080 105820 150120 105860
rect 75392 105064 75432 105104
rect 75474 105064 75514 105104
rect 75556 105064 75596 105104
rect 75638 105064 75678 105104
rect 75720 105064 75760 105104
rect 90512 105064 90552 105104
rect 90594 105064 90634 105104
rect 90676 105064 90716 105104
rect 90758 105064 90798 105104
rect 90840 105064 90880 105104
rect 105632 105064 105672 105104
rect 105714 105064 105754 105104
rect 105796 105064 105836 105104
rect 105878 105064 105918 105104
rect 105960 105064 106000 105104
rect 120752 105064 120792 105104
rect 120834 105064 120874 105104
rect 120916 105064 120956 105104
rect 120998 105064 121038 105104
rect 121080 105064 121120 105104
rect 135872 105064 135912 105104
rect 135954 105064 135994 105104
rect 136036 105064 136076 105104
rect 136118 105064 136158 105104
rect 136200 105064 136240 105104
rect 150992 105064 151032 105104
rect 151074 105064 151114 105104
rect 151156 105064 151196 105104
rect 151238 105064 151278 105104
rect 151320 105064 151360 105104
rect 74152 104308 74192 104348
rect 74234 104308 74274 104348
rect 74316 104308 74356 104348
rect 74398 104308 74438 104348
rect 74480 104308 74520 104348
rect 89272 104308 89312 104348
rect 89354 104308 89394 104348
rect 89436 104308 89476 104348
rect 89518 104308 89558 104348
rect 89600 104308 89640 104348
rect 104392 104308 104432 104348
rect 104474 104308 104514 104348
rect 104556 104308 104596 104348
rect 104638 104308 104678 104348
rect 104720 104308 104760 104348
rect 119512 104308 119552 104348
rect 119594 104308 119634 104348
rect 119676 104308 119716 104348
rect 119758 104308 119798 104348
rect 119840 104308 119880 104348
rect 134632 104308 134672 104348
rect 134714 104308 134754 104348
rect 134796 104308 134836 104348
rect 134878 104308 134918 104348
rect 134960 104308 135000 104348
rect 149752 104308 149792 104348
rect 149834 104308 149874 104348
rect 149916 104308 149956 104348
rect 149998 104308 150038 104348
rect 150080 104308 150120 104348
rect 75392 103552 75432 103592
rect 75474 103552 75514 103592
rect 75556 103552 75596 103592
rect 75638 103552 75678 103592
rect 75720 103552 75760 103592
rect 90512 103552 90552 103592
rect 90594 103552 90634 103592
rect 90676 103552 90716 103592
rect 90758 103552 90798 103592
rect 90840 103552 90880 103592
rect 105632 103552 105672 103592
rect 105714 103552 105754 103592
rect 105796 103552 105836 103592
rect 105878 103552 105918 103592
rect 105960 103552 106000 103592
rect 120752 103552 120792 103592
rect 120834 103552 120874 103592
rect 120916 103552 120956 103592
rect 120998 103552 121038 103592
rect 121080 103552 121120 103592
rect 135872 103552 135912 103592
rect 135954 103552 135994 103592
rect 136036 103552 136076 103592
rect 136118 103552 136158 103592
rect 136200 103552 136240 103592
rect 150992 103552 151032 103592
rect 151074 103552 151114 103592
rect 151156 103552 151196 103592
rect 151238 103552 151278 103592
rect 151320 103552 151360 103592
rect 74152 102796 74192 102836
rect 74234 102796 74274 102836
rect 74316 102796 74356 102836
rect 74398 102796 74438 102836
rect 74480 102796 74520 102836
rect 89272 102796 89312 102836
rect 89354 102796 89394 102836
rect 89436 102796 89476 102836
rect 89518 102796 89558 102836
rect 89600 102796 89640 102836
rect 104392 102796 104432 102836
rect 104474 102796 104514 102836
rect 104556 102796 104596 102836
rect 104638 102796 104678 102836
rect 104720 102796 104760 102836
rect 119512 102796 119552 102836
rect 119594 102796 119634 102836
rect 119676 102796 119716 102836
rect 119758 102796 119798 102836
rect 119840 102796 119880 102836
rect 134632 102796 134672 102836
rect 134714 102796 134754 102836
rect 134796 102796 134836 102836
rect 134878 102796 134918 102836
rect 134960 102796 135000 102836
rect 149752 102796 149792 102836
rect 149834 102796 149874 102836
rect 149916 102796 149956 102836
rect 149998 102796 150038 102836
rect 150080 102796 150120 102836
rect 75392 102040 75432 102080
rect 75474 102040 75514 102080
rect 75556 102040 75596 102080
rect 75638 102040 75678 102080
rect 75720 102040 75760 102080
rect 90512 102040 90552 102080
rect 90594 102040 90634 102080
rect 90676 102040 90716 102080
rect 90758 102040 90798 102080
rect 90840 102040 90880 102080
rect 105632 102040 105672 102080
rect 105714 102040 105754 102080
rect 105796 102040 105836 102080
rect 105878 102040 105918 102080
rect 105960 102040 106000 102080
rect 120752 102040 120792 102080
rect 120834 102040 120874 102080
rect 120916 102040 120956 102080
rect 120998 102040 121038 102080
rect 121080 102040 121120 102080
rect 135872 102040 135912 102080
rect 135954 102040 135994 102080
rect 136036 102040 136076 102080
rect 136118 102040 136158 102080
rect 136200 102040 136240 102080
rect 150992 102040 151032 102080
rect 151074 102040 151114 102080
rect 151156 102040 151196 102080
rect 151238 102040 151278 102080
rect 151320 102040 151360 102080
rect 74152 101284 74192 101324
rect 74234 101284 74274 101324
rect 74316 101284 74356 101324
rect 74398 101284 74438 101324
rect 74480 101284 74520 101324
rect 89272 101284 89312 101324
rect 89354 101284 89394 101324
rect 89436 101284 89476 101324
rect 89518 101284 89558 101324
rect 89600 101284 89640 101324
rect 104392 101284 104432 101324
rect 104474 101284 104514 101324
rect 104556 101284 104596 101324
rect 104638 101284 104678 101324
rect 104720 101284 104760 101324
rect 119512 101284 119552 101324
rect 119594 101284 119634 101324
rect 119676 101284 119716 101324
rect 119758 101284 119798 101324
rect 119840 101284 119880 101324
rect 134632 101284 134672 101324
rect 134714 101284 134754 101324
rect 134796 101284 134836 101324
rect 134878 101284 134918 101324
rect 134960 101284 135000 101324
rect 149752 101284 149792 101324
rect 149834 101284 149874 101324
rect 149916 101284 149956 101324
rect 149998 101284 150038 101324
rect 150080 101284 150120 101324
rect 75392 100528 75432 100568
rect 75474 100528 75514 100568
rect 75556 100528 75596 100568
rect 75638 100528 75678 100568
rect 75720 100528 75760 100568
rect 90512 100528 90552 100568
rect 90594 100528 90634 100568
rect 90676 100528 90716 100568
rect 90758 100528 90798 100568
rect 90840 100528 90880 100568
rect 105632 100528 105672 100568
rect 105714 100528 105754 100568
rect 105796 100528 105836 100568
rect 105878 100528 105918 100568
rect 105960 100528 106000 100568
rect 120752 100528 120792 100568
rect 120834 100528 120874 100568
rect 120916 100528 120956 100568
rect 120998 100528 121038 100568
rect 121080 100528 121120 100568
rect 135872 100528 135912 100568
rect 135954 100528 135994 100568
rect 136036 100528 136076 100568
rect 136118 100528 136158 100568
rect 136200 100528 136240 100568
rect 150992 100528 151032 100568
rect 151074 100528 151114 100568
rect 151156 100528 151196 100568
rect 151238 100528 151278 100568
rect 151320 100528 151360 100568
rect 74152 99772 74192 99812
rect 74234 99772 74274 99812
rect 74316 99772 74356 99812
rect 74398 99772 74438 99812
rect 74480 99772 74520 99812
rect 89272 99772 89312 99812
rect 89354 99772 89394 99812
rect 89436 99772 89476 99812
rect 89518 99772 89558 99812
rect 89600 99772 89640 99812
rect 104392 99772 104432 99812
rect 104474 99772 104514 99812
rect 104556 99772 104596 99812
rect 104638 99772 104678 99812
rect 104720 99772 104760 99812
rect 119512 99772 119552 99812
rect 119594 99772 119634 99812
rect 119676 99772 119716 99812
rect 119758 99772 119798 99812
rect 119840 99772 119880 99812
rect 134632 99772 134672 99812
rect 134714 99772 134754 99812
rect 134796 99772 134836 99812
rect 134878 99772 134918 99812
rect 134960 99772 135000 99812
rect 149752 99772 149792 99812
rect 149834 99772 149874 99812
rect 149916 99772 149956 99812
rect 149998 99772 150038 99812
rect 150080 99772 150120 99812
rect 75392 99016 75432 99056
rect 75474 99016 75514 99056
rect 75556 99016 75596 99056
rect 75638 99016 75678 99056
rect 75720 99016 75760 99056
rect 90512 99016 90552 99056
rect 90594 99016 90634 99056
rect 90676 99016 90716 99056
rect 90758 99016 90798 99056
rect 90840 99016 90880 99056
rect 105632 99016 105672 99056
rect 105714 99016 105754 99056
rect 105796 99016 105836 99056
rect 105878 99016 105918 99056
rect 105960 99016 106000 99056
rect 120752 99016 120792 99056
rect 120834 99016 120874 99056
rect 120916 99016 120956 99056
rect 120998 99016 121038 99056
rect 121080 99016 121120 99056
rect 135872 99016 135912 99056
rect 135954 99016 135994 99056
rect 136036 99016 136076 99056
rect 136118 99016 136158 99056
rect 136200 99016 136240 99056
rect 150992 99016 151032 99056
rect 151074 99016 151114 99056
rect 151156 99016 151196 99056
rect 151238 99016 151278 99056
rect 151320 99016 151360 99056
rect 74152 98260 74192 98300
rect 74234 98260 74274 98300
rect 74316 98260 74356 98300
rect 74398 98260 74438 98300
rect 74480 98260 74520 98300
rect 89272 98260 89312 98300
rect 89354 98260 89394 98300
rect 89436 98260 89476 98300
rect 89518 98260 89558 98300
rect 89600 98260 89640 98300
rect 104392 98260 104432 98300
rect 104474 98260 104514 98300
rect 104556 98260 104596 98300
rect 104638 98260 104678 98300
rect 104720 98260 104760 98300
rect 119512 98260 119552 98300
rect 119594 98260 119634 98300
rect 119676 98260 119716 98300
rect 119758 98260 119798 98300
rect 119840 98260 119880 98300
rect 134632 98260 134672 98300
rect 134714 98260 134754 98300
rect 134796 98260 134836 98300
rect 134878 98260 134918 98300
rect 134960 98260 135000 98300
rect 149752 98260 149792 98300
rect 149834 98260 149874 98300
rect 149916 98260 149956 98300
rect 149998 98260 150038 98300
rect 150080 98260 150120 98300
rect 75392 97504 75432 97544
rect 75474 97504 75514 97544
rect 75556 97504 75596 97544
rect 75638 97504 75678 97544
rect 75720 97504 75760 97544
rect 90512 97504 90552 97544
rect 90594 97504 90634 97544
rect 90676 97504 90716 97544
rect 90758 97504 90798 97544
rect 90840 97504 90880 97544
rect 105632 97504 105672 97544
rect 105714 97504 105754 97544
rect 105796 97504 105836 97544
rect 105878 97504 105918 97544
rect 105960 97504 106000 97544
rect 120752 97504 120792 97544
rect 120834 97504 120874 97544
rect 120916 97504 120956 97544
rect 120998 97504 121038 97544
rect 121080 97504 121120 97544
rect 135872 97504 135912 97544
rect 135954 97504 135994 97544
rect 136036 97504 136076 97544
rect 136118 97504 136158 97544
rect 136200 97504 136240 97544
rect 150992 97504 151032 97544
rect 151074 97504 151114 97544
rect 151156 97504 151196 97544
rect 151238 97504 151278 97544
rect 151320 97504 151360 97544
rect 74152 96748 74192 96788
rect 74234 96748 74274 96788
rect 74316 96748 74356 96788
rect 74398 96748 74438 96788
rect 74480 96748 74520 96788
rect 89272 96748 89312 96788
rect 89354 96748 89394 96788
rect 89436 96748 89476 96788
rect 89518 96748 89558 96788
rect 89600 96748 89640 96788
rect 104392 96748 104432 96788
rect 104474 96748 104514 96788
rect 104556 96748 104596 96788
rect 104638 96748 104678 96788
rect 104720 96748 104760 96788
rect 119512 96748 119552 96788
rect 119594 96748 119634 96788
rect 119676 96748 119716 96788
rect 119758 96748 119798 96788
rect 119840 96748 119880 96788
rect 134632 96748 134672 96788
rect 134714 96748 134754 96788
rect 134796 96748 134836 96788
rect 134878 96748 134918 96788
rect 134960 96748 135000 96788
rect 149752 96748 149792 96788
rect 149834 96748 149874 96788
rect 149916 96748 149956 96788
rect 149998 96748 150038 96788
rect 150080 96748 150120 96788
rect 75392 95992 75432 96032
rect 75474 95992 75514 96032
rect 75556 95992 75596 96032
rect 75638 95992 75678 96032
rect 75720 95992 75760 96032
rect 90512 95992 90552 96032
rect 90594 95992 90634 96032
rect 90676 95992 90716 96032
rect 90758 95992 90798 96032
rect 90840 95992 90880 96032
rect 105632 95992 105672 96032
rect 105714 95992 105754 96032
rect 105796 95992 105836 96032
rect 105878 95992 105918 96032
rect 105960 95992 106000 96032
rect 120752 95992 120792 96032
rect 120834 95992 120874 96032
rect 120916 95992 120956 96032
rect 120998 95992 121038 96032
rect 121080 95992 121120 96032
rect 135872 95992 135912 96032
rect 135954 95992 135994 96032
rect 136036 95992 136076 96032
rect 136118 95992 136158 96032
rect 136200 95992 136240 96032
rect 150992 95992 151032 96032
rect 151074 95992 151114 96032
rect 151156 95992 151196 96032
rect 151238 95992 151278 96032
rect 151320 95992 151360 96032
rect 74152 95236 74192 95276
rect 74234 95236 74274 95276
rect 74316 95236 74356 95276
rect 74398 95236 74438 95276
rect 74480 95236 74520 95276
rect 89272 95236 89312 95276
rect 89354 95236 89394 95276
rect 89436 95236 89476 95276
rect 89518 95236 89558 95276
rect 89600 95236 89640 95276
rect 104392 95236 104432 95276
rect 104474 95236 104514 95276
rect 104556 95236 104596 95276
rect 104638 95236 104678 95276
rect 104720 95236 104760 95276
rect 119512 95236 119552 95276
rect 119594 95236 119634 95276
rect 119676 95236 119716 95276
rect 119758 95236 119798 95276
rect 119840 95236 119880 95276
rect 134632 95236 134672 95276
rect 134714 95236 134754 95276
rect 134796 95236 134836 95276
rect 134878 95236 134918 95276
rect 134960 95236 135000 95276
rect 149752 95236 149792 95276
rect 149834 95236 149874 95276
rect 149916 95236 149956 95276
rect 149998 95236 150038 95276
rect 150080 95236 150120 95276
rect 75392 94480 75432 94520
rect 75474 94480 75514 94520
rect 75556 94480 75596 94520
rect 75638 94480 75678 94520
rect 75720 94480 75760 94520
rect 90512 94480 90552 94520
rect 90594 94480 90634 94520
rect 90676 94480 90716 94520
rect 90758 94480 90798 94520
rect 90840 94480 90880 94520
rect 105632 94480 105672 94520
rect 105714 94480 105754 94520
rect 105796 94480 105836 94520
rect 105878 94480 105918 94520
rect 105960 94480 106000 94520
rect 120752 94480 120792 94520
rect 120834 94480 120874 94520
rect 120916 94480 120956 94520
rect 120998 94480 121038 94520
rect 121080 94480 121120 94520
rect 135872 94480 135912 94520
rect 135954 94480 135994 94520
rect 136036 94480 136076 94520
rect 136118 94480 136158 94520
rect 136200 94480 136240 94520
rect 150992 94480 151032 94520
rect 151074 94480 151114 94520
rect 151156 94480 151196 94520
rect 151238 94480 151278 94520
rect 151320 94480 151360 94520
rect 74152 93724 74192 93764
rect 74234 93724 74274 93764
rect 74316 93724 74356 93764
rect 74398 93724 74438 93764
rect 74480 93724 74520 93764
rect 89272 93724 89312 93764
rect 89354 93724 89394 93764
rect 89436 93724 89476 93764
rect 89518 93724 89558 93764
rect 89600 93724 89640 93764
rect 104392 93724 104432 93764
rect 104474 93724 104514 93764
rect 104556 93724 104596 93764
rect 104638 93724 104678 93764
rect 104720 93724 104760 93764
rect 119512 93724 119552 93764
rect 119594 93724 119634 93764
rect 119676 93724 119716 93764
rect 119758 93724 119798 93764
rect 119840 93724 119880 93764
rect 134632 93724 134672 93764
rect 134714 93724 134754 93764
rect 134796 93724 134836 93764
rect 134878 93724 134918 93764
rect 134960 93724 135000 93764
rect 149752 93724 149792 93764
rect 149834 93724 149874 93764
rect 149916 93724 149956 93764
rect 149998 93724 150038 93764
rect 150080 93724 150120 93764
rect 75392 92968 75432 93008
rect 75474 92968 75514 93008
rect 75556 92968 75596 93008
rect 75638 92968 75678 93008
rect 75720 92968 75760 93008
rect 90512 92968 90552 93008
rect 90594 92968 90634 93008
rect 90676 92968 90716 93008
rect 90758 92968 90798 93008
rect 90840 92968 90880 93008
rect 105632 92968 105672 93008
rect 105714 92968 105754 93008
rect 105796 92968 105836 93008
rect 105878 92968 105918 93008
rect 105960 92968 106000 93008
rect 120752 92968 120792 93008
rect 120834 92968 120874 93008
rect 120916 92968 120956 93008
rect 120998 92968 121038 93008
rect 121080 92968 121120 93008
rect 135872 92968 135912 93008
rect 135954 92968 135994 93008
rect 136036 92968 136076 93008
rect 136118 92968 136158 93008
rect 136200 92968 136240 93008
rect 150992 92968 151032 93008
rect 151074 92968 151114 93008
rect 151156 92968 151196 93008
rect 151238 92968 151278 93008
rect 151320 92968 151360 93008
rect 74152 92212 74192 92252
rect 74234 92212 74274 92252
rect 74316 92212 74356 92252
rect 74398 92212 74438 92252
rect 74480 92212 74520 92252
rect 89272 92212 89312 92252
rect 89354 92212 89394 92252
rect 89436 92212 89476 92252
rect 89518 92212 89558 92252
rect 89600 92212 89640 92252
rect 104392 92212 104432 92252
rect 104474 92212 104514 92252
rect 104556 92212 104596 92252
rect 104638 92212 104678 92252
rect 104720 92212 104760 92252
rect 119512 92212 119552 92252
rect 119594 92212 119634 92252
rect 119676 92212 119716 92252
rect 119758 92212 119798 92252
rect 119840 92212 119880 92252
rect 134632 92212 134672 92252
rect 134714 92212 134754 92252
rect 134796 92212 134836 92252
rect 134878 92212 134918 92252
rect 134960 92212 135000 92252
rect 149752 92212 149792 92252
rect 149834 92212 149874 92252
rect 149916 92212 149956 92252
rect 149998 92212 150038 92252
rect 150080 92212 150120 92252
rect 75392 91456 75432 91496
rect 75474 91456 75514 91496
rect 75556 91456 75596 91496
rect 75638 91456 75678 91496
rect 75720 91456 75760 91496
rect 90512 91456 90552 91496
rect 90594 91456 90634 91496
rect 90676 91456 90716 91496
rect 90758 91456 90798 91496
rect 90840 91456 90880 91496
rect 105632 91456 105672 91496
rect 105714 91456 105754 91496
rect 105796 91456 105836 91496
rect 105878 91456 105918 91496
rect 105960 91456 106000 91496
rect 120752 91456 120792 91496
rect 120834 91456 120874 91496
rect 120916 91456 120956 91496
rect 120998 91456 121038 91496
rect 121080 91456 121120 91496
rect 135872 91456 135912 91496
rect 135954 91456 135994 91496
rect 136036 91456 136076 91496
rect 136118 91456 136158 91496
rect 136200 91456 136240 91496
rect 150992 91456 151032 91496
rect 151074 91456 151114 91496
rect 151156 91456 151196 91496
rect 151238 91456 151278 91496
rect 151320 91456 151360 91496
rect 74152 90700 74192 90740
rect 74234 90700 74274 90740
rect 74316 90700 74356 90740
rect 74398 90700 74438 90740
rect 74480 90700 74520 90740
rect 89272 90700 89312 90740
rect 89354 90700 89394 90740
rect 89436 90700 89476 90740
rect 89518 90700 89558 90740
rect 89600 90700 89640 90740
rect 104392 90700 104432 90740
rect 104474 90700 104514 90740
rect 104556 90700 104596 90740
rect 104638 90700 104678 90740
rect 104720 90700 104760 90740
rect 119512 90700 119552 90740
rect 119594 90700 119634 90740
rect 119676 90700 119716 90740
rect 119758 90700 119798 90740
rect 119840 90700 119880 90740
rect 134632 90700 134672 90740
rect 134714 90700 134754 90740
rect 134796 90700 134836 90740
rect 134878 90700 134918 90740
rect 134960 90700 135000 90740
rect 149752 90700 149792 90740
rect 149834 90700 149874 90740
rect 149916 90700 149956 90740
rect 149998 90700 150038 90740
rect 150080 90700 150120 90740
rect 75392 89944 75432 89984
rect 75474 89944 75514 89984
rect 75556 89944 75596 89984
rect 75638 89944 75678 89984
rect 75720 89944 75760 89984
rect 90512 89944 90552 89984
rect 90594 89944 90634 89984
rect 90676 89944 90716 89984
rect 90758 89944 90798 89984
rect 90840 89944 90880 89984
rect 105632 89944 105672 89984
rect 105714 89944 105754 89984
rect 105796 89944 105836 89984
rect 105878 89944 105918 89984
rect 105960 89944 106000 89984
rect 120752 89944 120792 89984
rect 120834 89944 120874 89984
rect 120916 89944 120956 89984
rect 120998 89944 121038 89984
rect 121080 89944 121120 89984
rect 135872 89944 135912 89984
rect 135954 89944 135994 89984
rect 136036 89944 136076 89984
rect 136118 89944 136158 89984
rect 136200 89944 136240 89984
rect 150992 89944 151032 89984
rect 151074 89944 151114 89984
rect 151156 89944 151196 89984
rect 151238 89944 151278 89984
rect 151320 89944 151360 89984
rect 74152 89188 74192 89228
rect 74234 89188 74274 89228
rect 74316 89188 74356 89228
rect 74398 89188 74438 89228
rect 74480 89188 74520 89228
rect 89272 89188 89312 89228
rect 89354 89188 89394 89228
rect 89436 89188 89476 89228
rect 89518 89188 89558 89228
rect 89600 89188 89640 89228
rect 104392 89188 104432 89228
rect 104474 89188 104514 89228
rect 104556 89188 104596 89228
rect 104638 89188 104678 89228
rect 104720 89188 104760 89228
rect 119512 89188 119552 89228
rect 119594 89188 119634 89228
rect 119676 89188 119716 89228
rect 119758 89188 119798 89228
rect 119840 89188 119880 89228
rect 134632 89188 134672 89228
rect 134714 89188 134754 89228
rect 134796 89188 134836 89228
rect 134878 89188 134918 89228
rect 134960 89188 135000 89228
rect 149752 89188 149792 89228
rect 149834 89188 149874 89228
rect 149916 89188 149956 89228
rect 149998 89188 150038 89228
rect 150080 89188 150120 89228
rect 75392 88432 75432 88472
rect 75474 88432 75514 88472
rect 75556 88432 75596 88472
rect 75638 88432 75678 88472
rect 75720 88432 75760 88472
rect 90512 88432 90552 88472
rect 90594 88432 90634 88472
rect 90676 88432 90716 88472
rect 90758 88432 90798 88472
rect 90840 88432 90880 88472
rect 105632 88432 105672 88472
rect 105714 88432 105754 88472
rect 105796 88432 105836 88472
rect 105878 88432 105918 88472
rect 105960 88432 106000 88472
rect 120752 88432 120792 88472
rect 120834 88432 120874 88472
rect 120916 88432 120956 88472
rect 120998 88432 121038 88472
rect 121080 88432 121120 88472
rect 135872 88432 135912 88472
rect 135954 88432 135994 88472
rect 136036 88432 136076 88472
rect 136118 88432 136158 88472
rect 136200 88432 136240 88472
rect 150992 88432 151032 88472
rect 151074 88432 151114 88472
rect 151156 88432 151196 88472
rect 151238 88432 151278 88472
rect 151320 88432 151360 88472
rect 74152 87676 74192 87716
rect 74234 87676 74274 87716
rect 74316 87676 74356 87716
rect 74398 87676 74438 87716
rect 74480 87676 74520 87716
rect 89272 87676 89312 87716
rect 89354 87676 89394 87716
rect 89436 87676 89476 87716
rect 89518 87676 89558 87716
rect 89600 87676 89640 87716
rect 104392 87676 104432 87716
rect 104474 87676 104514 87716
rect 104556 87676 104596 87716
rect 104638 87676 104678 87716
rect 104720 87676 104760 87716
rect 119512 87676 119552 87716
rect 119594 87676 119634 87716
rect 119676 87676 119716 87716
rect 119758 87676 119798 87716
rect 119840 87676 119880 87716
rect 134632 87676 134672 87716
rect 134714 87676 134754 87716
rect 134796 87676 134836 87716
rect 134878 87676 134918 87716
rect 134960 87676 135000 87716
rect 149752 87676 149792 87716
rect 149834 87676 149874 87716
rect 149916 87676 149956 87716
rect 149998 87676 150038 87716
rect 150080 87676 150120 87716
rect 75392 86920 75432 86960
rect 75474 86920 75514 86960
rect 75556 86920 75596 86960
rect 75638 86920 75678 86960
rect 75720 86920 75760 86960
rect 90512 86920 90552 86960
rect 90594 86920 90634 86960
rect 90676 86920 90716 86960
rect 90758 86920 90798 86960
rect 90840 86920 90880 86960
rect 105632 86920 105672 86960
rect 105714 86920 105754 86960
rect 105796 86920 105836 86960
rect 105878 86920 105918 86960
rect 105960 86920 106000 86960
rect 120752 86920 120792 86960
rect 120834 86920 120874 86960
rect 120916 86920 120956 86960
rect 120998 86920 121038 86960
rect 121080 86920 121120 86960
rect 135872 86920 135912 86960
rect 135954 86920 135994 86960
rect 136036 86920 136076 86960
rect 136118 86920 136158 86960
rect 136200 86920 136240 86960
rect 150992 86920 151032 86960
rect 151074 86920 151114 86960
rect 151156 86920 151196 86960
rect 151238 86920 151278 86960
rect 151320 86920 151360 86960
rect 74152 86164 74192 86204
rect 74234 86164 74274 86204
rect 74316 86164 74356 86204
rect 74398 86164 74438 86204
rect 74480 86164 74520 86204
rect 89272 86164 89312 86204
rect 89354 86164 89394 86204
rect 89436 86164 89476 86204
rect 89518 86164 89558 86204
rect 89600 86164 89640 86204
rect 104392 86164 104432 86204
rect 104474 86164 104514 86204
rect 104556 86164 104596 86204
rect 104638 86164 104678 86204
rect 104720 86164 104760 86204
rect 119512 86164 119552 86204
rect 119594 86164 119634 86204
rect 119676 86164 119716 86204
rect 119758 86164 119798 86204
rect 119840 86164 119880 86204
rect 134632 86164 134672 86204
rect 134714 86164 134754 86204
rect 134796 86164 134836 86204
rect 134878 86164 134918 86204
rect 134960 86164 135000 86204
rect 149752 86164 149792 86204
rect 149834 86164 149874 86204
rect 149916 86164 149956 86204
rect 149998 86164 150038 86204
rect 150080 86164 150120 86204
rect 75392 85408 75432 85448
rect 75474 85408 75514 85448
rect 75556 85408 75596 85448
rect 75638 85408 75678 85448
rect 75720 85408 75760 85448
rect 90512 85408 90552 85448
rect 90594 85408 90634 85448
rect 90676 85408 90716 85448
rect 90758 85408 90798 85448
rect 90840 85408 90880 85448
rect 105632 85408 105672 85448
rect 105714 85408 105754 85448
rect 105796 85408 105836 85448
rect 105878 85408 105918 85448
rect 105960 85408 106000 85448
rect 120752 85408 120792 85448
rect 120834 85408 120874 85448
rect 120916 85408 120956 85448
rect 120998 85408 121038 85448
rect 121080 85408 121120 85448
rect 135872 85408 135912 85448
rect 135954 85408 135994 85448
rect 136036 85408 136076 85448
rect 136118 85408 136158 85448
rect 136200 85408 136240 85448
rect 150992 85408 151032 85448
rect 151074 85408 151114 85448
rect 151156 85408 151196 85448
rect 151238 85408 151278 85448
rect 151320 85408 151360 85448
rect 74152 84652 74192 84692
rect 74234 84652 74274 84692
rect 74316 84652 74356 84692
rect 74398 84652 74438 84692
rect 74480 84652 74520 84692
rect 89272 84652 89312 84692
rect 89354 84652 89394 84692
rect 89436 84652 89476 84692
rect 89518 84652 89558 84692
rect 89600 84652 89640 84692
rect 104392 84652 104432 84692
rect 104474 84652 104514 84692
rect 104556 84652 104596 84692
rect 104638 84652 104678 84692
rect 104720 84652 104760 84692
rect 119512 84652 119552 84692
rect 119594 84652 119634 84692
rect 119676 84652 119716 84692
rect 119758 84652 119798 84692
rect 119840 84652 119880 84692
rect 134632 84652 134672 84692
rect 134714 84652 134754 84692
rect 134796 84652 134836 84692
rect 134878 84652 134918 84692
rect 134960 84652 135000 84692
rect 149752 84652 149792 84692
rect 149834 84652 149874 84692
rect 149916 84652 149956 84692
rect 149998 84652 150038 84692
rect 150080 84652 150120 84692
rect 75392 83896 75432 83936
rect 75474 83896 75514 83936
rect 75556 83896 75596 83936
rect 75638 83896 75678 83936
rect 75720 83896 75760 83936
rect 90512 83896 90552 83936
rect 90594 83896 90634 83936
rect 90676 83896 90716 83936
rect 90758 83896 90798 83936
rect 90840 83896 90880 83936
rect 105632 83896 105672 83936
rect 105714 83896 105754 83936
rect 105796 83896 105836 83936
rect 105878 83896 105918 83936
rect 105960 83896 106000 83936
rect 120752 83896 120792 83936
rect 120834 83896 120874 83936
rect 120916 83896 120956 83936
rect 120998 83896 121038 83936
rect 121080 83896 121120 83936
rect 135872 83896 135912 83936
rect 135954 83896 135994 83936
rect 136036 83896 136076 83936
rect 136118 83896 136158 83936
rect 136200 83896 136240 83936
rect 150992 83896 151032 83936
rect 151074 83896 151114 83936
rect 151156 83896 151196 83936
rect 151238 83896 151278 83936
rect 151320 83896 151360 83936
rect 74152 83140 74192 83180
rect 74234 83140 74274 83180
rect 74316 83140 74356 83180
rect 74398 83140 74438 83180
rect 74480 83140 74520 83180
rect 89272 83140 89312 83180
rect 89354 83140 89394 83180
rect 89436 83140 89476 83180
rect 89518 83140 89558 83180
rect 89600 83140 89640 83180
rect 104392 83140 104432 83180
rect 104474 83140 104514 83180
rect 104556 83140 104596 83180
rect 104638 83140 104678 83180
rect 104720 83140 104760 83180
rect 119512 83140 119552 83180
rect 119594 83140 119634 83180
rect 119676 83140 119716 83180
rect 119758 83140 119798 83180
rect 119840 83140 119880 83180
rect 134632 83140 134672 83180
rect 134714 83140 134754 83180
rect 134796 83140 134836 83180
rect 134878 83140 134918 83180
rect 134960 83140 135000 83180
rect 149752 83140 149792 83180
rect 149834 83140 149874 83180
rect 149916 83140 149956 83180
rect 149998 83140 150038 83180
rect 150080 83140 150120 83180
rect 75392 82384 75432 82424
rect 75474 82384 75514 82424
rect 75556 82384 75596 82424
rect 75638 82384 75678 82424
rect 75720 82384 75760 82424
rect 90512 82384 90552 82424
rect 90594 82384 90634 82424
rect 90676 82384 90716 82424
rect 90758 82384 90798 82424
rect 90840 82384 90880 82424
rect 105632 82384 105672 82424
rect 105714 82384 105754 82424
rect 105796 82384 105836 82424
rect 105878 82384 105918 82424
rect 105960 82384 106000 82424
rect 120752 82384 120792 82424
rect 120834 82384 120874 82424
rect 120916 82384 120956 82424
rect 120998 82384 121038 82424
rect 121080 82384 121120 82424
rect 135872 82384 135912 82424
rect 135954 82384 135994 82424
rect 136036 82384 136076 82424
rect 136118 82384 136158 82424
rect 136200 82384 136240 82424
rect 150992 82384 151032 82424
rect 151074 82384 151114 82424
rect 151156 82384 151196 82424
rect 151238 82384 151278 82424
rect 151320 82384 151360 82424
rect 74152 81628 74192 81668
rect 74234 81628 74274 81668
rect 74316 81628 74356 81668
rect 74398 81628 74438 81668
rect 74480 81628 74520 81668
rect 89272 81628 89312 81668
rect 89354 81628 89394 81668
rect 89436 81628 89476 81668
rect 89518 81628 89558 81668
rect 89600 81628 89640 81668
rect 104392 81628 104432 81668
rect 104474 81628 104514 81668
rect 104556 81628 104596 81668
rect 104638 81628 104678 81668
rect 104720 81628 104760 81668
rect 119512 81628 119552 81668
rect 119594 81628 119634 81668
rect 119676 81628 119716 81668
rect 119758 81628 119798 81668
rect 119840 81628 119880 81668
rect 134632 81628 134672 81668
rect 134714 81628 134754 81668
rect 134796 81628 134836 81668
rect 134878 81628 134918 81668
rect 134960 81628 135000 81668
rect 149752 81628 149792 81668
rect 149834 81628 149874 81668
rect 149916 81628 149956 81668
rect 149998 81628 150038 81668
rect 150080 81628 150120 81668
rect 75392 80872 75432 80912
rect 75474 80872 75514 80912
rect 75556 80872 75596 80912
rect 75638 80872 75678 80912
rect 75720 80872 75760 80912
rect 90512 80872 90552 80912
rect 90594 80872 90634 80912
rect 90676 80872 90716 80912
rect 90758 80872 90798 80912
rect 90840 80872 90880 80912
rect 105632 80872 105672 80912
rect 105714 80872 105754 80912
rect 105796 80872 105836 80912
rect 105878 80872 105918 80912
rect 105960 80872 106000 80912
rect 120752 80872 120792 80912
rect 120834 80872 120874 80912
rect 120916 80872 120956 80912
rect 120998 80872 121038 80912
rect 121080 80872 121120 80912
rect 135872 80872 135912 80912
rect 135954 80872 135994 80912
rect 136036 80872 136076 80912
rect 136118 80872 136158 80912
rect 136200 80872 136240 80912
rect 150992 80872 151032 80912
rect 151074 80872 151114 80912
rect 151156 80872 151196 80912
rect 151238 80872 151278 80912
rect 151320 80872 151360 80912
rect 74152 80116 74192 80156
rect 74234 80116 74274 80156
rect 74316 80116 74356 80156
rect 74398 80116 74438 80156
rect 74480 80116 74520 80156
rect 89272 80116 89312 80156
rect 89354 80116 89394 80156
rect 89436 80116 89476 80156
rect 89518 80116 89558 80156
rect 89600 80116 89640 80156
rect 104392 80116 104432 80156
rect 104474 80116 104514 80156
rect 104556 80116 104596 80156
rect 104638 80116 104678 80156
rect 104720 80116 104760 80156
rect 119512 80116 119552 80156
rect 119594 80116 119634 80156
rect 119676 80116 119716 80156
rect 119758 80116 119798 80156
rect 119840 80116 119880 80156
rect 134632 80116 134672 80156
rect 134714 80116 134754 80156
rect 134796 80116 134836 80156
rect 134878 80116 134918 80156
rect 134960 80116 135000 80156
rect 149752 80116 149792 80156
rect 149834 80116 149874 80156
rect 149916 80116 149956 80156
rect 149998 80116 150038 80156
rect 150080 80116 150120 80156
rect 75392 79360 75432 79400
rect 75474 79360 75514 79400
rect 75556 79360 75596 79400
rect 75638 79360 75678 79400
rect 75720 79360 75760 79400
rect 90512 79360 90552 79400
rect 90594 79360 90634 79400
rect 90676 79360 90716 79400
rect 90758 79360 90798 79400
rect 90840 79360 90880 79400
rect 105632 79360 105672 79400
rect 105714 79360 105754 79400
rect 105796 79360 105836 79400
rect 105878 79360 105918 79400
rect 105960 79360 106000 79400
rect 120752 79360 120792 79400
rect 120834 79360 120874 79400
rect 120916 79360 120956 79400
rect 120998 79360 121038 79400
rect 121080 79360 121120 79400
rect 135872 79360 135912 79400
rect 135954 79360 135994 79400
rect 136036 79360 136076 79400
rect 136118 79360 136158 79400
rect 136200 79360 136240 79400
rect 150992 79360 151032 79400
rect 151074 79360 151114 79400
rect 151156 79360 151196 79400
rect 151238 79360 151278 79400
rect 151320 79360 151360 79400
rect 74152 78604 74192 78644
rect 74234 78604 74274 78644
rect 74316 78604 74356 78644
rect 74398 78604 74438 78644
rect 74480 78604 74520 78644
rect 89272 78604 89312 78644
rect 89354 78604 89394 78644
rect 89436 78604 89476 78644
rect 89518 78604 89558 78644
rect 89600 78604 89640 78644
rect 104392 78604 104432 78644
rect 104474 78604 104514 78644
rect 104556 78604 104596 78644
rect 104638 78604 104678 78644
rect 104720 78604 104760 78644
rect 119512 78604 119552 78644
rect 119594 78604 119634 78644
rect 119676 78604 119716 78644
rect 119758 78604 119798 78644
rect 119840 78604 119880 78644
rect 134632 78604 134672 78644
rect 134714 78604 134754 78644
rect 134796 78604 134836 78644
rect 134878 78604 134918 78644
rect 134960 78604 135000 78644
rect 149752 78604 149792 78644
rect 149834 78604 149874 78644
rect 149916 78604 149956 78644
rect 149998 78604 150038 78644
rect 150080 78604 150120 78644
rect 75392 77848 75432 77888
rect 75474 77848 75514 77888
rect 75556 77848 75596 77888
rect 75638 77848 75678 77888
rect 75720 77848 75760 77888
rect 90512 77848 90552 77888
rect 90594 77848 90634 77888
rect 90676 77848 90716 77888
rect 90758 77848 90798 77888
rect 90840 77848 90880 77888
rect 105632 77848 105672 77888
rect 105714 77848 105754 77888
rect 105796 77848 105836 77888
rect 105878 77848 105918 77888
rect 105960 77848 106000 77888
rect 120752 77848 120792 77888
rect 120834 77848 120874 77888
rect 120916 77848 120956 77888
rect 120998 77848 121038 77888
rect 121080 77848 121120 77888
rect 135872 77848 135912 77888
rect 135954 77848 135994 77888
rect 136036 77848 136076 77888
rect 136118 77848 136158 77888
rect 136200 77848 136240 77888
rect 150992 77848 151032 77888
rect 151074 77848 151114 77888
rect 151156 77848 151196 77888
rect 151238 77848 151278 77888
rect 151320 77848 151360 77888
rect 74152 77092 74192 77132
rect 74234 77092 74274 77132
rect 74316 77092 74356 77132
rect 74398 77092 74438 77132
rect 74480 77092 74520 77132
rect 89272 77092 89312 77132
rect 89354 77092 89394 77132
rect 89436 77092 89476 77132
rect 89518 77092 89558 77132
rect 89600 77092 89640 77132
rect 104392 77092 104432 77132
rect 104474 77092 104514 77132
rect 104556 77092 104596 77132
rect 104638 77092 104678 77132
rect 104720 77092 104760 77132
rect 119512 77092 119552 77132
rect 119594 77092 119634 77132
rect 119676 77092 119716 77132
rect 119758 77092 119798 77132
rect 119840 77092 119880 77132
rect 134632 77092 134672 77132
rect 134714 77092 134754 77132
rect 134796 77092 134836 77132
rect 134878 77092 134918 77132
rect 134960 77092 135000 77132
rect 149752 77092 149792 77132
rect 149834 77092 149874 77132
rect 149916 77092 149956 77132
rect 149998 77092 150038 77132
rect 150080 77092 150120 77132
rect 75392 76336 75432 76376
rect 75474 76336 75514 76376
rect 75556 76336 75596 76376
rect 75638 76336 75678 76376
rect 75720 76336 75760 76376
rect 90512 76336 90552 76376
rect 90594 76336 90634 76376
rect 90676 76336 90716 76376
rect 90758 76336 90798 76376
rect 90840 76336 90880 76376
rect 105632 76336 105672 76376
rect 105714 76336 105754 76376
rect 105796 76336 105836 76376
rect 105878 76336 105918 76376
rect 105960 76336 106000 76376
rect 120752 76336 120792 76376
rect 120834 76336 120874 76376
rect 120916 76336 120956 76376
rect 120998 76336 121038 76376
rect 121080 76336 121120 76376
rect 135872 76336 135912 76376
rect 135954 76336 135994 76376
rect 136036 76336 136076 76376
rect 136118 76336 136158 76376
rect 136200 76336 136240 76376
rect 150992 76336 151032 76376
rect 151074 76336 151114 76376
rect 151156 76336 151196 76376
rect 151238 76336 151278 76376
rect 151320 76336 151360 76376
rect 74152 75580 74192 75620
rect 74234 75580 74274 75620
rect 74316 75580 74356 75620
rect 74398 75580 74438 75620
rect 74480 75580 74520 75620
rect 89272 75580 89312 75620
rect 89354 75580 89394 75620
rect 89436 75580 89476 75620
rect 89518 75580 89558 75620
rect 89600 75580 89640 75620
rect 104392 75580 104432 75620
rect 104474 75580 104514 75620
rect 104556 75580 104596 75620
rect 104638 75580 104678 75620
rect 104720 75580 104760 75620
rect 119512 75580 119552 75620
rect 119594 75580 119634 75620
rect 119676 75580 119716 75620
rect 119758 75580 119798 75620
rect 119840 75580 119880 75620
rect 134632 75580 134672 75620
rect 134714 75580 134754 75620
rect 134796 75580 134836 75620
rect 134878 75580 134918 75620
rect 134960 75580 135000 75620
rect 149752 75580 149792 75620
rect 149834 75580 149874 75620
rect 149916 75580 149956 75620
rect 149998 75580 150038 75620
rect 150080 75580 150120 75620
rect 75392 74824 75432 74864
rect 75474 74824 75514 74864
rect 75556 74824 75596 74864
rect 75638 74824 75678 74864
rect 75720 74824 75760 74864
rect 90512 74824 90552 74864
rect 90594 74824 90634 74864
rect 90676 74824 90716 74864
rect 90758 74824 90798 74864
rect 90840 74824 90880 74864
rect 105632 74824 105672 74864
rect 105714 74824 105754 74864
rect 105796 74824 105836 74864
rect 105878 74824 105918 74864
rect 105960 74824 106000 74864
rect 120752 74824 120792 74864
rect 120834 74824 120874 74864
rect 120916 74824 120956 74864
rect 120998 74824 121038 74864
rect 121080 74824 121120 74864
rect 135872 74824 135912 74864
rect 135954 74824 135994 74864
rect 136036 74824 136076 74864
rect 136118 74824 136158 74864
rect 136200 74824 136240 74864
rect 150992 74824 151032 74864
rect 151074 74824 151114 74864
rect 151156 74824 151196 74864
rect 151238 74824 151278 74864
rect 151320 74824 151360 74864
rect 74152 74068 74192 74108
rect 74234 74068 74274 74108
rect 74316 74068 74356 74108
rect 74398 74068 74438 74108
rect 74480 74068 74520 74108
rect 89272 74068 89312 74108
rect 89354 74068 89394 74108
rect 89436 74068 89476 74108
rect 89518 74068 89558 74108
rect 89600 74068 89640 74108
rect 104392 74068 104432 74108
rect 104474 74068 104514 74108
rect 104556 74068 104596 74108
rect 104638 74068 104678 74108
rect 104720 74068 104760 74108
rect 119512 74068 119552 74108
rect 119594 74068 119634 74108
rect 119676 74068 119716 74108
rect 119758 74068 119798 74108
rect 119840 74068 119880 74108
rect 134632 74068 134672 74108
rect 134714 74068 134754 74108
rect 134796 74068 134836 74108
rect 134878 74068 134918 74108
rect 134960 74068 135000 74108
rect 149752 74068 149792 74108
rect 149834 74068 149874 74108
rect 149916 74068 149956 74108
rect 149998 74068 150038 74108
rect 150080 74068 150120 74108
rect 75392 73312 75432 73352
rect 75474 73312 75514 73352
rect 75556 73312 75596 73352
rect 75638 73312 75678 73352
rect 75720 73312 75760 73352
rect 90512 73312 90552 73352
rect 90594 73312 90634 73352
rect 90676 73312 90716 73352
rect 90758 73312 90798 73352
rect 90840 73312 90880 73352
rect 105632 73312 105672 73352
rect 105714 73312 105754 73352
rect 105796 73312 105836 73352
rect 105878 73312 105918 73352
rect 105960 73312 106000 73352
rect 120752 73312 120792 73352
rect 120834 73312 120874 73352
rect 120916 73312 120956 73352
rect 120998 73312 121038 73352
rect 121080 73312 121120 73352
rect 135872 73312 135912 73352
rect 135954 73312 135994 73352
rect 136036 73312 136076 73352
rect 136118 73312 136158 73352
rect 136200 73312 136240 73352
rect 150992 73312 151032 73352
rect 151074 73312 151114 73352
rect 151156 73312 151196 73352
rect 151238 73312 151278 73352
rect 151320 73312 151360 73352
rect 74152 72556 74192 72596
rect 74234 72556 74274 72596
rect 74316 72556 74356 72596
rect 74398 72556 74438 72596
rect 74480 72556 74520 72596
rect 89272 72556 89312 72596
rect 89354 72556 89394 72596
rect 89436 72556 89476 72596
rect 89518 72556 89558 72596
rect 89600 72556 89640 72596
rect 104392 72556 104432 72596
rect 104474 72556 104514 72596
rect 104556 72556 104596 72596
rect 104638 72556 104678 72596
rect 104720 72556 104760 72596
rect 119512 72556 119552 72596
rect 119594 72556 119634 72596
rect 119676 72556 119716 72596
rect 119758 72556 119798 72596
rect 119840 72556 119880 72596
rect 134632 72556 134672 72596
rect 134714 72556 134754 72596
rect 134796 72556 134836 72596
rect 134878 72556 134918 72596
rect 134960 72556 135000 72596
rect 149752 72556 149792 72596
rect 149834 72556 149874 72596
rect 149916 72556 149956 72596
rect 149998 72556 150038 72596
rect 150080 72556 150120 72596
rect 75392 71800 75432 71840
rect 75474 71800 75514 71840
rect 75556 71800 75596 71840
rect 75638 71800 75678 71840
rect 75720 71800 75760 71840
rect 90512 71800 90552 71840
rect 90594 71800 90634 71840
rect 90676 71800 90716 71840
rect 90758 71800 90798 71840
rect 90840 71800 90880 71840
rect 105632 71800 105672 71840
rect 105714 71800 105754 71840
rect 105796 71800 105836 71840
rect 105878 71800 105918 71840
rect 105960 71800 106000 71840
rect 120752 71800 120792 71840
rect 120834 71800 120874 71840
rect 120916 71800 120956 71840
rect 120998 71800 121038 71840
rect 121080 71800 121120 71840
rect 135872 71800 135912 71840
rect 135954 71800 135994 71840
rect 136036 71800 136076 71840
rect 136118 71800 136158 71840
rect 136200 71800 136240 71840
rect 150992 71800 151032 71840
rect 151074 71800 151114 71840
rect 151156 71800 151196 71840
rect 151238 71800 151278 71840
rect 151320 71800 151360 71840
<< metal2 >>
rect 103660 159461 103700 160020
rect 71979 159452 72021 159461
rect 71979 159412 71980 159452
rect 72020 159412 72021 159452
rect 71979 159403 72021 159412
rect 103659 159452 103701 159461
rect 103659 159412 103660 159452
rect 103700 159412 103701 159452
rect 103659 159403 103701 159412
rect 104043 159452 104085 159461
rect 104043 159412 104044 159452
rect 104084 159412 104085 159452
rect 104043 159403 104085 159412
rect 64107 152060 64149 152069
rect 64107 152020 64108 152060
rect 64148 152020 64149 152060
rect 64107 152018 64149 152020
rect 63984 152011 64149 152018
rect 63984 151978 64148 152011
rect 64107 136016 64149 136025
rect 63984 135976 64108 136016
rect 64148 135976 64149 136016
rect 64107 135967 64149 135976
rect 64107 120056 64149 120065
rect 64107 120016 64108 120056
rect 64148 120016 64149 120056
rect 64107 120014 64149 120016
rect 63984 120007 64149 120014
rect 63984 119974 64148 120007
rect 64107 104012 64149 104021
rect 63984 103972 64108 104012
rect 64148 103972 64149 104012
rect 64107 103963 64149 103972
rect 64107 88052 64149 88061
rect 64107 88012 64108 88052
rect 64148 88012 64149 88052
rect 64107 88010 64149 88012
rect 63984 88003 64149 88010
rect 63984 87970 64148 88003
rect 64107 72008 64149 72017
rect 63984 71968 64108 72008
rect 64148 71968 64149 72008
rect 64107 71959 64149 71968
rect 71980 64364 72020 159403
rect 88011 159368 88053 159377
rect 88011 159328 88012 159368
rect 88052 159328 88053 159368
rect 88011 159319 88053 159328
rect 75392 151976 75760 151985
rect 75432 151936 75474 151976
rect 75514 151936 75556 151976
rect 75596 151936 75638 151976
rect 75678 151936 75720 151976
rect 75392 151927 75760 151936
rect 74152 151220 74520 151229
rect 74192 151180 74234 151220
rect 74274 151180 74316 151220
rect 74356 151180 74398 151220
rect 74438 151180 74480 151220
rect 74152 151171 74520 151180
rect 75392 150464 75760 150473
rect 75432 150424 75474 150464
rect 75514 150424 75556 150464
rect 75596 150424 75638 150464
rect 75678 150424 75720 150464
rect 75392 150415 75760 150424
rect 74152 149708 74520 149717
rect 74192 149668 74234 149708
rect 74274 149668 74316 149708
rect 74356 149668 74398 149708
rect 74438 149668 74480 149708
rect 74152 149659 74520 149668
rect 75392 148952 75760 148961
rect 75432 148912 75474 148952
rect 75514 148912 75556 148952
rect 75596 148912 75638 148952
rect 75678 148912 75720 148952
rect 75392 148903 75760 148912
rect 74152 148196 74520 148205
rect 74192 148156 74234 148196
rect 74274 148156 74316 148196
rect 74356 148156 74398 148196
rect 74438 148156 74480 148196
rect 74152 148147 74520 148156
rect 75392 147440 75760 147449
rect 75432 147400 75474 147440
rect 75514 147400 75556 147440
rect 75596 147400 75638 147440
rect 75678 147400 75720 147440
rect 75392 147391 75760 147400
rect 74152 146684 74520 146693
rect 74192 146644 74234 146684
rect 74274 146644 74316 146684
rect 74356 146644 74398 146684
rect 74438 146644 74480 146684
rect 74152 146635 74520 146644
rect 75392 145928 75760 145937
rect 75432 145888 75474 145928
rect 75514 145888 75556 145928
rect 75596 145888 75638 145928
rect 75678 145888 75720 145928
rect 75392 145879 75760 145888
rect 74152 145172 74520 145181
rect 74192 145132 74234 145172
rect 74274 145132 74316 145172
rect 74356 145132 74398 145172
rect 74438 145132 74480 145172
rect 74152 145123 74520 145132
rect 75392 144416 75760 144425
rect 75432 144376 75474 144416
rect 75514 144376 75556 144416
rect 75596 144376 75638 144416
rect 75678 144376 75720 144416
rect 75392 144367 75760 144376
rect 74152 143660 74520 143669
rect 74192 143620 74234 143660
rect 74274 143620 74316 143660
rect 74356 143620 74398 143660
rect 74438 143620 74480 143660
rect 74152 143611 74520 143620
rect 75392 142904 75760 142913
rect 75432 142864 75474 142904
rect 75514 142864 75556 142904
rect 75596 142864 75638 142904
rect 75678 142864 75720 142904
rect 75392 142855 75760 142864
rect 74152 142148 74520 142157
rect 74192 142108 74234 142148
rect 74274 142108 74316 142148
rect 74356 142108 74398 142148
rect 74438 142108 74480 142148
rect 74152 142099 74520 142108
rect 75392 141392 75760 141401
rect 75432 141352 75474 141392
rect 75514 141352 75556 141392
rect 75596 141352 75638 141392
rect 75678 141352 75720 141392
rect 75392 141343 75760 141352
rect 74152 140636 74520 140645
rect 74192 140596 74234 140636
rect 74274 140596 74316 140636
rect 74356 140596 74398 140636
rect 74438 140596 74480 140636
rect 74152 140587 74520 140596
rect 75392 139880 75760 139889
rect 75432 139840 75474 139880
rect 75514 139840 75556 139880
rect 75596 139840 75638 139880
rect 75678 139840 75720 139880
rect 75392 139831 75760 139840
rect 74152 139124 74520 139133
rect 74192 139084 74234 139124
rect 74274 139084 74316 139124
rect 74356 139084 74398 139124
rect 74438 139084 74480 139124
rect 74152 139075 74520 139084
rect 75392 138368 75760 138377
rect 75432 138328 75474 138368
rect 75514 138328 75556 138368
rect 75596 138328 75638 138368
rect 75678 138328 75720 138368
rect 75392 138319 75760 138328
rect 74152 137612 74520 137621
rect 74192 137572 74234 137612
rect 74274 137572 74316 137612
rect 74356 137572 74398 137612
rect 74438 137572 74480 137612
rect 74152 137563 74520 137572
rect 75392 136856 75760 136865
rect 75432 136816 75474 136856
rect 75514 136816 75556 136856
rect 75596 136816 75638 136856
rect 75678 136816 75720 136856
rect 75392 136807 75760 136816
rect 74152 136100 74520 136109
rect 74192 136060 74234 136100
rect 74274 136060 74316 136100
rect 74356 136060 74398 136100
rect 74438 136060 74480 136100
rect 74152 136051 74520 136060
rect 75392 135344 75760 135353
rect 75432 135304 75474 135344
rect 75514 135304 75556 135344
rect 75596 135304 75638 135344
rect 75678 135304 75720 135344
rect 75392 135295 75760 135304
rect 74152 134588 74520 134597
rect 74192 134548 74234 134588
rect 74274 134548 74316 134588
rect 74356 134548 74398 134588
rect 74438 134548 74480 134588
rect 74152 134539 74520 134548
rect 75392 133832 75760 133841
rect 75432 133792 75474 133832
rect 75514 133792 75556 133832
rect 75596 133792 75638 133832
rect 75678 133792 75720 133832
rect 75392 133783 75760 133792
rect 74152 133076 74520 133085
rect 74192 133036 74234 133076
rect 74274 133036 74316 133076
rect 74356 133036 74398 133076
rect 74438 133036 74480 133076
rect 74152 133027 74520 133036
rect 75392 132320 75760 132329
rect 75432 132280 75474 132320
rect 75514 132280 75556 132320
rect 75596 132280 75638 132320
rect 75678 132280 75720 132320
rect 75392 132271 75760 132280
rect 74152 131564 74520 131573
rect 74192 131524 74234 131564
rect 74274 131524 74316 131564
rect 74356 131524 74398 131564
rect 74438 131524 74480 131564
rect 74152 131515 74520 131524
rect 75392 130808 75760 130817
rect 75432 130768 75474 130808
rect 75514 130768 75556 130808
rect 75596 130768 75638 130808
rect 75678 130768 75720 130808
rect 75392 130759 75760 130768
rect 74152 130052 74520 130061
rect 74192 130012 74234 130052
rect 74274 130012 74316 130052
rect 74356 130012 74398 130052
rect 74438 130012 74480 130052
rect 74152 130003 74520 130012
rect 75392 129296 75760 129305
rect 75432 129256 75474 129296
rect 75514 129256 75556 129296
rect 75596 129256 75638 129296
rect 75678 129256 75720 129296
rect 75392 129247 75760 129256
rect 74152 128540 74520 128549
rect 74192 128500 74234 128540
rect 74274 128500 74316 128540
rect 74356 128500 74398 128540
rect 74438 128500 74480 128540
rect 74152 128491 74520 128500
rect 75392 127784 75760 127793
rect 75432 127744 75474 127784
rect 75514 127744 75556 127784
rect 75596 127744 75638 127784
rect 75678 127744 75720 127784
rect 75392 127735 75760 127744
rect 74152 127028 74520 127037
rect 74192 126988 74234 127028
rect 74274 126988 74316 127028
rect 74356 126988 74398 127028
rect 74438 126988 74480 127028
rect 74152 126979 74520 126988
rect 75392 126272 75760 126281
rect 75432 126232 75474 126272
rect 75514 126232 75556 126272
rect 75596 126232 75638 126272
rect 75678 126232 75720 126272
rect 75392 126223 75760 126232
rect 74152 125516 74520 125525
rect 74192 125476 74234 125516
rect 74274 125476 74316 125516
rect 74356 125476 74398 125516
rect 74438 125476 74480 125516
rect 74152 125467 74520 125476
rect 75392 124760 75760 124769
rect 75432 124720 75474 124760
rect 75514 124720 75556 124760
rect 75596 124720 75638 124760
rect 75678 124720 75720 124760
rect 75392 124711 75760 124720
rect 74152 124004 74520 124013
rect 74192 123964 74234 124004
rect 74274 123964 74316 124004
rect 74356 123964 74398 124004
rect 74438 123964 74480 124004
rect 74152 123955 74520 123964
rect 75392 123248 75760 123257
rect 75432 123208 75474 123248
rect 75514 123208 75556 123248
rect 75596 123208 75638 123248
rect 75678 123208 75720 123248
rect 75392 123199 75760 123208
rect 74152 122492 74520 122501
rect 74192 122452 74234 122492
rect 74274 122452 74316 122492
rect 74356 122452 74398 122492
rect 74438 122452 74480 122492
rect 74152 122443 74520 122452
rect 75392 121736 75760 121745
rect 75432 121696 75474 121736
rect 75514 121696 75556 121736
rect 75596 121696 75638 121736
rect 75678 121696 75720 121736
rect 75392 121687 75760 121696
rect 74152 120980 74520 120989
rect 74192 120940 74234 120980
rect 74274 120940 74316 120980
rect 74356 120940 74398 120980
rect 74438 120940 74480 120980
rect 74152 120931 74520 120940
rect 75392 120224 75760 120233
rect 75432 120184 75474 120224
rect 75514 120184 75556 120224
rect 75596 120184 75638 120224
rect 75678 120184 75720 120224
rect 75392 120175 75760 120184
rect 74152 119468 74520 119477
rect 74192 119428 74234 119468
rect 74274 119428 74316 119468
rect 74356 119428 74398 119468
rect 74438 119428 74480 119468
rect 74152 119419 74520 119428
rect 75392 118712 75760 118721
rect 75432 118672 75474 118712
rect 75514 118672 75556 118712
rect 75596 118672 75638 118712
rect 75678 118672 75720 118712
rect 75392 118663 75760 118672
rect 74152 117956 74520 117965
rect 74192 117916 74234 117956
rect 74274 117916 74316 117956
rect 74356 117916 74398 117956
rect 74438 117916 74480 117956
rect 74152 117907 74520 117916
rect 75392 117200 75760 117209
rect 75432 117160 75474 117200
rect 75514 117160 75556 117200
rect 75596 117160 75638 117200
rect 75678 117160 75720 117200
rect 75392 117151 75760 117160
rect 74152 116444 74520 116453
rect 74192 116404 74234 116444
rect 74274 116404 74316 116444
rect 74356 116404 74398 116444
rect 74438 116404 74480 116444
rect 74152 116395 74520 116404
rect 75392 115688 75760 115697
rect 75432 115648 75474 115688
rect 75514 115648 75556 115688
rect 75596 115648 75638 115688
rect 75678 115648 75720 115688
rect 75392 115639 75760 115648
rect 74152 114932 74520 114941
rect 74192 114892 74234 114932
rect 74274 114892 74316 114932
rect 74356 114892 74398 114932
rect 74438 114892 74480 114932
rect 74152 114883 74520 114892
rect 75392 114176 75760 114185
rect 75432 114136 75474 114176
rect 75514 114136 75556 114176
rect 75596 114136 75638 114176
rect 75678 114136 75720 114176
rect 75392 114127 75760 114136
rect 74152 113420 74520 113429
rect 74192 113380 74234 113420
rect 74274 113380 74316 113420
rect 74356 113380 74398 113420
rect 74438 113380 74480 113420
rect 74152 113371 74520 113380
rect 75392 112664 75760 112673
rect 75432 112624 75474 112664
rect 75514 112624 75556 112664
rect 75596 112624 75638 112664
rect 75678 112624 75720 112664
rect 75392 112615 75760 112624
rect 74152 111908 74520 111917
rect 74192 111868 74234 111908
rect 74274 111868 74316 111908
rect 74356 111868 74398 111908
rect 74438 111868 74480 111908
rect 74152 111859 74520 111868
rect 75392 111152 75760 111161
rect 75432 111112 75474 111152
rect 75514 111112 75556 111152
rect 75596 111112 75638 111152
rect 75678 111112 75720 111152
rect 75392 111103 75760 111112
rect 74152 110396 74520 110405
rect 74192 110356 74234 110396
rect 74274 110356 74316 110396
rect 74356 110356 74398 110396
rect 74438 110356 74480 110396
rect 74152 110347 74520 110356
rect 75392 109640 75760 109649
rect 75432 109600 75474 109640
rect 75514 109600 75556 109640
rect 75596 109600 75638 109640
rect 75678 109600 75720 109640
rect 75392 109591 75760 109600
rect 74152 108884 74520 108893
rect 74192 108844 74234 108884
rect 74274 108844 74316 108884
rect 74356 108844 74398 108884
rect 74438 108844 74480 108884
rect 74152 108835 74520 108844
rect 75392 108128 75760 108137
rect 75432 108088 75474 108128
rect 75514 108088 75556 108128
rect 75596 108088 75638 108128
rect 75678 108088 75720 108128
rect 75392 108079 75760 108088
rect 74152 107372 74520 107381
rect 74192 107332 74234 107372
rect 74274 107332 74316 107372
rect 74356 107332 74398 107372
rect 74438 107332 74480 107372
rect 74152 107323 74520 107332
rect 75392 106616 75760 106625
rect 75432 106576 75474 106616
rect 75514 106576 75556 106616
rect 75596 106576 75638 106616
rect 75678 106576 75720 106616
rect 75392 106567 75760 106576
rect 74152 105860 74520 105869
rect 74192 105820 74234 105860
rect 74274 105820 74316 105860
rect 74356 105820 74398 105860
rect 74438 105820 74480 105860
rect 74152 105811 74520 105820
rect 75392 105104 75760 105113
rect 75432 105064 75474 105104
rect 75514 105064 75556 105104
rect 75596 105064 75638 105104
rect 75678 105064 75720 105104
rect 75392 105055 75760 105064
rect 74152 104348 74520 104357
rect 74192 104308 74234 104348
rect 74274 104308 74316 104348
rect 74356 104308 74398 104348
rect 74438 104308 74480 104348
rect 74152 104299 74520 104308
rect 75392 103592 75760 103601
rect 75432 103552 75474 103592
rect 75514 103552 75556 103592
rect 75596 103552 75638 103592
rect 75678 103552 75720 103592
rect 75392 103543 75760 103552
rect 74152 102836 74520 102845
rect 74192 102796 74234 102836
rect 74274 102796 74316 102836
rect 74356 102796 74398 102836
rect 74438 102796 74480 102836
rect 74152 102787 74520 102796
rect 75392 102080 75760 102089
rect 75432 102040 75474 102080
rect 75514 102040 75556 102080
rect 75596 102040 75638 102080
rect 75678 102040 75720 102080
rect 75392 102031 75760 102040
rect 74152 101324 74520 101333
rect 74192 101284 74234 101324
rect 74274 101284 74316 101324
rect 74356 101284 74398 101324
rect 74438 101284 74480 101324
rect 74152 101275 74520 101284
rect 75392 100568 75760 100577
rect 75432 100528 75474 100568
rect 75514 100528 75556 100568
rect 75596 100528 75638 100568
rect 75678 100528 75720 100568
rect 75392 100519 75760 100528
rect 74152 99812 74520 99821
rect 74192 99772 74234 99812
rect 74274 99772 74316 99812
rect 74356 99772 74398 99812
rect 74438 99772 74480 99812
rect 74152 99763 74520 99772
rect 75392 99056 75760 99065
rect 75432 99016 75474 99056
rect 75514 99016 75556 99056
rect 75596 99016 75638 99056
rect 75678 99016 75720 99056
rect 75392 99007 75760 99016
rect 74152 98300 74520 98309
rect 74192 98260 74234 98300
rect 74274 98260 74316 98300
rect 74356 98260 74398 98300
rect 74438 98260 74480 98300
rect 74152 98251 74520 98260
rect 75392 97544 75760 97553
rect 75432 97504 75474 97544
rect 75514 97504 75556 97544
rect 75596 97504 75638 97544
rect 75678 97504 75720 97544
rect 75392 97495 75760 97504
rect 74152 96788 74520 96797
rect 74192 96748 74234 96788
rect 74274 96748 74316 96788
rect 74356 96748 74398 96788
rect 74438 96748 74480 96788
rect 74152 96739 74520 96748
rect 75392 96032 75760 96041
rect 75432 95992 75474 96032
rect 75514 95992 75556 96032
rect 75596 95992 75638 96032
rect 75678 95992 75720 96032
rect 75392 95983 75760 95992
rect 74152 95276 74520 95285
rect 74192 95236 74234 95276
rect 74274 95236 74316 95276
rect 74356 95236 74398 95276
rect 74438 95236 74480 95276
rect 74152 95227 74520 95236
rect 75392 94520 75760 94529
rect 75432 94480 75474 94520
rect 75514 94480 75556 94520
rect 75596 94480 75638 94520
rect 75678 94480 75720 94520
rect 75392 94471 75760 94480
rect 74152 93764 74520 93773
rect 74192 93724 74234 93764
rect 74274 93724 74316 93764
rect 74356 93724 74398 93764
rect 74438 93724 74480 93764
rect 74152 93715 74520 93724
rect 75392 93008 75760 93017
rect 75432 92968 75474 93008
rect 75514 92968 75556 93008
rect 75596 92968 75638 93008
rect 75678 92968 75720 93008
rect 75392 92959 75760 92968
rect 74152 92252 74520 92261
rect 74192 92212 74234 92252
rect 74274 92212 74316 92252
rect 74356 92212 74398 92252
rect 74438 92212 74480 92252
rect 74152 92203 74520 92212
rect 75392 91496 75760 91505
rect 75432 91456 75474 91496
rect 75514 91456 75556 91496
rect 75596 91456 75638 91496
rect 75678 91456 75720 91496
rect 75392 91447 75760 91456
rect 74152 90740 74520 90749
rect 74192 90700 74234 90740
rect 74274 90700 74316 90740
rect 74356 90700 74398 90740
rect 74438 90700 74480 90740
rect 74152 90691 74520 90700
rect 75392 89984 75760 89993
rect 75432 89944 75474 89984
rect 75514 89944 75556 89984
rect 75596 89944 75638 89984
rect 75678 89944 75720 89984
rect 75392 89935 75760 89944
rect 74152 89228 74520 89237
rect 74192 89188 74234 89228
rect 74274 89188 74316 89228
rect 74356 89188 74398 89228
rect 74438 89188 74480 89228
rect 74152 89179 74520 89188
rect 75392 88472 75760 88481
rect 75432 88432 75474 88472
rect 75514 88432 75556 88472
rect 75596 88432 75638 88472
rect 75678 88432 75720 88472
rect 75392 88423 75760 88432
rect 74152 87716 74520 87725
rect 74192 87676 74234 87716
rect 74274 87676 74316 87716
rect 74356 87676 74398 87716
rect 74438 87676 74480 87716
rect 74152 87667 74520 87676
rect 75392 86960 75760 86969
rect 75432 86920 75474 86960
rect 75514 86920 75556 86960
rect 75596 86920 75638 86960
rect 75678 86920 75720 86960
rect 75392 86911 75760 86920
rect 74152 86204 74520 86213
rect 74192 86164 74234 86204
rect 74274 86164 74316 86204
rect 74356 86164 74398 86204
rect 74438 86164 74480 86204
rect 74152 86155 74520 86164
rect 75392 85448 75760 85457
rect 75432 85408 75474 85448
rect 75514 85408 75556 85448
rect 75596 85408 75638 85448
rect 75678 85408 75720 85448
rect 75392 85399 75760 85408
rect 74152 84692 74520 84701
rect 74192 84652 74234 84692
rect 74274 84652 74316 84692
rect 74356 84652 74398 84692
rect 74438 84652 74480 84692
rect 74152 84643 74520 84652
rect 75392 83936 75760 83945
rect 75432 83896 75474 83936
rect 75514 83896 75556 83936
rect 75596 83896 75638 83936
rect 75678 83896 75720 83936
rect 75392 83887 75760 83896
rect 74152 83180 74520 83189
rect 74192 83140 74234 83180
rect 74274 83140 74316 83180
rect 74356 83140 74398 83180
rect 74438 83140 74480 83180
rect 74152 83131 74520 83140
rect 75392 82424 75760 82433
rect 75432 82384 75474 82424
rect 75514 82384 75556 82424
rect 75596 82384 75638 82424
rect 75678 82384 75720 82424
rect 75392 82375 75760 82384
rect 74152 81668 74520 81677
rect 74192 81628 74234 81668
rect 74274 81628 74316 81668
rect 74356 81628 74398 81668
rect 74438 81628 74480 81668
rect 74152 81619 74520 81628
rect 75392 80912 75760 80921
rect 75432 80872 75474 80912
rect 75514 80872 75556 80912
rect 75596 80872 75638 80912
rect 75678 80872 75720 80912
rect 75392 80863 75760 80872
rect 74152 80156 74520 80165
rect 74192 80116 74234 80156
rect 74274 80116 74316 80156
rect 74356 80116 74398 80156
rect 74438 80116 74480 80156
rect 74152 80107 74520 80116
rect 75392 79400 75760 79409
rect 75432 79360 75474 79400
rect 75514 79360 75556 79400
rect 75596 79360 75638 79400
rect 75678 79360 75720 79400
rect 75392 79351 75760 79360
rect 74152 78644 74520 78653
rect 74192 78604 74234 78644
rect 74274 78604 74316 78644
rect 74356 78604 74398 78644
rect 74438 78604 74480 78644
rect 74152 78595 74520 78604
rect 75392 77888 75760 77897
rect 75432 77848 75474 77888
rect 75514 77848 75556 77888
rect 75596 77848 75638 77888
rect 75678 77848 75720 77888
rect 75392 77839 75760 77848
rect 74152 77132 74520 77141
rect 74192 77092 74234 77132
rect 74274 77092 74316 77132
rect 74356 77092 74398 77132
rect 74438 77092 74480 77132
rect 74152 77083 74520 77092
rect 75392 76376 75760 76385
rect 75432 76336 75474 76376
rect 75514 76336 75556 76376
rect 75596 76336 75638 76376
rect 75678 76336 75720 76376
rect 75392 76327 75760 76336
rect 74152 75620 74520 75629
rect 74192 75580 74234 75620
rect 74274 75580 74316 75620
rect 74356 75580 74398 75620
rect 74438 75580 74480 75620
rect 74152 75571 74520 75580
rect 75392 74864 75760 74873
rect 75432 74824 75474 74864
rect 75514 74824 75556 74864
rect 75596 74824 75638 74864
rect 75678 74824 75720 74864
rect 75392 74815 75760 74824
rect 74152 74108 74520 74117
rect 74192 74068 74234 74108
rect 74274 74068 74316 74108
rect 74356 74068 74398 74108
rect 74438 74068 74480 74108
rect 74152 74059 74520 74068
rect 75392 73352 75760 73361
rect 75432 73312 75474 73352
rect 75514 73312 75556 73352
rect 75596 73312 75638 73352
rect 75678 73312 75720 73352
rect 75392 73303 75760 73312
rect 74152 72596 74520 72605
rect 74192 72556 74234 72596
rect 74274 72556 74316 72596
rect 74356 72556 74398 72596
rect 74438 72556 74480 72596
rect 74152 72547 74520 72556
rect 75392 71840 75760 71849
rect 75432 71800 75474 71840
rect 75514 71800 75556 71840
rect 75596 71800 75638 71840
rect 75678 71800 75720 71840
rect 75392 71791 75760 71800
rect 88012 64364 88052 159319
rect 90512 151976 90880 151985
rect 90552 151936 90594 151976
rect 90634 151936 90676 151976
rect 90716 151936 90758 151976
rect 90798 151936 90840 151976
rect 90512 151927 90880 151936
rect 89272 151220 89640 151229
rect 89312 151180 89354 151220
rect 89394 151180 89436 151220
rect 89476 151180 89518 151220
rect 89558 151180 89600 151220
rect 89272 151171 89640 151180
rect 90512 150464 90880 150473
rect 90552 150424 90594 150464
rect 90634 150424 90676 150464
rect 90716 150424 90758 150464
rect 90798 150424 90840 150464
rect 90512 150415 90880 150424
rect 89272 149708 89640 149717
rect 89312 149668 89354 149708
rect 89394 149668 89436 149708
rect 89476 149668 89518 149708
rect 89558 149668 89600 149708
rect 89272 149659 89640 149668
rect 90512 148952 90880 148961
rect 90552 148912 90594 148952
rect 90634 148912 90676 148952
rect 90716 148912 90758 148952
rect 90798 148912 90840 148952
rect 90512 148903 90880 148912
rect 89272 148196 89640 148205
rect 89312 148156 89354 148196
rect 89394 148156 89436 148196
rect 89476 148156 89518 148196
rect 89558 148156 89600 148196
rect 89272 148147 89640 148156
rect 90512 147440 90880 147449
rect 90552 147400 90594 147440
rect 90634 147400 90676 147440
rect 90716 147400 90758 147440
rect 90798 147400 90840 147440
rect 90512 147391 90880 147400
rect 89272 146684 89640 146693
rect 89312 146644 89354 146684
rect 89394 146644 89436 146684
rect 89476 146644 89518 146684
rect 89558 146644 89600 146684
rect 89272 146635 89640 146644
rect 90512 145928 90880 145937
rect 90552 145888 90594 145928
rect 90634 145888 90676 145928
rect 90716 145888 90758 145928
rect 90798 145888 90840 145928
rect 90512 145879 90880 145888
rect 89272 145172 89640 145181
rect 89312 145132 89354 145172
rect 89394 145132 89436 145172
rect 89476 145132 89518 145172
rect 89558 145132 89600 145172
rect 89272 145123 89640 145132
rect 90512 144416 90880 144425
rect 90552 144376 90594 144416
rect 90634 144376 90676 144416
rect 90716 144376 90758 144416
rect 90798 144376 90840 144416
rect 90512 144367 90880 144376
rect 89272 143660 89640 143669
rect 89312 143620 89354 143660
rect 89394 143620 89436 143660
rect 89476 143620 89518 143660
rect 89558 143620 89600 143660
rect 89272 143611 89640 143620
rect 90512 142904 90880 142913
rect 90552 142864 90594 142904
rect 90634 142864 90676 142904
rect 90716 142864 90758 142904
rect 90798 142864 90840 142904
rect 90512 142855 90880 142864
rect 89272 142148 89640 142157
rect 89312 142108 89354 142148
rect 89394 142108 89436 142148
rect 89476 142108 89518 142148
rect 89558 142108 89600 142148
rect 89272 142099 89640 142108
rect 90512 141392 90880 141401
rect 90552 141352 90594 141392
rect 90634 141352 90676 141392
rect 90716 141352 90758 141392
rect 90798 141352 90840 141392
rect 90512 141343 90880 141352
rect 89272 140636 89640 140645
rect 89312 140596 89354 140636
rect 89394 140596 89436 140636
rect 89476 140596 89518 140636
rect 89558 140596 89600 140636
rect 89272 140587 89640 140596
rect 90512 139880 90880 139889
rect 90552 139840 90594 139880
rect 90634 139840 90676 139880
rect 90716 139840 90758 139880
rect 90798 139840 90840 139880
rect 90512 139831 90880 139840
rect 89272 139124 89640 139133
rect 89312 139084 89354 139124
rect 89394 139084 89436 139124
rect 89476 139084 89518 139124
rect 89558 139084 89600 139124
rect 89272 139075 89640 139084
rect 90512 138368 90880 138377
rect 90552 138328 90594 138368
rect 90634 138328 90676 138368
rect 90716 138328 90758 138368
rect 90798 138328 90840 138368
rect 90512 138319 90880 138328
rect 89272 137612 89640 137621
rect 89312 137572 89354 137612
rect 89394 137572 89436 137612
rect 89476 137572 89518 137612
rect 89558 137572 89600 137612
rect 89272 137563 89640 137572
rect 90512 136856 90880 136865
rect 90552 136816 90594 136856
rect 90634 136816 90676 136856
rect 90716 136816 90758 136856
rect 90798 136816 90840 136856
rect 90512 136807 90880 136816
rect 89272 136100 89640 136109
rect 89312 136060 89354 136100
rect 89394 136060 89436 136100
rect 89476 136060 89518 136100
rect 89558 136060 89600 136100
rect 89272 136051 89640 136060
rect 90512 135344 90880 135353
rect 90552 135304 90594 135344
rect 90634 135304 90676 135344
rect 90716 135304 90758 135344
rect 90798 135304 90840 135344
rect 90512 135295 90880 135304
rect 89272 134588 89640 134597
rect 89312 134548 89354 134588
rect 89394 134548 89436 134588
rect 89476 134548 89518 134588
rect 89558 134548 89600 134588
rect 89272 134539 89640 134548
rect 90512 133832 90880 133841
rect 90552 133792 90594 133832
rect 90634 133792 90676 133832
rect 90716 133792 90758 133832
rect 90798 133792 90840 133832
rect 90512 133783 90880 133792
rect 89272 133076 89640 133085
rect 89312 133036 89354 133076
rect 89394 133036 89436 133076
rect 89476 133036 89518 133076
rect 89558 133036 89600 133076
rect 89272 133027 89640 133036
rect 90512 132320 90880 132329
rect 90552 132280 90594 132320
rect 90634 132280 90676 132320
rect 90716 132280 90758 132320
rect 90798 132280 90840 132320
rect 90512 132271 90880 132280
rect 89272 131564 89640 131573
rect 89312 131524 89354 131564
rect 89394 131524 89436 131564
rect 89476 131524 89518 131564
rect 89558 131524 89600 131564
rect 89272 131515 89640 131524
rect 90512 130808 90880 130817
rect 90552 130768 90594 130808
rect 90634 130768 90676 130808
rect 90716 130768 90758 130808
rect 90798 130768 90840 130808
rect 90512 130759 90880 130768
rect 89272 130052 89640 130061
rect 89312 130012 89354 130052
rect 89394 130012 89436 130052
rect 89476 130012 89518 130052
rect 89558 130012 89600 130052
rect 89272 130003 89640 130012
rect 90512 129296 90880 129305
rect 90552 129256 90594 129296
rect 90634 129256 90676 129296
rect 90716 129256 90758 129296
rect 90798 129256 90840 129296
rect 90512 129247 90880 129256
rect 89272 128540 89640 128549
rect 89312 128500 89354 128540
rect 89394 128500 89436 128540
rect 89476 128500 89518 128540
rect 89558 128500 89600 128540
rect 89272 128491 89640 128500
rect 90512 127784 90880 127793
rect 90552 127744 90594 127784
rect 90634 127744 90676 127784
rect 90716 127744 90758 127784
rect 90798 127744 90840 127784
rect 90512 127735 90880 127744
rect 89272 127028 89640 127037
rect 89312 126988 89354 127028
rect 89394 126988 89436 127028
rect 89476 126988 89518 127028
rect 89558 126988 89600 127028
rect 89272 126979 89640 126988
rect 90512 126272 90880 126281
rect 90552 126232 90594 126272
rect 90634 126232 90676 126272
rect 90716 126232 90758 126272
rect 90798 126232 90840 126272
rect 90512 126223 90880 126232
rect 89272 125516 89640 125525
rect 89312 125476 89354 125516
rect 89394 125476 89436 125516
rect 89476 125476 89518 125516
rect 89558 125476 89600 125516
rect 89272 125467 89640 125476
rect 90512 124760 90880 124769
rect 90552 124720 90594 124760
rect 90634 124720 90676 124760
rect 90716 124720 90758 124760
rect 90798 124720 90840 124760
rect 90512 124711 90880 124720
rect 89272 124004 89640 124013
rect 89312 123964 89354 124004
rect 89394 123964 89436 124004
rect 89476 123964 89518 124004
rect 89558 123964 89600 124004
rect 89272 123955 89640 123964
rect 90512 123248 90880 123257
rect 90552 123208 90594 123248
rect 90634 123208 90676 123248
rect 90716 123208 90758 123248
rect 90798 123208 90840 123248
rect 90512 123199 90880 123208
rect 89272 122492 89640 122501
rect 89312 122452 89354 122492
rect 89394 122452 89436 122492
rect 89476 122452 89518 122492
rect 89558 122452 89600 122492
rect 89272 122443 89640 122452
rect 90512 121736 90880 121745
rect 90552 121696 90594 121736
rect 90634 121696 90676 121736
rect 90716 121696 90758 121736
rect 90798 121696 90840 121736
rect 90512 121687 90880 121696
rect 89272 120980 89640 120989
rect 89312 120940 89354 120980
rect 89394 120940 89436 120980
rect 89476 120940 89518 120980
rect 89558 120940 89600 120980
rect 89272 120931 89640 120940
rect 90512 120224 90880 120233
rect 90552 120184 90594 120224
rect 90634 120184 90676 120224
rect 90716 120184 90758 120224
rect 90798 120184 90840 120224
rect 90512 120175 90880 120184
rect 89272 119468 89640 119477
rect 89312 119428 89354 119468
rect 89394 119428 89436 119468
rect 89476 119428 89518 119468
rect 89558 119428 89600 119468
rect 89272 119419 89640 119428
rect 90512 118712 90880 118721
rect 90552 118672 90594 118712
rect 90634 118672 90676 118712
rect 90716 118672 90758 118712
rect 90798 118672 90840 118712
rect 90512 118663 90880 118672
rect 89272 117956 89640 117965
rect 89312 117916 89354 117956
rect 89394 117916 89436 117956
rect 89476 117916 89518 117956
rect 89558 117916 89600 117956
rect 89272 117907 89640 117916
rect 90512 117200 90880 117209
rect 90552 117160 90594 117200
rect 90634 117160 90676 117200
rect 90716 117160 90758 117200
rect 90798 117160 90840 117200
rect 90512 117151 90880 117160
rect 89272 116444 89640 116453
rect 89312 116404 89354 116444
rect 89394 116404 89436 116444
rect 89476 116404 89518 116444
rect 89558 116404 89600 116444
rect 89272 116395 89640 116404
rect 90512 115688 90880 115697
rect 90552 115648 90594 115688
rect 90634 115648 90676 115688
rect 90716 115648 90758 115688
rect 90798 115648 90840 115688
rect 90512 115639 90880 115648
rect 89272 114932 89640 114941
rect 89312 114892 89354 114932
rect 89394 114892 89436 114932
rect 89476 114892 89518 114932
rect 89558 114892 89600 114932
rect 89272 114883 89640 114892
rect 90512 114176 90880 114185
rect 90552 114136 90594 114176
rect 90634 114136 90676 114176
rect 90716 114136 90758 114176
rect 90798 114136 90840 114176
rect 90512 114127 90880 114136
rect 89272 113420 89640 113429
rect 89312 113380 89354 113420
rect 89394 113380 89436 113420
rect 89476 113380 89518 113420
rect 89558 113380 89600 113420
rect 89272 113371 89640 113380
rect 90512 112664 90880 112673
rect 90552 112624 90594 112664
rect 90634 112624 90676 112664
rect 90716 112624 90758 112664
rect 90798 112624 90840 112664
rect 90512 112615 90880 112624
rect 89272 111908 89640 111917
rect 89312 111868 89354 111908
rect 89394 111868 89436 111908
rect 89476 111868 89518 111908
rect 89558 111868 89600 111908
rect 89272 111859 89640 111868
rect 90512 111152 90880 111161
rect 90552 111112 90594 111152
rect 90634 111112 90676 111152
rect 90716 111112 90758 111152
rect 90798 111112 90840 111152
rect 90512 111103 90880 111112
rect 89272 110396 89640 110405
rect 89312 110356 89354 110396
rect 89394 110356 89436 110396
rect 89476 110356 89518 110396
rect 89558 110356 89600 110396
rect 89272 110347 89640 110356
rect 90512 109640 90880 109649
rect 90552 109600 90594 109640
rect 90634 109600 90676 109640
rect 90716 109600 90758 109640
rect 90798 109600 90840 109640
rect 90512 109591 90880 109600
rect 89272 108884 89640 108893
rect 89312 108844 89354 108884
rect 89394 108844 89436 108884
rect 89476 108844 89518 108884
rect 89558 108844 89600 108884
rect 89272 108835 89640 108844
rect 90512 108128 90880 108137
rect 90552 108088 90594 108128
rect 90634 108088 90676 108128
rect 90716 108088 90758 108128
rect 90798 108088 90840 108128
rect 90512 108079 90880 108088
rect 89272 107372 89640 107381
rect 89312 107332 89354 107372
rect 89394 107332 89436 107372
rect 89476 107332 89518 107372
rect 89558 107332 89600 107372
rect 89272 107323 89640 107332
rect 90512 106616 90880 106625
rect 90552 106576 90594 106616
rect 90634 106576 90676 106616
rect 90716 106576 90758 106616
rect 90798 106576 90840 106616
rect 90512 106567 90880 106576
rect 89272 105860 89640 105869
rect 89312 105820 89354 105860
rect 89394 105820 89436 105860
rect 89476 105820 89518 105860
rect 89558 105820 89600 105860
rect 89272 105811 89640 105820
rect 90512 105104 90880 105113
rect 90552 105064 90594 105104
rect 90634 105064 90676 105104
rect 90716 105064 90758 105104
rect 90798 105064 90840 105104
rect 90512 105055 90880 105064
rect 89272 104348 89640 104357
rect 89312 104308 89354 104348
rect 89394 104308 89436 104348
rect 89476 104308 89518 104348
rect 89558 104308 89600 104348
rect 89272 104299 89640 104308
rect 90512 103592 90880 103601
rect 90552 103552 90594 103592
rect 90634 103552 90676 103592
rect 90716 103552 90758 103592
rect 90798 103552 90840 103592
rect 90512 103543 90880 103552
rect 89272 102836 89640 102845
rect 89312 102796 89354 102836
rect 89394 102796 89436 102836
rect 89476 102796 89518 102836
rect 89558 102796 89600 102836
rect 89272 102787 89640 102796
rect 90512 102080 90880 102089
rect 90552 102040 90594 102080
rect 90634 102040 90676 102080
rect 90716 102040 90758 102080
rect 90798 102040 90840 102080
rect 90512 102031 90880 102040
rect 89272 101324 89640 101333
rect 89312 101284 89354 101324
rect 89394 101284 89436 101324
rect 89476 101284 89518 101324
rect 89558 101284 89600 101324
rect 89272 101275 89640 101284
rect 90512 100568 90880 100577
rect 90552 100528 90594 100568
rect 90634 100528 90676 100568
rect 90716 100528 90758 100568
rect 90798 100528 90840 100568
rect 90512 100519 90880 100528
rect 89272 99812 89640 99821
rect 89312 99772 89354 99812
rect 89394 99772 89436 99812
rect 89476 99772 89518 99812
rect 89558 99772 89600 99812
rect 89272 99763 89640 99772
rect 90512 99056 90880 99065
rect 90552 99016 90594 99056
rect 90634 99016 90676 99056
rect 90716 99016 90758 99056
rect 90798 99016 90840 99056
rect 90512 99007 90880 99016
rect 89272 98300 89640 98309
rect 89312 98260 89354 98300
rect 89394 98260 89436 98300
rect 89476 98260 89518 98300
rect 89558 98260 89600 98300
rect 89272 98251 89640 98260
rect 90512 97544 90880 97553
rect 90552 97504 90594 97544
rect 90634 97504 90676 97544
rect 90716 97504 90758 97544
rect 90798 97504 90840 97544
rect 90512 97495 90880 97504
rect 89272 96788 89640 96797
rect 89312 96748 89354 96788
rect 89394 96748 89436 96788
rect 89476 96748 89518 96788
rect 89558 96748 89600 96788
rect 89272 96739 89640 96748
rect 90512 96032 90880 96041
rect 90552 95992 90594 96032
rect 90634 95992 90676 96032
rect 90716 95992 90758 96032
rect 90798 95992 90840 96032
rect 90512 95983 90880 95992
rect 89272 95276 89640 95285
rect 89312 95236 89354 95276
rect 89394 95236 89436 95276
rect 89476 95236 89518 95276
rect 89558 95236 89600 95276
rect 89272 95227 89640 95236
rect 90512 94520 90880 94529
rect 90552 94480 90594 94520
rect 90634 94480 90676 94520
rect 90716 94480 90758 94520
rect 90798 94480 90840 94520
rect 90512 94471 90880 94480
rect 89272 93764 89640 93773
rect 89312 93724 89354 93764
rect 89394 93724 89436 93764
rect 89476 93724 89518 93764
rect 89558 93724 89600 93764
rect 89272 93715 89640 93724
rect 90512 93008 90880 93017
rect 90552 92968 90594 93008
rect 90634 92968 90676 93008
rect 90716 92968 90758 93008
rect 90798 92968 90840 93008
rect 90512 92959 90880 92968
rect 89272 92252 89640 92261
rect 89312 92212 89354 92252
rect 89394 92212 89436 92252
rect 89476 92212 89518 92252
rect 89558 92212 89600 92252
rect 89272 92203 89640 92212
rect 90512 91496 90880 91505
rect 90552 91456 90594 91496
rect 90634 91456 90676 91496
rect 90716 91456 90758 91496
rect 90798 91456 90840 91496
rect 90512 91447 90880 91456
rect 89272 90740 89640 90749
rect 89312 90700 89354 90740
rect 89394 90700 89436 90740
rect 89476 90700 89518 90740
rect 89558 90700 89600 90740
rect 89272 90691 89640 90700
rect 90512 89984 90880 89993
rect 90552 89944 90594 89984
rect 90634 89944 90676 89984
rect 90716 89944 90758 89984
rect 90798 89944 90840 89984
rect 90512 89935 90880 89944
rect 89272 89228 89640 89237
rect 89312 89188 89354 89228
rect 89394 89188 89436 89228
rect 89476 89188 89518 89228
rect 89558 89188 89600 89228
rect 89272 89179 89640 89188
rect 90512 88472 90880 88481
rect 90552 88432 90594 88472
rect 90634 88432 90676 88472
rect 90716 88432 90758 88472
rect 90798 88432 90840 88472
rect 90512 88423 90880 88432
rect 89272 87716 89640 87725
rect 89312 87676 89354 87716
rect 89394 87676 89436 87716
rect 89476 87676 89518 87716
rect 89558 87676 89600 87716
rect 89272 87667 89640 87676
rect 90512 86960 90880 86969
rect 90552 86920 90594 86960
rect 90634 86920 90676 86960
rect 90716 86920 90758 86960
rect 90798 86920 90840 86960
rect 90512 86911 90880 86920
rect 89272 86204 89640 86213
rect 89312 86164 89354 86204
rect 89394 86164 89436 86204
rect 89476 86164 89518 86204
rect 89558 86164 89600 86204
rect 89272 86155 89640 86164
rect 90512 85448 90880 85457
rect 90552 85408 90594 85448
rect 90634 85408 90676 85448
rect 90716 85408 90758 85448
rect 90798 85408 90840 85448
rect 90512 85399 90880 85408
rect 89272 84692 89640 84701
rect 89312 84652 89354 84692
rect 89394 84652 89436 84692
rect 89476 84652 89518 84692
rect 89558 84652 89600 84692
rect 89272 84643 89640 84652
rect 90512 83936 90880 83945
rect 90552 83896 90594 83936
rect 90634 83896 90676 83936
rect 90716 83896 90758 83936
rect 90798 83896 90840 83936
rect 90512 83887 90880 83896
rect 89272 83180 89640 83189
rect 89312 83140 89354 83180
rect 89394 83140 89436 83180
rect 89476 83140 89518 83180
rect 89558 83140 89600 83180
rect 89272 83131 89640 83140
rect 90512 82424 90880 82433
rect 90552 82384 90594 82424
rect 90634 82384 90676 82424
rect 90716 82384 90758 82424
rect 90798 82384 90840 82424
rect 90512 82375 90880 82384
rect 89272 81668 89640 81677
rect 89312 81628 89354 81668
rect 89394 81628 89436 81668
rect 89476 81628 89518 81668
rect 89558 81628 89600 81668
rect 89272 81619 89640 81628
rect 90512 80912 90880 80921
rect 90552 80872 90594 80912
rect 90634 80872 90676 80912
rect 90716 80872 90758 80912
rect 90798 80872 90840 80912
rect 90512 80863 90880 80872
rect 89272 80156 89640 80165
rect 89312 80116 89354 80156
rect 89394 80116 89436 80156
rect 89476 80116 89518 80156
rect 89558 80116 89600 80156
rect 89272 80107 89640 80116
rect 90512 79400 90880 79409
rect 90552 79360 90594 79400
rect 90634 79360 90676 79400
rect 90716 79360 90758 79400
rect 90798 79360 90840 79400
rect 90512 79351 90880 79360
rect 89272 78644 89640 78653
rect 89312 78604 89354 78644
rect 89394 78604 89436 78644
rect 89476 78604 89518 78644
rect 89558 78604 89600 78644
rect 89272 78595 89640 78604
rect 90512 77888 90880 77897
rect 90552 77848 90594 77888
rect 90634 77848 90676 77888
rect 90716 77848 90758 77888
rect 90798 77848 90840 77888
rect 90512 77839 90880 77848
rect 89272 77132 89640 77141
rect 89312 77092 89354 77132
rect 89394 77092 89436 77132
rect 89476 77092 89518 77132
rect 89558 77092 89600 77132
rect 89272 77083 89640 77092
rect 90512 76376 90880 76385
rect 90552 76336 90594 76376
rect 90634 76336 90676 76376
rect 90716 76336 90758 76376
rect 90798 76336 90840 76376
rect 90512 76327 90880 76336
rect 89272 75620 89640 75629
rect 89312 75580 89354 75620
rect 89394 75580 89436 75620
rect 89476 75580 89518 75620
rect 89558 75580 89600 75620
rect 89272 75571 89640 75580
rect 90512 74864 90880 74873
rect 90552 74824 90594 74864
rect 90634 74824 90676 74864
rect 90716 74824 90758 74864
rect 90798 74824 90840 74864
rect 90512 74815 90880 74824
rect 89272 74108 89640 74117
rect 89312 74068 89354 74108
rect 89394 74068 89436 74108
rect 89476 74068 89518 74108
rect 89558 74068 89600 74108
rect 89272 74059 89640 74068
rect 90512 73352 90880 73361
rect 90552 73312 90594 73352
rect 90634 73312 90676 73352
rect 90716 73312 90758 73352
rect 90798 73312 90840 73352
rect 90512 73303 90880 73312
rect 89272 72596 89640 72605
rect 89312 72556 89354 72596
rect 89394 72556 89436 72596
rect 89476 72556 89518 72596
rect 89558 72556 89600 72596
rect 89272 72547 89640 72556
rect 90512 71840 90880 71849
rect 90552 71800 90594 71840
rect 90634 71800 90676 71840
rect 90716 71800 90758 71840
rect 90798 71800 90840 71840
rect 90512 71791 90880 71800
rect 104044 64364 104084 159403
rect 119692 159377 119732 160020
rect 135724 159461 135764 160020
rect 135723 159452 135765 159461
rect 135723 159412 135724 159452
rect 135764 159412 135765 159452
rect 135723 159403 135765 159412
rect 119691 159368 119733 159377
rect 119691 159328 119692 159368
rect 119732 159328 119733 159368
rect 119691 159319 119733 159328
rect 151660 158780 151700 160020
rect 151564 158740 151700 158780
rect 105632 151976 106000 151985
rect 105672 151936 105714 151976
rect 105754 151936 105796 151976
rect 105836 151936 105878 151976
rect 105918 151936 105960 151976
rect 105632 151927 106000 151936
rect 120752 151976 121120 151985
rect 120792 151936 120834 151976
rect 120874 151936 120916 151976
rect 120956 151936 120998 151976
rect 121038 151936 121080 151976
rect 120752 151927 121120 151936
rect 135872 151976 136240 151985
rect 135912 151936 135954 151976
rect 135994 151936 136036 151976
rect 136076 151936 136118 151976
rect 136158 151936 136200 151976
rect 135872 151927 136240 151936
rect 150992 151976 151360 151985
rect 151032 151936 151074 151976
rect 151114 151936 151156 151976
rect 151196 151936 151238 151976
rect 151278 151936 151320 151976
rect 150992 151927 151360 151936
rect 104392 151220 104760 151229
rect 104432 151180 104474 151220
rect 104514 151180 104556 151220
rect 104596 151180 104638 151220
rect 104678 151180 104720 151220
rect 104392 151171 104760 151180
rect 119512 151220 119880 151229
rect 119552 151180 119594 151220
rect 119634 151180 119676 151220
rect 119716 151180 119758 151220
rect 119798 151180 119840 151220
rect 119512 151171 119880 151180
rect 134632 151220 135000 151229
rect 134672 151180 134714 151220
rect 134754 151180 134796 151220
rect 134836 151180 134878 151220
rect 134918 151180 134960 151220
rect 134632 151171 135000 151180
rect 149752 151220 150120 151229
rect 149792 151180 149834 151220
rect 149874 151180 149916 151220
rect 149956 151180 149998 151220
rect 150038 151180 150080 151220
rect 149752 151171 150120 151180
rect 105632 150464 106000 150473
rect 105672 150424 105714 150464
rect 105754 150424 105796 150464
rect 105836 150424 105878 150464
rect 105918 150424 105960 150464
rect 105632 150415 106000 150424
rect 120752 150464 121120 150473
rect 120792 150424 120834 150464
rect 120874 150424 120916 150464
rect 120956 150424 120998 150464
rect 121038 150424 121080 150464
rect 120752 150415 121120 150424
rect 135872 150464 136240 150473
rect 135912 150424 135954 150464
rect 135994 150424 136036 150464
rect 136076 150424 136118 150464
rect 136158 150424 136200 150464
rect 135872 150415 136240 150424
rect 150992 150464 151360 150473
rect 151032 150424 151074 150464
rect 151114 150424 151156 150464
rect 151196 150424 151238 150464
rect 151278 150424 151320 150464
rect 150992 150415 151360 150424
rect 104392 149708 104760 149717
rect 104432 149668 104474 149708
rect 104514 149668 104556 149708
rect 104596 149668 104638 149708
rect 104678 149668 104720 149708
rect 104392 149659 104760 149668
rect 119512 149708 119880 149717
rect 119552 149668 119594 149708
rect 119634 149668 119676 149708
rect 119716 149668 119758 149708
rect 119798 149668 119840 149708
rect 119512 149659 119880 149668
rect 134632 149708 135000 149717
rect 134672 149668 134714 149708
rect 134754 149668 134796 149708
rect 134836 149668 134878 149708
rect 134918 149668 134960 149708
rect 134632 149659 135000 149668
rect 149752 149708 150120 149717
rect 149792 149668 149834 149708
rect 149874 149668 149916 149708
rect 149956 149668 149998 149708
rect 150038 149668 150080 149708
rect 149752 149659 150120 149668
rect 105632 148952 106000 148961
rect 105672 148912 105714 148952
rect 105754 148912 105796 148952
rect 105836 148912 105878 148952
rect 105918 148912 105960 148952
rect 105632 148903 106000 148912
rect 120752 148952 121120 148961
rect 120792 148912 120834 148952
rect 120874 148912 120916 148952
rect 120956 148912 120998 148952
rect 121038 148912 121080 148952
rect 120752 148903 121120 148912
rect 135872 148952 136240 148961
rect 135912 148912 135954 148952
rect 135994 148912 136036 148952
rect 136076 148912 136118 148952
rect 136158 148912 136200 148952
rect 135872 148903 136240 148912
rect 150992 148952 151360 148961
rect 151032 148912 151074 148952
rect 151114 148912 151156 148952
rect 151196 148912 151238 148952
rect 151278 148912 151320 148952
rect 150992 148903 151360 148912
rect 104392 148196 104760 148205
rect 104432 148156 104474 148196
rect 104514 148156 104556 148196
rect 104596 148156 104638 148196
rect 104678 148156 104720 148196
rect 104392 148147 104760 148156
rect 119512 148196 119880 148205
rect 119552 148156 119594 148196
rect 119634 148156 119676 148196
rect 119716 148156 119758 148196
rect 119798 148156 119840 148196
rect 119512 148147 119880 148156
rect 134632 148196 135000 148205
rect 134672 148156 134714 148196
rect 134754 148156 134796 148196
rect 134836 148156 134878 148196
rect 134918 148156 134960 148196
rect 134632 148147 135000 148156
rect 149752 148196 150120 148205
rect 149792 148156 149834 148196
rect 149874 148156 149916 148196
rect 149956 148156 149998 148196
rect 150038 148156 150080 148196
rect 149752 148147 150120 148156
rect 105632 147440 106000 147449
rect 105672 147400 105714 147440
rect 105754 147400 105796 147440
rect 105836 147400 105878 147440
rect 105918 147400 105960 147440
rect 105632 147391 106000 147400
rect 120752 147440 121120 147449
rect 120792 147400 120834 147440
rect 120874 147400 120916 147440
rect 120956 147400 120998 147440
rect 121038 147400 121080 147440
rect 120752 147391 121120 147400
rect 135872 147440 136240 147449
rect 135912 147400 135954 147440
rect 135994 147400 136036 147440
rect 136076 147400 136118 147440
rect 136158 147400 136200 147440
rect 135872 147391 136240 147400
rect 150992 147440 151360 147449
rect 151032 147400 151074 147440
rect 151114 147400 151156 147440
rect 151196 147400 151238 147440
rect 151278 147400 151320 147440
rect 150992 147391 151360 147400
rect 104392 146684 104760 146693
rect 104432 146644 104474 146684
rect 104514 146644 104556 146684
rect 104596 146644 104638 146684
rect 104678 146644 104720 146684
rect 104392 146635 104760 146644
rect 119512 146684 119880 146693
rect 119552 146644 119594 146684
rect 119634 146644 119676 146684
rect 119716 146644 119758 146684
rect 119798 146644 119840 146684
rect 119512 146635 119880 146644
rect 134632 146684 135000 146693
rect 134672 146644 134714 146684
rect 134754 146644 134796 146684
rect 134836 146644 134878 146684
rect 134918 146644 134960 146684
rect 134632 146635 135000 146644
rect 149752 146684 150120 146693
rect 149792 146644 149834 146684
rect 149874 146644 149916 146684
rect 149956 146644 149998 146684
rect 150038 146644 150080 146684
rect 149752 146635 150120 146644
rect 105632 145928 106000 145937
rect 105672 145888 105714 145928
rect 105754 145888 105796 145928
rect 105836 145888 105878 145928
rect 105918 145888 105960 145928
rect 105632 145879 106000 145888
rect 120752 145928 121120 145937
rect 120792 145888 120834 145928
rect 120874 145888 120916 145928
rect 120956 145888 120998 145928
rect 121038 145888 121080 145928
rect 120752 145879 121120 145888
rect 135872 145928 136240 145937
rect 135912 145888 135954 145928
rect 135994 145888 136036 145928
rect 136076 145888 136118 145928
rect 136158 145888 136200 145928
rect 135872 145879 136240 145888
rect 150992 145928 151360 145937
rect 151032 145888 151074 145928
rect 151114 145888 151156 145928
rect 151196 145888 151238 145928
rect 151278 145888 151320 145928
rect 150992 145879 151360 145888
rect 104392 145172 104760 145181
rect 104432 145132 104474 145172
rect 104514 145132 104556 145172
rect 104596 145132 104638 145172
rect 104678 145132 104720 145172
rect 104392 145123 104760 145132
rect 119512 145172 119880 145181
rect 119552 145132 119594 145172
rect 119634 145132 119676 145172
rect 119716 145132 119758 145172
rect 119798 145132 119840 145172
rect 119512 145123 119880 145132
rect 134632 145172 135000 145181
rect 134672 145132 134714 145172
rect 134754 145132 134796 145172
rect 134836 145132 134878 145172
rect 134918 145132 134960 145172
rect 134632 145123 135000 145132
rect 149752 145172 150120 145181
rect 149792 145132 149834 145172
rect 149874 145132 149916 145172
rect 149956 145132 149998 145172
rect 150038 145132 150080 145172
rect 149752 145123 150120 145132
rect 105632 144416 106000 144425
rect 105672 144376 105714 144416
rect 105754 144376 105796 144416
rect 105836 144376 105878 144416
rect 105918 144376 105960 144416
rect 105632 144367 106000 144376
rect 120752 144416 121120 144425
rect 120792 144376 120834 144416
rect 120874 144376 120916 144416
rect 120956 144376 120998 144416
rect 121038 144376 121080 144416
rect 120752 144367 121120 144376
rect 135872 144416 136240 144425
rect 135912 144376 135954 144416
rect 135994 144376 136036 144416
rect 136076 144376 136118 144416
rect 136158 144376 136200 144416
rect 135872 144367 136240 144376
rect 150992 144416 151360 144425
rect 151032 144376 151074 144416
rect 151114 144376 151156 144416
rect 151196 144376 151238 144416
rect 151278 144376 151320 144416
rect 150992 144367 151360 144376
rect 104392 143660 104760 143669
rect 104432 143620 104474 143660
rect 104514 143620 104556 143660
rect 104596 143620 104638 143660
rect 104678 143620 104720 143660
rect 104392 143611 104760 143620
rect 119512 143660 119880 143669
rect 119552 143620 119594 143660
rect 119634 143620 119676 143660
rect 119716 143620 119758 143660
rect 119798 143620 119840 143660
rect 119512 143611 119880 143620
rect 134632 143660 135000 143669
rect 134672 143620 134714 143660
rect 134754 143620 134796 143660
rect 134836 143620 134878 143660
rect 134918 143620 134960 143660
rect 134632 143611 135000 143620
rect 149752 143660 150120 143669
rect 149792 143620 149834 143660
rect 149874 143620 149916 143660
rect 149956 143620 149998 143660
rect 150038 143620 150080 143660
rect 149752 143611 150120 143620
rect 105632 142904 106000 142913
rect 105672 142864 105714 142904
rect 105754 142864 105796 142904
rect 105836 142864 105878 142904
rect 105918 142864 105960 142904
rect 105632 142855 106000 142864
rect 120752 142904 121120 142913
rect 120792 142864 120834 142904
rect 120874 142864 120916 142904
rect 120956 142864 120998 142904
rect 121038 142864 121080 142904
rect 120752 142855 121120 142864
rect 135872 142904 136240 142913
rect 135912 142864 135954 142904
rect 135994 142864 136036 142904
rect 136076 142864 136118 142904
rect 136158 142864 136200 142904
rect 135872 142855 136240 142864
rect 150992 142904 151360 142913
rect 151032 142864 151074 142904
rect 151114 142864 151156 142904
rect 151196 142864 151238 142904
rect 151278 142864 151320 142904
rect 150992 142855 151360 142864
rect 104392 142148 104760 142157
rect 104432 142108 104474 142148
rect 104514 142108 104556 142148
rect 104596 142108 104638 142148
rect 104678 142108 104720 142148
rect 104392 142099 104760 142108
rect 119512 142148 119880 142157
rect 119552 142108 119594 142148
rect 119634 142108 119676 142148
rect 119716 142108 119758 142148
rect 119798 142108 119840 142148
rect 119512 142099 119880 142108
rect 134632 142148 135000 142157
rect 134672 142108 134714 142148
rect 134754 142108 134796 142148
rect 134836 142108 134878 142148
rect 134918 142108 134960 142148
rect 134632 142099 135000 142108
rect 149752 142148 150120 142157
rect 149792 142108 149834 142148
rect 149874 142108 149916 142148
rect 149956 142108 149998 142148
rect 150038 142108 150080 142148
rect 149752 142099 150120 142108
rect 105632 141392 106000 141401
rect 105672 141352 105714 141392
rect 105754 141352 105796 141392
rect 105836 141352 105878 141392
rect 105918 141352 105960 141392
rect 105632 141343 106000 141352
rect 120752 141392 121120 141401
rect 120792 141352 120834 141392
rect 120874 141352 120916 141392
rect 120956 141352 120998 141392
rect 121038 141352 121080 141392
rect 120752 141343 121120 141352
rect 135872 141392 136240 141401
rect 135912 141352 135954 141392
rect 135994 141352 136036 141392
rect 136076 141352 136118 141392
rect 136158 141352 136200 141392
rect 135872 141343 136240 141352
rect 150992 141392 151360 141401
rect 151032 141352 151074 141392
rect 151114 141352 151156 141392
rect 151196 141352 151238 141392
rect 151278 141352 151320 141392
rect 150992 141343 151360 141352
rect 104392 140636 104760 140645
rect 104432 140596 104474 140636
rect 104514 140596 104556 140636
rect 104596 140596 104638 140636
rect 104678 140596 104720 140636
rect 104392 140587 104760 140596
rect 119512 140636 119880 140645
rect 119552 140596 119594 140636
rect 119634 140596 119676 140636
rect 119716 140596 119758 140636
rect 119798 140596 119840 140636
rect 119512 140587 119880 140596
rect 134632 140636 135000 140645
rect 134672 140596 134714 140636
rect 134754 140596 134796 140636
rect 134836 140596 134878 140636
rect 134918 140596 134960 140636
rect 134632 140587 135000 140596
rect 149752 140636 150120 140645
rect 149792 140596 149834 140636
rect 149874 140596 149916 140636
rect 149956 140596 149998 140636
rect 150038 140596 150080 140636
rect 149752 140587 150120 140596
rect 105632 139880 106000 139889
rect 105672 139840 105714 139880
rect 105754 139840 105796 139880
rect 105836 139840 105878 139880
rect 105918 139840 105960 139880
rect 105632 139831 106000 139840
rect 120752 139880 121120 139889
rect 120792 139840 120834 139880
rect 120874 139840 120916 139880
rect 120956 139840 120998 139880
rect 121038 139840 121080 139880
rect 120752 139831 121120 139840
rect 135872 139880 136240 139889
rect 135912 139840 135954 139880
rect 135994 139840 136036 139880
rect 136076 139840 136118 139880
rect 136158 139840 136200 139880
rect 135872 139831 136240 139840
rect 150992 139880 151360 139889
rect 151032 139840 151074 139880
rect 151114 139840 151156 139880
rect 151196 139840 151238 139880
rect 151278 139840 151320 139880
rect 150992 139831 151360 139840
rect 104392 139124 104760 139133
rect 104432 139084 104474 139124
rect 104514 139084 104556 139124
rect 104596 139084 104638 139124
rect 104678 139084 104720 139124
rect 104392 139075 104760 139084
rect 119512 139124 119880 139133
rect 119552 139084 119594 139124
rect 119634 139084 119676 139124
rect 119716 139084 119758 139124
rect 119798 139084 119840 139124
rect 119512 139075 119880 139084
rect 134632 139124 135000 139133
rect 134672 139084 134714 139124
rect 134754 139084 134796 139124
rect 134836 139084 134878 139124
rect 134918 139084 134960 139124
rect 134632 139075 135000 139084
rect 149752 139124 150120 139133
rect 149792 139084 149834 139124
rect 149874 139084 149916 139124
rect 149956 139084 149998 139124
rect 150038 139084 150080 139124
rect 149752 139075 150120 139084
rect 105632 138368 106000 138377
rect 105672 138328 105714 138368
rect 105754 138328 105796 138368
rect 105836 138328 105878 138368
rect 105918 138328 105960 138368
rect 105632 138319 106000 138328
rect 120752 138368 121120 138377
rect 120792 138328 120834 138368
rect 120874 138328 120916 138368
rect 120956 138328 120998 138368
rect 121038 138328 121080 138368
rect 120752 138319 121120 138328
rect 135872 138368 136240 138377
rect 135912 138328 135954 138368
rect 135994 138328 136036 138368
rect 136076 138328 136118 138368
rect 136158 138328 136200 138368
rect 135872 138319 136240 138328
rect 150992 138368 151360 138377
rect 151032 138328 151074 138368
rect 151114 138328 151156 138368
rect 151196 138328 151238 138368
rect 151278 138328 151320 138368
rect 150992 138319 151360 138328
rect 104392 137612 104760 137621
rect 104432 137572 104474 137612
rect 104514 137572 104556 137612
rect 104596 137572 104638 137612
rect 104678 137572 104720 137612
rect 104392 137563 104760 137572
rect 119512 137612 119880 137621
rect 119552 137572 119594 137612
rect 119634 137572 119676 137612
rect 119716 137572 119758 137612
rect 119798 137572 119840 137612
rect 119512 137563 119880 137572
rect 134632 137612 135000 137621
rect 134672 137572 134714 137612
rect 134754 137572 134796 137612
rect 134836 137572 134878 137612
rect 134918 137572 134960 137612
rect 134632 137563 135000 137572
rect 149752 137612 150120 137621
rect 149792 137572 149834 137612
rect 149874 137572 149916 137612
rect 149956 137572 149998 137612
rect 150038 137572 150080 137612
rect 149752 137563 150120 137572
rect 105632 136856 106000 136865
rect 105672 136816 105714 136856
rect 105754 136816 105796 136856
rect 105836 136816 105878 136856
rect 105918 136816 105960 136856
rect 105632 136807 106000 136816
rect 120752 136856 121120 136865
rect 120792 136816 120834 136856
rect 120874 136816 120916 136856
rect 120956 136816 120998 136856
rect 121038 136816 121080 136856
rect 120752 136807 121120 136816
rect 135872 136856 136240 136865
rect 135912 136816 135954 136856
rect 135994 136816 136036 136856
rect 136076 136816 136118 136856
rect 136158 136816 136200 136856
rect 135872 136807 136240 136816
rect 150992 136856 151360 136865
rect 151032 136816 151074 136856
rect 151114 136816 151156 136856
rect 151196 136816 151238 136856
rect 151278 136816 151320 136856
rect 150992 136807 151360 136816
rect 104392 136100 104760 136109
rect 104432 136060 104474 136100
rect 104514 136060 104556 136100
rect 104596 136060 104638 136100
rect 104678 136060 104720 136100
rect 104392 136051 104760 136060
rect 119512 136100 119880 136109
rect 119552 136060 119594 136100
rect 119634 136060 119676 136100
rect 119716 136060 119758 136100
rect 119798 136060 119840 136100
rect 119512 136051 119880 136060
rect 134632 136100 135000 136109
rect 134672 136060 134714 136100
rect 134754 136060 134796 136100
rect 134836 136060 134878 136100
rect 134918 136060 134960 136100
rect 134632 136051 135000 136060
rect 149752 136100 150120 136109
rect 149792 136060 149834 136100
rect 149874 136060 149916 136100
rect 149956 136060 149998 136100
rect 150038 136060 150080 136100
rect 149752 136051 150120 136060
rect 105632 135344 106000 135353
rect 105672 135304 105714 135344
rect 105754 135304 105796 135344
rect 105836 135304 105878 135344
rect 105918 135304 105960 135344
rect 105632 135295 106000 135304
rect 120752 135344 121120 135353
rect 120792 135304 120834 135344
rect 120874 135304 120916 135344
rect 120956 135304 120998 135344
rect 121038 135304 121080 135344
rect 120752 135295 121120 135304
rect 135872 135344 136240 135353
rect 135912 135304 135954 135344
rect 135994 135304 136036 135344
rect 136076 135304 136118 135344
rect 136158 135304 136200 135344
rect 135872 135295 136240 135304
rect 150992 135344 151360 135353
rect 151032 135304 151074 135344
rect 151114 135304 151156 135344
rect 151196 135304 151238 135344
rect 151278 135304 151320 135344
rect 150992 135295 151360 135304
rect 104392 134588 104760 134597
rect 104432 134548 104474 134588
rect 104514 134548 104556 134588
rect 104596 134548 104638 134588
rect 104678 134548 104720 134588
rect 104392 134539 104760 134548
rect 119512 134588 119880 134597
rect 119552 134548 119594 134588
rect 119634 134548 119676 134588
rect 119716 134548 119758 134588
rect 119798 134548 119840 134588
rect 119512 134539 119880 134548
rect 134632 134588 135000 134597
rect 134672 134548 134714 134588
rect 134754 134548 134796 134588
rect 134836 134548 134878 134588
rect 134918 134548 134960 134588
rect 134632 134539 135000 134548
rect 149752 134588 150120 134597
rect 149792 134548 149834 134588
rect 149874 134548 149916 134588
rect 149956 134548 149998 134588
rect 150038 134548 150080 134588
rect 149752 134539 150120 134548
rect 105632 133832 106000 133841
rect 105672 133792 105714 133832
rect 105754 133792 105796 133832
rect 105836 133792 105878 133832
rect 105918 133792 105960 133832
rect 105632 133783 106000 133792
rect 120752 133832 121120 133841
rect 120792 133792 120834 133832
rect 120874 133792 120916 133832
rect 120956 133792 120998 133832
rect 121038 133792 121080 133832
rect 120752 133783 121120 133792
rect 135872 133832 136240 133841
rect 135912 133792 135954 133832
rect 135994 133792 136036 133832
rect 136076 133792 136118 133832
rect 136158 133792 136200 133832
rect 135872 133783 136240 133792
rect 150992 133832 151360 133841
rect 151032 133792 151074 133832
rect 151114 133792 151156 133832
rect 151196 133792 151238 133832
rect 151278 133792 151320 133832
rect 150992 133783 151360 133792
rect 104392 133076 104760 133085
rect 104432 133036 104474 133076
rect 104514 133036 104556 133076
rect 104596 133036 104638 133076
rect 104678 133036 104720 133076
rect 104392 133027 104760 133036
rect 119512 133076 119880 133085
rect 119552 133036 119594 133076
rect 119634 133036 119676 133076
rect 119716 133036 119758 133076
rect 119798 133036 119840 133076
rect 119512 133027 119880 133036
rect 134632 133076 135000 133085
rect 134672 133036 134714 133076
rect 134754 133036 134796 133076
rect 134836 133036 134878 133076
rect 134918 133036 134960 133076
rect 134632 133027 135000 133036
rect 149752 133076 150120 133085
rect 149792 133036 149834 133076
rect 149874 133036 149916 133076
rect 149956 133036 149998 133076
rect 150038 133036 150080 133076
rect 149752 133027 150120 133036
rect 105632 132320 106000 132329
rect 105672 132280 105714 132320
rect 105754 132280 105796 132320
rect 105836 132280 105878 132320
rect 105918 132280 105960 132320
rect 105632 132271 106000 132280
rect 120752 132320 121120 132329
rect 120792 132280 120834 132320
rect 120874 132280 120916 132320
rect 120956 132280 120998 132320
rect 121038 132280 121080 132320
rect 120752 132271 121120 132280
rect 135872 132320 136240 132329
rect 135912 132280 135954 132320
rect 135994 132280 136036 132320
rect 136076 132280 136118 132320
rect 136158 132280 136200 132320
rect 135872 132271 136240 132280
rect 150992 132320 151360 132329
rect 151032 132280 151074 132320
rect 151114 132280 151156 132320
rect 151196 132280 151238 132320
rect 151278 132280 151320 132320
rect 150992 132271 151360 132280
rect 104392 131564 104760 131573
rect 104432 131524 104474 131564
rect 104514 131524 104556 131564
rect 104596 131524 104638 131564
rect 104678 131524 104720 131564
rect 104392 131515 104760 131524
rect 119512 131564 119880 131573
rect 119552 131524 119594 131564
rect 119634 131524 119676 131564
rect 119716 131524 119758 131564
rect 119798 131524 119840 131564
rect 119512 131515 119880 131524
rect 134632 131564 135000 131573
rect 134672 131524 134714 131564
rect 134754 131524 134796 131564
rect 134836 131524 134878 131564
rect 134918 131524 134960 131564
rect 134632 131515 135000 131524
rect 149752 131564 150120 131573
rect 149792 131524 149834 131564
rect 149874 131524 149916 131564
rect 149956 131524 149998 131564
rect 150038 131524 150080 131564
rect 149752 131515 150120 131524
rect 105632 130808 106000 130817
rect 105672 130768 105714 130808
rect 105754 130768 105796 130808
rect 105836 130768 105878 130808
rect 105918 130768 105960 130808
rect 105632 130759 106000 130768
rect 120752 130808 121120 130817
rect 120792 130768 120834 130808
rect 120874 130768 120916 130808
rect 120956 130768 120998 130808
rect 121038 130768 121080 130808
rect 120752 130759 121120 130768
rect 135872 130808 136240 130817
rect 135912 130768 135954 130808
rect 135994 130768 136036 130808
rect 136076 130768 136118 130808
rect 136158 130768 136200 130808
rect 135872 130759 136240 130768
rect 150992 130808 151360 130817
rect 151032 130768 151074 130808
rect 151114 130768 151156 130808
rect 151196 130768 151238 130808
rect 151278 130768 151320 130808
rect 150992 130759 151360 130768
rect 104392 130052 104760 130061
rect 104432 130012 104474 130052
rect 104514 130012 104556 130052
rect 104596 130012 104638 130052
rect 104678 130012 104720 130052
rect 104392 130003 104760 130012
rect 119512 130052 119880 130061
rect 119552 130012 119594 130052
rect 119634 130012 119676 130052
rect 119716 130012 119758 130052
rect 119798 130012 119840 130052
rect 119512 130003 119880 130012
rect 134632 130052 135000 130061
rect 134672 130012 134714 130052
rect 134754 130012 134796 130052
rect 134836 130012 134878 130052
rect 134918 130012 134960 130052
rect 134632 130003 135000 130012
rect 149752 130052 150120 130061
rect 149792 130012 149834 130052
rect 149874 130012 149916 130052
rect 149956 130012 149998 130052
rect 150038 130012 150080 130052
rect 149752 130003 150120 130012
rect 105632 129296 106000 129305
rect 105672 129256 105714 129296
rect 105754 129256 105796 129296
rect 105836 129256 105878 129296
rect 105918 129256 105960 129296
rect 105632 129247 106000 129256
rect 120752 129296 121120 129305
rect 120792 129256 120834 129296
rect 120874 129256 120916 129296
rect 120956 129256 120998 129296
rect 121038 129256 121080 129296
rect 120752 129247 121120 129256
rect 135872 129296 136240 129305
rect 135912 129256 135954 129296
rect 135994 129256 136036 129296
rect 136076 129256 136118 129296
rect 136158 129256 136200 129296
rect 135872 129247 136240 129256
rect 150992 129296 151360 129305
rect 151032 129256 151074 129296
rect 151114 129256 151156 129296
rect 151196 129256 151238 129296
rect 151278 129256 151320 129296
rect 150992 129247 151360 129256
rect 104392 128540 104760 128549
rect 104432 128500 104474 128540
rect 104514 128500 104556 128540
rect 104596 128500 104638 128540
rect 104678 128500 104720 128540
rect 104392 128491 104760 128500
rect 119512 128540 119880 128549
rect 119552 128500 119594 128540
rect 119634 128500 119676 128540
rect 119716 128500 119758 128540
rect 119798 128500 119840 128540
rect 119512 128491 119880 128500
rect 134632 128540 135000 128549
rect 134672 128500 134714 128540
rect 134754 128500 134796 128540
rect 134836 128500 134878 128540
rect 134918 128500 134960 128540
rect 134632 128491 135000 128500
rect 149752 128540 150120 128549
rect 149792 128500 149834 128540
rect 149874 128500 149916 128540
rect 149956 128500 149998 128540
rect 150038 128500 150080 128540
rect 149752 128491 150120 128500
rect 105632 127784 106000 127793
rect 105672 127744 105714 127784
rect 105754 127744 105796 127784
rect 105836 127744 105878 127784
rect 105918 127744 105960 127784
rect 105632 127735 106000 127744
rect 120752 127784 121120 127793
rect 120792 127744 120834 127784
rect 120874 127744 120916 127784
rect 120956 127744 120998 127784
rect 121038 127744 121080 127784
rect 120752 127735 121120 127744
rect 135872 127784 136240 127793
rect 135912 127744 135954 127784
rect 135994 127744 136036 127784
rect 136076 127744 136118 127784
rect 136158 127744 136200 127784
rect 135872 127735 136240 127744
rect 150992 127784 151360 127793
rect 151032 127744 151074 127784
rect 151114 127744 151156 127784
rect 151196 127744 151238 127784
rect 151278 127744 151320 127784
rect 150992 127735 151360 127744
rect 104392 127028 104760 127037
rect 104432 126988 104474 127028
rect 104514 126988 104556 127028
rect 104596 126988 104638 127028
rect 104678 126988 104720 127028
rect 104392 126979 104760 126988
rect 119512 127028 119880 127037
rect 119552 126988 119594 127028
rect 119634 126988 119676 127028
rect 119716 126988 119758 127028
rect 119798 126988 119840 127028
rect 119512 126979 119880 126988
rect 134632 127028 135000 127037
rect 134672 126988 134714 127028
rect 134754 126988 134796 127028
rect 134836 126988 134878 127028
rect 134918 126988 134960 127028
rect 134632 126979 135000 126988
rect 149752 127028 150120 127037
rect 149792 126988 149834 127028
rect 149874 126988 149916 127028
rect 149956 126988 149998 127028
rect 150038 126988 150080 127028
rect 149752 126979 150120 126988
rect 105632 126272 106000 126281
rect 105672 126232 105714 126272
rect 105754 126232 105796 126272
rect 105836 126232 105878 126272
rect 105918 126232 105960 126272
rect 105632 126223 106000 126232
rect 120752 126272 121120 126281
rect 120792 126232 120834 126272
rect 120874 126232 120916 126272
rect 120956 126232 120998 126272
rect 121038 126232 121080 126272
rect 120752 126223 121120 126232
rect 135872 126272 136240 126281
rect 135912 126232 135954 126272
rect 135994 126232 136036 126272
rect 136076 126232 136118 126272
rect 136158 126232 136200 126272
rect 135872 126223 136240 126232
rect 150992 126272 151360 126281
rect 151032 126232 151074 126272
rect 151114 126232 151156 126272
rect 151196 126232 151238 126272
rect 151278 126232 151320 126272
rect 150992 126223 151360 126232
rect 104392 125516 104760 125525
rect 104432 125476 104474 125516
rect 104514 125476 104556 125516
rect 104596 125476 104638 125516
rect 104678 125476 104720 125516
rect 104392 125467 104760 125476
rect 119512 125516 119880 125525
rect 119552 125476 119594 125516
rect 119634 125476 119676 125516
rect 119716 125476 119758 125516
rect 119798 125476 119840 125516
rect 119512 125467 119880 125476
rect 134632 125516 135000 125525
rect 134672 125476 134714 125516
rect 134754 125476 134796 125516
rect 134836 125476 134878 125516
rect 134918 125476 134960 125516
rect 134632 125467 135000 125476
rect 149752 125516 150120 125525
rect 149792 125476 149834 125516
rect 149874 125476 149916 125516
rect 149956 125476 149998 125516
rect 150038 125476 150080 125516
rect 149752 125467 150120 125476
rect 105632 124760 106000 124769
rect 105672 124720 105714 124760
rect 105754 124720 105796 124760
rect 105836 124720 105878 124760
rect 105918 124720 105960 124760
rect 105632 124711 106000 124720
rect 120752 124760 121120 124769
rect 120792 124720 120834 124760
rect 120874 124720 120916 124760
rect 120956 124720 120998 124760
rect 121038 124720 121080 124760
rect 120752 124711 121120 124720
rect 135872 124760 136240 124769
rect 135912 124720 135954 124760
rect 135994 124720 136036 124760
rect 136076 124720 136118 124760
rect 136158 124720 136200 124760
rect 135872 124711 136240 124720
rect 150992 124760 151360 124769
rect 151032 124720 151074 124760
rect 151114 124720 151156 124760
rect 151196 124720 151238 124760
rect 151278 124720 151320 124760
rect 150992 124711 151360 124720
rect 104392 124004 104760 124013
rect 104432 123964 104474 124004
rect 104514 123964 104556 124004
rect 104596 123964 104638 124004
rect 104678 123964 104720 124004
rect 104392 123955 104760 123964
rect 119512 124004 119880 124013
rect 119552 123964 119594 124004
rect 119634 123964 119676 124004
rect 119716 123964 119758 124004
rect 119798 123964 119840 124004
rect 119512 123955 119880 123964
rect 134632 124004 135000 124013
rect 134672 123964 134714 124004
rect 134754 123964 134796 124004
rect 134836 123964 134878 124004
rect 134918 123964 134960 124004
rect 134632 123955 135000 123964
rect 149752 124004 150120 124013
rect 149792 123964 149834 124004
rect 149874 123964 149916 124004
rect 149956 123964 149998 124004
rect 150038 123964 150080 124004
rect 149752 123955 150120 123964
rect 105632 123248 106000 123257
rect 105672 123208 105714 123248
rect 105754 123208 105796 123248
rect 105836 123208 105878 123248
rect 105918 123208 105960 123248
rect 105632 123199 106000 123208
rect 120752 123248 121120 123257
rect 120792 123208 120834 123248
rect 120874 123208 120916 123248
rect 120956 123208 120998 123248
rect 121038 123208 121080 123248
rect 120752 123199 121120 123208
rect 135872 123248 136240 123257
rect 135912 123208 135954 123248
rect 135994 123208 136036 123248
rect 136076 123208 136118 123248
rect 136158 123208 136200 123248
rect 135872 123199 136240 123208
rect 150992 123248 151360 123257
rect 151032 123208 151074 123248
rect 151114 123208 151156 123248
rect 151196 123208 151238 123248
rect 151278 123208 151320 123248
rect 150992 123199 151360 123208
rect 104392 122492 104760 122501
rect 104432 122452 104474 122492
rect 104514 122452 104556 122492
rect 104596 122452 104638 122492
rect 104678 122452 104720 122492
rect 104392 122443 104760 122452
rect 119512 122492 119880 122501
rect 119552 122452 119594 122492
rect 119634 122452 119676 122492
rect 119716 122452 119758 122492
rect 119798 122452 119840 122492
rect 119512 122443 119880 122452
rect 134632 122492 135000 122501
rect 134672 122452 134714 122492
rect 134754 122452 134796 122492
rect 134836 122452 134878 122492
rect 134918 122452 134960 122492
rect 134632 122443 135000 122452
rect 149752 122492 150120 122501
rect 149792 122452 149834 122492
rect 149874 122452 149916 122492
rect 149956 122452 149998 122492
rect 150038 122452 150080 122492
rect 149752 122443 150120 122452
rect 105632 121736 106000 121745
rect 105672 121696 105714 121736
rect 105754 121696 105796 121736
rect 105836 121696 105878 121736
rect 105918 121696 105960 121736
rect 105632 121687 106000 121696
rect 120752 121736 121120 121745
rect 120792 121696 120834 121736
rect 120874 121696 120916 121736
rect 120956 121696 120998 121736
rect 121038 121696 121080 121736
rect 120752 121687 121120 121696
rect 135872 121736 136240 121745
rect 135912 121696 135954 121736
rect 135994 121696 136036 121736
rect 136076 121696 136118 121736
rect 136158 121696 136200 121736
rect 135872 121687 136240 121696
rect 150992 121736 151360 121745
rect 151032 121696 151074 121736
rect 151114 121696 151156 121736
rect 151196 121696 151238 121736
rect 151278 121696 151320 121736
rect 150992 121687 151360 121696
rect 104392 120980 104760 120989
rect 104432 120940 104474 120980
rect 104514 120940 104556 120980
rect 104596 120940 104638 120980
rect 104678 120940 104720 120980
rect 104392 120931 104760 120940
rect 119512 120980 119880 120989
rect 119552 120940 119594 120980
rect 119634 120940 119676 120980
rect 119716 120940 119758 120980
rect 119798 120940 119840 120980
rect 119512 120931 119880 120940
rect 134632 120980 135000 120989
rect 134672 120940 134714 120980
rect 134754 120940 134796 120980
rect 134836 120940 134878 120980
rect 134918 120940 134960 120980
rect 134632 120931 135000 120940
rect 149752 120980 150120 120989
rect 149792 120940 149834 120980
rect 149874 120940 149916 120980
rect 149956 120940 149998 120980
rect 150038 120940 150080 120980
rect 149752 120931 150120 120940
rect 105632 120224 106000 120233
rect 105672 120184 105714 120224
rect 105754 120184 105796 120224
rect 105836 120184 105878 120224
rect 105918 120184 105960 120224
rect 105632 120175 106000 120184
rect 120752 120224 121120 120233
rect 120792 120184 120834 120224
rect 120874 120184 120916 120224
rect 120956 120184 120998 120224
rect 121038 120184 121080 120224
rect 120752 120175 121120 120184
rect 135872 120224 136240 120233
rect 135912 120184 135954 120224
rect 135994 120184 136036 120224
rect 136076 120184 136118 120224
rect 136158 120184 136200 120224
rect 135872 120175 136240 120184
rect 150992 120224 151360 120233
rect 151032 120184 151074 120224
rect 151114 120184 151156 120224
rect 151196 120184 151238 120224
rect 151278 120184 151320 120224
rect 150992 120175 151360 120184
rect 104392 119468 104760 119477
rect 104432 119428 104474 119468
rect 104514 119428 104556 119468
rect 104596 119428 104638 119468
rect 104678 119428 104720 119468
rect 104392 119419 104760 119428
rect 119512 119468 119880 119477
rect 119552 119428 119594 119468
rect 119634 119428 119676 119468
rect 119716 119428 119758 119468
rect 119798 119428 119840 119468
rect 119512 119419 119880 119428
rect 134632 119468 135000 119477
rect 134672 119428 134714 119468
rect 134754 119428 134796 119468
rect 134836 119428 134878 119468
rect 134918 119428 134960 119468
rect 134632 119419 135000 119428
rect 149752 119468 150120 119477
rect 149792 119428 149834 119468
rect 149874 119428 149916 119468
rect 149956 119428 149998 119468
rect 150038 119428 150080 119468
rect 149752 119419 150120 119428
rect 105632 118712 106000 118721
rect 105672 118672 105714 118712
rect 105754 118672 105796 118712
rect 105836 118672 105878 118712
rect 105918 118672 105960 118712
rect 105632 118663 106000 118672
rect 120752 118712 121120 118721
rect 120792 118672 120834 118712
rect 120874 118672 120916 118712
rect 120956 118672 120998 118712
rect 121038 118672 121080 118712
rect 120752 118663 121120 118672
rect 135872 118712 136240 118721
rect 135912 118672 135954 118712
rect 135994 118672 136036 118712
rect 136076 118672 136118 118712
rect 136158 118672 136200 118712
rect 135872 118663 136240 118672
rect 150992 118712 151360 118721
rect 151032 118672 151074 118712
rect 151114 118672 151156 118712
rect 151196 118672 151238 118712
rect 151278 118672 151320 118712
rect 150992 118663 151360 118672
rect 104392 117956 104760 117965
rect 104432 117916 104474 117956
rect 104514 117916 104556 117956
rect 104596 117916 104638 117956
rect 104678 117916 104720 117956
rect 104392 117907 104760 117916
rect 119512 117956 119880 117965
rect 119552 117916 119594 117956
rect 119634 117916 119676 117956
rect 119716 117916 119758 117956
rect 119798 117916 119840 117956
rect 119512 117907 119880 117916
rect 134632 117956 135000 117965
rect 134672 117916 134714 117956
rect 134754 117916 134796 117956
rect 134836 117916 134878 117956
rect 134918 117916 134960 117956
rect 134632 117907 135000 117916
rect 149752 117956 150120 117965
rect 149792 117916 149834 117956
rect 149874 117916 149916 117956
rect 149956 117916 149998 117956
rect 150038 117916 150080 117956
rect 149752 117907 150120 117916
rect 105632 117200 106000 117209
rect 105672 117160 105714 117200
rect 105754 117160 105796 117200
rect 105836 117160 105878 117200
rect 105918 117160 105960 117200
rect 105632 117151 106000 117160
rect 120752 117200 121120 117209
rect 120792 117160 120834 117200
rect 120874 117160 120916 117200
rect 120956 117160 120998 117200
rect 121038 117160 121080 117200
rect 120752 117151 121120 117160
rect 135872 117200 136240 117209
rect 135912 117160 135954 117200
rect 135994 117160 136036 117200
rect 136076 117160 136118 117200
rect 136158 117160 136200 117200
rect 135872 117151 136240 117160
rect 150992 117200 151360 117209
rect 151032 117160 151074 117200
rect 151114 117160 151156 117200
rect 151196 117160 151238 117200
rect 151278 117160 151320 117200
rect 150992 117151 151360 117160
rect 104392 116444 104760 116453
rect 104432 116404 104474 116444
rect 104514 116404 104556 116444
rect 104596 116404 104638 116444
rect 104678 116404 104720 116444
rect 104392 116395 104760 116404
rect 119512 116444 119880 116453
rect 119552 116404 119594 116444
rect 119634 116404 119676 116444
rect 119716 116404 119758 116444
rect 119798 116404 119840 116444
rect 119512 116395 119880 116404
rect 134632 116444 135000 116453
rect 134672 116404 134714 116444
rect 134754 116404 134796 116444
rect 134836 116404 134878 116444
rect 134918 116404 134960 116444
rect 134632 116395 135000 116404
rect 149752 116444 150120 116453
rect 149792 116404 149834 116444
rect 149874 116404 149916 116444
rect 149956 116404 149998 116444
rect 150038 116404 150080 116444
rect 149752 116395 150120 116404
rect 105632 115688 106000 115697
rect 105672 115648 105714 115688
rect 105754 115648 105796 115688
rect 105836 115648 105878 115688
rect 105918 115648 105960 115688
rect 105632 115639 106000 115648
rect 120752 115688 121120 115697
rect 120792 115648 120834 115688
rect 120874 115648 120916 115688
rect 120956 115648 120998 115688
rect 121038 115648 121080 115688
rect 120752 115639 121120 115648
rect 135872 115688 136240 115697
rect 135912 115648 135954 115688
rect 135994 115648 136036 115688
rect 136076 115648 136118 115688
rect 136158 115648 136200 115688
rect 135872 115639 136240 115648
rect 150992 115688 151360 115697
rect 151032 115648 151074 115688
rect 151114 115648 151156 115688
rect 151196 115648 151238 115688
rect 151278 115648 151320 115688
rect 150992 115639 151360 115648
rect 104392 114932 104760 114941
rect 104432 114892 104474 114932
rect 104514 114892 104556 114932
rect 104596 114892 104638 114932
rect 104678 114892 104720 114932
rect 104392 114883 104760 114892
rect 119512 114932 119880 114941
rect 119552 114892 119594 114932
rect 119634 114892 119676 114932
rect 119716 114892 119758 114932
rect 119798 114892 119840 114932
rect 119512 114883 119880 114892
rect 134632 114932 135000 114941
rect 134672 114892 134714 114932
rect 134754 114892 134796 114932
rect 134836 114892 134878 114932
rect 134918 114892 134960 114932
rect 134632 114883 135000 114892
rect 149752 114932 150120 114941
rect 149792 114892 149834 114932
rect 149874 114892 149916 114932
rect 149956 114892 149998 114932
rect 150038 114892 150080 114932
rect 149752 114883 150120 114892
rect 105632 114176 106000 114185
rect 105672 114136 105714 114176
rect 105754 114136 105796 114176
rect 105836 114136 105878 114176
rect 105918 114136 105960 114176
rect 105632 114127 106000 114136
rect 120752 114176 121120 114185
rect 120792 114136 120834 114176
rect 120874 114136 120916 114176
rect 120956 114136 120998 114176
rect 121038 114136 121080 114176
rect 120752 114127 121120 114136
rect 135872 114176 136240 114185
rect 135912 114136 135954 114176
rect 135994 114136 136036 114176
rect 136076 114136 136118 114176
rect 136158 114136 136200 114176
rect 135872 114127 136240 114136
rect 150992 114176 151360 114185
rect 151032 114136 151074 114176
rect 151114 114136 151156 114176
rect 151196 114136 151238 114176
rect 151278 114136 151320 114176
rect 150992 114127 151360 114136
rect 104392 113420 104760 113429
rect 104432 113380 104474 113420
rect 104514 113380 104556 113420
rect 104596 113380 104638 113420
rect 104678 113380 104720 113420
rect 104392 113371 104760 113380
rect 119512 113420 119880 113429
rect 119552 113380 119594 113420
rect 119634 113380 119676 113420
rect 119716 113380 119758 113420
rect 119798 113380 119840 113420
rect 119512 113371 119880 113380
rect 134632 113420 135000 113429
rect 134672 113380 134714 113420
rect 134754 113380 134796 113420
rect 134836 113380 134878 113420
rect 134918 113380 134960 113420
rect 134632 113371 135000 113380
rect 149752 113420 150120 113429
rect 149792 113380 149834 113420
rect 149874 113380 149916 113420
rect 149956 113380 149998 113420
rect 150038 113380 150080 113420
rect 149752 113371 150120 113380
rect 105632 112664 106000 112673
rect 105672 112624 105714 112664
rect 105754 112624 105796 112664
rect 105836 112624 105878 112664
rect 105918 112624 105960 112664
rect 105632 112615 106000 112624
rect 120752 112664 121120 112673
rect 120792 112624 120834 112664
rect 120874 112624 120916 112664
rect 120956 112624 120998 112664
rect 121038 112624 121080 112664
rect 120752 112615 121120 112624
rect 135872 112664 136240 112673
rect 135912 112624 135954 112664
rect 135994 112624 136036 112664
rect 136076 112624 136118 112664
rect 136158 112624 136200 112664
rect 135872 112615 136240 112624
rect 150992 112664 151360 112673
rect 151032 112624 151074 112664
rect 151114 112624 151156 112664
rect 151196 112624 151238 112664
rect 151278 112624 151320 112664
rect 150992 112615 151360 112624
rect 104392 111908 104760 111917
rect 104432 111868 104474 111908
rect 104514 111868 104556 111908
rect 104596 111868 104638 111908
rect 104678 111868 104720 111908
rect 104392 111859 104760 111868
rect 119512 111908 119880 111917
rect 119552 111868 119594 111908
rect 119634 111868 119676 111908
rect 119716 111868 119758 111908
rect 119798 111868 119840 111908
rect 119512 111859 119880 111868
rect 134632 111908 135000 111917
rect 134672 111868 134714 111908
rect 134754 111868 134796 111908
rect 134836 111868 134878 111908
rect 134918 111868 134960 111908
rect 134632 111859 135000 111868
rect 149752 111908 150120 111917
rect 149792 111868 149834 111908
rect 149874 111868 149916 111908
rect 149956 111868 149998 111908
rect 150038 111868 150080 111908
rect 149752 111859 150120 111868
rect 105632 111152 106000 111161
rect 105672 111112 105714 111152
rect 105754 111112 105796 111152
rect 105836 111112 105878 111152
rect 105918 111112 105960 111152
rect 105632 111103 106000 111112
rect 120752 111152 121120 111161
rect 120792 111112 120834 111152
rect 120874 111112 120916 111152
rect 120956 111112 120998 111152
rect 121038 111112 121080 111152
rect 120752 111103 121120 111112
rect 135872 111152 136240 111161
rect 135912 111112 135954 111152
rect 135994 111112 136036 111152
rect 136076 111112 136118 111152
rect 136158 111112 136200 111152
rect 135872 111103 136240 111112
rect 150992 111152 151360 111161
rect 151032 111112 151074 111152
rect 151114 111112 151156 111152
rect 151196 111112 151238 111152
rect 151278 111112 151320 111152
rect 150992 111103 151360 111112
rect 104392 110396 104760 110405
rect 104432 110356 104474 110396
rect 104514 110356 104556 110396
rect 104596 110356 104638 110396
rect 104678 110356 104720 110396
rect 104392 110347 104760 110356
rect 119512 110396 119880 110405
rect 119552 110356 119594 110396
rect 119634 110356 119676 110396
rect 119716 110356 119758 110396
rect 119798 110356 119840 110396
rect 119512 110347 119880 110356
rect 134632 110396 135000 110405
rect 134672 110356 134714 110396
rect 134754 110356 134796 110396
rect 134836 110356 134878 110396
rect 134918 110356 134960 110396
rect 134632 110347 135000 110356
rect 149752 110396 150120 110405
rect 149792 110356 149834 110396
rect 149874 110356 149916 110396
rect 149956 110356 149998 110396
rect 150038 110356 150080 110396
rect 149752 110347 150120 110356
rect 105632 109640 106000 109649
rect 105672 109600 105714 109640
rect 105754 109600 105796 109640
rect 105836 109600 105878 109640
rect 105918 109600 105960 109640
rect 105632 109591 106000 109600
rect 120752 109640 121120 109649
rect 120792 109600 120834 109640
rect 120874 109600 120916 109640
rect 120956 109600 120998 109640
rect 121038 109600 121080 109640
rect 120752 109591 121120 109600
rect 135872 109640 136240 109649
rect 135912 109600 135954 109640
rect 135994 109600 136036 109640
rect 136076 109600 136118 109640
rect 136158 109600 136200 109640
rect 135872 109591 136240 109600
rect 150992 109640 151360 109649
rect 151032 109600 151074 109640
rect 151114 109600 151156 109640
rect 151196 109600 151238 109640
rect 151278 109600 151320 109640
rect 150992 109591 151360 109600
rect 104392 108884 104760 108893
rect 104432 108844 104474 108884
rect 104514 108844 104556 108884
rect 104596 108844 104638 108884
rect 104678 108844 104720 108884
rect 104392 108835 104760 108844
rect 119512 108884 119880 108893
rect 119552 108844 119594 108884
rect 119634 108844 119676 108884
rect 119716 108844 119758 108884
rect 119798 108844 119840 108884
rect 119512 108835 119880 108844
rect 134632 108884 135000 108893
rect 134672 108844 134714 108884
rect 134754 108844 134796 108884
rect 134836 108844 134878 108884
rect 134918 108844 134960 108884
rect 134632 108835 135000 108844
rect 149752 108884 150120 108893
rect 149792 108844 149834 108884
rect 149874 108844 149916 108884
rect 149956 108844 149998 108884
rect 150038 108844 150080 108884
rect 149752 108835 150120 108844
rect 105632 108128 106000 108137
rect 105672 108088 105714 108128
rect 105754 108088 105796 108128
rect 105836 108088 105878 108128
rect 105918 108088 105960 108128
rect 105632 108079 106000 108088
rect 120752 108128 121120 108137
rect 120792 108088 120834 108128
rect 120874 108088 120916 108128
rect 120956 108088 120998 108128
rect 121038 108088 121080 108128
rect 120752 108079 121120 108088
rect 135872 108128 136240 108137
rect 135912 108088 135954 108128
rect 135994 108088 136036 108128
rect 136076 108088 136118 108128
rect 136158 108088 136200 108128
rect 135872 108079 136240 108088
rect 150992 108128 151360 108137
rect 151032 108088 151074 108128
rect 151114 108088 151156 108128
rect 151196 108088 151238 108128
rect 151278 108088 151320 108128
rect 150992 108079 151360 108088
rect 104392 107372 104760 107381
rect 104432 107332 104474 107372
rect 104514 107332 104556 107372
rect 104596 107332 104638 107372
rect 104678 107332 104720 107372
rect 104392 107323 104760 107332
rect 119512 107372 119880 107381
rect 119552 107332 119594 107372
rect 119634 107332 119676 107372
rect 119716 107332 119758 107372
rect 119798 107332 119840 107372
rect 119512 107323 119880 107332
rect 134632 107372 135000 107381
rect 134672 107332 134714 107372
rect 134754 107332 134796 107372
rect 134836 107332 134878 107372
rect 134918 107332 134960 107372
rect 134632 107323 135000 107332
rect 149752 107372 150120 107381
rect 149792 107332 149834 107372
rect 149874 107332 149916 107372
rect 149956 107332 149998 107372
rect 150038 107332 150080 107372
rect 149752 107323 150120 107332
rect 105632 106616 106000 106625
rect 105672 106576 105714 106616
rect 105754 106576 105796 106616
rect 105836 106576 105878 106616
rect 105918 106576 105960 106616
rect 105632 106567 106000 106576
rect 120752 106616 121120 106625
rect 120792 106576 120834 106616
rect 120874 106576 120916 106616
rect 120956 106576 120998 106616
rect 121038 106576 121080 106616
rect 120752 106567 121120 106576
rect 135872 106616 136240 106625
rect 135912 106576 135954 106616
rect 135994 106576 136036 106616
rect 136076 106576 136118 106616
rect 136158 106576 136200 106616
rect 135872 106567 136240 106576
rect 150992 106616 151360 106625
rect 151032 106576 151074 106616
rect 151114 106576 151156 106616
rect 151196 106576 151238 106616
rect 151278 106576 151320 106616
rect 150992 106567 151360 106576
rect 104392 105860 104760 105869
rect 104432 105820 104474 105860
rect 104514 105820 104556 105860
rect 104596 105820 104638 105860
rect 104678 105820 104720 105860
rect 104392 105811 104760 105820
rect 119512 105860 119880 105869
rect 119552 105820 119594 105860
rect 119634 105820 119676 105860
rect 119716 105820 119758 105860
rect 119798 105820 119840 105860
rect 119512 105811 119880 105820
rect 134632 105860 135000 105869
rect 134672 105820 134714 105860
rect 134754 105820 134796 105860
rect 134836 105820 134878 105860
rect 134918 105820 134960 105860
rect 134632 105811 135000 105820
rect 149752 105860 150120 105869
rect 149792 105820 149834 105860
rect 149874 105820 149916 105860
rect 149956 105820 149998 105860
rect 150038 105820 150080 105860
rect 149752 105811 150120 105820
rect 105632 105104 106000 105113
rect 105672 105064 105714 105104
rect 105754 105064 105796 105104
rect 105836 105064 105878 105104
rect 105918 105064 105960 105104
rect 105632 105055 106000 105064
rect 120752 105104 121120 105113
rect 120792 105064 120834 105104
rect 120874 105064 120916 105104
rect 120956 105064 120998 105104
rect 121038 105064 121080 105104
rect 120752 105055 121120 105064
rect 135872 105104 136240 105113
rect 135912 105064 135954 105104
rect 135994 105064 136036 105104
rect 136076 105064 136118 105104
rect 136158 105064 136200 105104
rect 135872 105055 136240 105064
rect 150992 105104 151360 105113
rect 151032 105064 151074 105104
rect 151114 105064 151156 105104
rect 151196 105064 151238 105104
rect 151278 105064 151320 105104
rect 150992 105055 151360 105064
rect 104392 104348 104760 104357
rect 104432 104308 104474 104348
rect 104514 104308 104556 104348
rect 104596 104308 104638 104348
rect 104678 104308 104720 104348
rect 104392 104299 104760 104308
rect 119512 104348 119880 104357
rect 119552 104308 119594 104348
rect 119634 104308 119676 104348
rect 119716 104308 119758 104348
rect 119798 104308 119840 104348
rect 119512 104299 119880 104308
rect 134632 104348 135000 104357
rect 134672 104308 134714 104348
rect 134754 104308 134796 104348
rect 134836 104308 134878 104348
rect 134918 104308 134960 104348
rect 134632 104299 135000 104308
rect 149752 104348 150120 104357
rect 149792 104308 149834 104348
rect 149874 104308 149916 104348
rect 149956 104308 149998 104348
rect 150038 104308 150080 104348
rect 149752 104299 150120 104308
rect 105632 103592 106000 103601
rect 105672 103552 105714 103592
rect 105754 103552 105796 103592
rect 105836 103552 105878 103592
rect 105918 103552 105960 103592
rect 105632 103543 106000 103552
rect 120752 103592 121120 103601
rect 120792 103552 120834 103592
rect 120874 103552 120916 103592
rect 120956 103552 120998 103592
rect 121038 103552 121080 103592
rect 120752 103543 121120 103552
rect 135872 103592 136240 103601
rect 135912 103552 135954 103592
rect 135994 103552 136036 103592
rect 136076 103552 136118 103592
rect 136158 103552 136200 103592
rect 135872 103543 136240 103552
rect 150992 103592 151360 103601
rect 151032 103552 151074 103592
rect 151114 103552 151156 103592
rect 151196 103552 151238 103592
rect 151278 103552 151320 103592
rect 150992 103543 151360 103552
rect 104392 102836 104760 102845
rect 104432 102796 104474 102836
rect 104514 102796 104556 102836
rect 104596 102796 104638 102836
rect 104678 102796 104720 102836
rect 104392 102787 104760 102796
rect 119512 102836 119880 102845
rect 119552 102796 119594 102836
rect 119634 102796 119676 102836
rect 119716 102796 119758 102836
rect 119798 102796 119840 102836
rect 119512 102787 119880 102796
rect 134632 102836 135000 102845
rect 134672 102796 134714 102836
rect 134754 102796 134796 102836
rect 134836 102796 134878 102836
rect 134918 102796 134960 102836
rect 134632 102787 135000 102796
rect 149752 102836 150120 102845
rect 149792 102796 149834 102836
rect 149874 102796 149916 102836
rect 149956 102796 149998 102836
rect 150038 102796 150080 102836
rect 149752 102787 150120 102796
rect 105632 102080 106000 102089
rect 105672 102040 105714 102080
rect 105754 102040 105796 102080
rect 105836 102040 105878 102080
rect 105918 102040 105960 102080
rect 105632 102031 106000 102040
rect 120752 102080 121120 102089
rect 120792 102040 120834 102080
rect 120874 102040 120916 102080
rect 120956 102040 120998 102080
rect 121038 102040 121080 102080
rect 120752 102031 121120 102040
rect 135872 102080 136240 102089
rect 135912 102040 135954 102080
rect 135994 102040 136036 102080
rect 136076 102040 136118 102080
rect 136158 102040 136200 102080
rect 135872 102031 136240 102040
rect 150992 102080 151360 102089
rect 151032 102040 151074 102080
rect 151114 102040 151156 102080
rect 151196 102040 151238 102080
rect 151278 102040 151320 102080
rect 150992 102031 151360 102040
rect 104392 101324 104760 101333
rect 104432 101284 104474 101324
rect 104514 101284 104556 101324
rect 104596 101284 104638 101324
rect 104678 101284 104720 101324
rect 104392 101275 104760 101284
rect 119512 101324 119880 101333
rect 119552 101284 119594 101324
rect 119634 101284 119676 101324
rect 119716 101284 119758 101324
rect 119798 101284 119840 101324
rect 119512 101275 119880 101284
rect 134632 101324 135000 101333
rect 134672 101284 134714 101324
rect 134754 101284 134796 101324
rect 134836 101284 134878 101324
rect 134918 101284 134960 101324
rect 134632 101275 135000 101284
rect 149752 101324 150120 101333
rect 149792 101284 149834 101324
rect 149874 101284 149916 101324
rect 149956 101284 149998 101324
rect 150038 101284 150080 101324
rect 149752 101275 150120 101284
rect 105632 100568 106000 100577
rect 105672 100528 105714 100568
rect 105754 100528 105796 100568
rect 105836 100528 105878 100568
rect 105918 100528 105960 100568
rect 105632 100519 106000 100528
rect 120752 100568 121120 100577
rect 120792 100528 120834 100568
rect 120874 100528 120916 100568
rect 120956 100528 120998 100568
rect 121038 100528 121080 100568
rect 120752 100519 121120 100528
rect 135872 100568 136240 100577
rect 135912 100528 135954 100568
rect 135994 100528 136036 100568
rect 136076 100528 136118 100568
rect 136158 100528 136200 100568
rect 135872 100519 136240 100528
rect 150992 100568 151360 100577
rect 151032 100528 151074 100568
rect 151114 100528 151156 100568
rect 151196 100528 151238 100568
rect 151278 100528 151320 100568
rect 150992 100519 151360 100528
rect 104392 99812 104760 99821
rect 104432 99772 104474 99812
rect 104514 99772 104556 99812
rect 104596 99772 104638 99812
rect 104678 99772 104720 99812
rect 104392 99763 104760 99772
rect 119512 99812 119880 99821
rect 119552 99772 119594 99812
rect 119634 99772 119676 99812
rect 119716 99772 119758 99812
rect 119798 99772 119840 99812
rect 119512 99763 119880 99772
rect 134632 99812 135000 99821
rect 134672 99772 134714 99812
rect 134754 99772 134796 99812
rect 134836 99772 134878 99812
rect 134918 99772 134960 99812
rect 134632 99763 135000 99772
rect 149752 99812 150120 99821
rect 149792 99772 149834 99812
rect 149874 99772 149916 99812
rect 149956 99772 149998 99812
rect 150038 99772 150080 99812
rect 149752 99763 150120 99772
rect 105632 99056 106000 99065
rect 105672 99016 105714 99056
rect 105754 99016 105796 99056
rect 105836 99016 105878 99056
rect 105918 99016 105960 99056
rect 105632 99007 106000 99016
rect 120752 99056 121120 99065
rect 120792 99016 120834 99056
rect 120874 99016 120916 99056
rect 120956 99016 120998 99056
rect 121038 99016 121080 99056
rect 120752 99007 121120 99016
rect 135872 99056 136240 99065
rect 135912 99016 135954 99056
rect 135994 99016 136036 99056
rect 136076 99016 136118 99056
rect 136158 99016 136200 99056
rect 135872 99007 136240 99016
rect 150992 99056 151360 99065
rect 151032 99016 151074 99056
rect 151114 99016 151156 99056
rect 151196 99016 151238 99056
rect 151278 99016 151320 99056
rect 150992 99007 151360 99016
rect 104392 98300 104760 98309
rect 104432 98260 104474 98300
rect 104514 98260 104556 98300
rect 104596 98260 104638 98300
rect 104678 98260 104720 98300
rect 104392 98251 104760 98260
rect 119512 98300 119880 98309
rect 119552 98260 119594 98300
rect 119634 98260 119676 98300
rect 119716 98260 119758 98300
rect 119798 98260 119840 98300
rect 119512 98251 119880 98260
rect 134632 98300 135000 98309
rect 134672 98260 134714 98300
rect 134754 98260 134796 98300
rect 134836 98260 134878 98300
rect 134918 98260 134960 98300
rect 134632 98251 135000 98260
rect 149752 98300 150120 98309
rect 149792 98260 149834 98300
rect 149874 98260 149916 98300
rect 149956 98260 149998 98300
rect 150038 98260 150080 98300
rect 149752 98251 150120 98260
rect 105632 97544 106000 97553
rect 105672 97504 105714 97544
rect 105754 97504 105796 97544
rect 105836 97504 105878 97544
rect 105918 97504 105960 97544
rect 105632 97495 106000 97504
rect 120752 97544 121120 97553
rect 120792 97504 120834 97544
rect 120874 97504 120916 97544
rect 120956 97504 120998 97544
rect 121038 97504 121080 97544
rect 120752 97495 121120 97504
rect 135872 97544 136240 97553
rect 135912 97504 135954 97544
rect 135994 97504 136036 97544
rect 136076 97504 136118 97544
rect 136158 97504 136200 97544
rect 135872 97495 136240 97504
rect 150992 97544 151360 97553
rect 151032 97504 151074 97544
rect 151114 97504 151156 97544
rect 151196 97504 151238 97544
rect 151278 97504 151320 97544
rect 150992 97495 151360 97504
rect 104392 96788 104760 96797
rect 104432 96748 104474 96788
rect 104514 96748 104556 96788
rect 104596 96748 104638 96788
rect 104678 96748 104720 96788
rect 104392 96739 104760 96748
rect 119512 96788 119880 96797
rect 119552 96748 119594 96788
rect 119634 96748 119676 96788
rect 119716 96748 119758 96788
rect 119798 96748 119840 96788
rect 119512 96739 119880 96748
rect 134632 96788 135000 96797
rect 134672 96748 134714 96788
rect 134754 96748 134796 96788
rect 134836 96748 134878 96788
rect 134918 96748 134960 96788
rect 134632 96739 135000 96748
rect 149752 96788 150120 96797
rect 149792 96748 149834 96788
rect 149874 96748 149916 96788
rect 149956 96748 149998 96788
rect 150038 96748 150080 96788
rect 149752 96739 150120 96748
rect 105632 96032 106000 96041
rect 105672 95992 105714 96032
rect 105754 95992 105796 96032
rect 105836 95992 105878 96032
rect 105918 95992 105960 96032
rect 105632 95983 106000 95992
rect 120752 96032 121120 96041
rect 120792 95992 120834 96032
rect 120874 95992 120916 96032
rect 120956 95992 120998 96032
rect 121038 95992 121080 96032
rect 120752 95983 121120 95992
rect 135872 96032 136240 96041
rect 135912 95992 135954 96032
rect 135994 95992 136036 96032
rect 136076 95992 136118 96032
rect 136158 95992 136200 96032
rect 135872 95983 136240 95992
rect 150992 96032 151360 96041
rect 151032 95992 151074 96032
rect 151114 95992 151156 96032
rect 151196 95992 151238 96032
rect 151278 95992 151320 96032
rect 150992 95983 151360 95992
rect 104392 95276 104760 95285
rect 104432 95236 104474 95276
rect 104514 95236 104556 95276
rect 104596 95236 104638 95276
rect 104678 95236 104720 95276
rect 104392 95227 104760 95236
rect 119512 95276 119880 95285
rect 119552 95236 119594 95276
rect 119634 95236 119676 95276
rect 119716 95236 119758 95276
rect 119798 95236 119840 95276
rect 119512 95227 119880 95236
rect 134632 95276 135000 95285
rect 134672 95236 134714 95276
rect 134754 95236 134796 95276
rect 134836 95236 134878 95276
rect 134918 95236 134960 95276
rect 134632 95227 135000 95236
rect 149752 95276 150120 95285
rect 149792 95236 149834 95276
rect 149874 95236 149916 95276
rect 149956 95236 149998 95276
rect 150038 95236 150080 95276
rect 149752 95227 150120 95236
rect 105632 94520 106000 94529
rect 105672 94480 105714 94520
rect 105754 94480 105796 94520
rect 105836 94480 105878 94520
rect 105918 94480 105960 94520
rect 105632 94471 106000 94480
rect 120752 94520 121120 94529
rect 120792 94480 120834 94520
rect 120874 94480 120916 94520
rect 120956 94480 120998 94520
rect 121038 94480 121080 94520
rect 120752 94471 121120 94480
rect 135872 94520 136240 94529
rect 135912 94480 135954 94520
rect 135994 94480 136036 94520
rect 136076 94480 136118 94520
rect 136158 94480 136200 94520
rect 135872 94471 136240 94480
rect 150992 94520 151360 94529
rect 151032 94480 151074 94520
rect 151114 94480 151156 94520
rect 151196 94480 151238 94520
rect 151278 94480 151320 94520
rect 150992 94471 151360 94480
rect 104392 93764 104760 93773
rect 104432 93724 104474 93764
rect 104514 93724 104556 93764
rect 104596 93724 104638 93764
rect 104678 93724 104720 93764
rect 104392 93715 104760 93724
rect 119512 93764 119880 93773
rect 119552 93724 119594 93764
rect 119634 93724 119676 93764
rect 119716 93724 119758 93764
rect 119798 93724 119840 93764
rect 119512 93715 119880 93724
rect 134632 93764 135000 93773
rect 134672 93724 134714 93764
rect 134754 93724 134796 93764
rect 134836 93724 134878 93764
rect 134918 93724 134960 93764
rect 134632 93715 135000 93724
rect 149752 93764 150120 93773
rect 149792 93724 149834 93764
rect 149874 93724 149916 93764
rect 149956 93724 149998 93764
rect 150038 93724 150080 93764
rect 149752 93715 150120 93724
rect 105632 93008 106000 93017
rect 105672 92968 105714 93008
rect 105754 92968 105796 93008
rect 105836 92968 105878 93008
rect 105918 92968 105960 93008
rect 105632 92959 106000 92968
rect 120752 93008 121120 93017
rect 120792 92968 120834 93008
rect 120874 92968 120916 93008
rect 120956 92968 120998 93008
rect 121038 92968 121080 93008
rect 120752 92959 121120 92968
rect 135872 93008 136240 93017
rect 135912 92968 135954 93008
rect 135994 92968 136036 93008
rect 136076 92968 136118 93008
rect 136158 92968 136200 93008
rect 135872 92959 136240 92968
rect 150992 93008 151360 93017
rect 151032 92968 151074 93008
rect 151114 92968 151156 93008
rect 151196 92968 151238 93008
rect 151278 92968 151320 93008
rect 150992 92959 151360 92968
rect 104392 92252 104760 92261
rect 104432 92212 104474 92252
rect 104514 92212 104556 92252
rect 104596 92212 104638 92252
rect 104678 92212 104720 92252
rect 104392 92203 104760 92212
rect 119512 92252 119880 92261
rect 119552 92212 119594 92252
rect 119634 92212 119676 92252
rect 119716 92212 119758 92252
rect 119798 92212 119840 92252
rect 119512 92203 119880 92212
rect 134632 92252 135000 92261
rect 134672 92212 134714 92252
rect 134754 92212 134796 92252
rect 134836 92212 134878 92252
rect 134918 92212 134960 92252
rect 134632 92203 135000 92212
rect 149752 92252 150120 92261
rect 149792 92212 149834 92252
rect 149874 92212 149916 92252
rect 149956 92212 149998 92252
rect 150038 92212 150080 92252
rect 149752 92203 150120 92212
rect 105632 91496 106000 91505
rect 105672 91456 105714 91496
rect 105754 91456 105796 91496
rect 105836 91456 105878 91496
rect 105918 91456 105960 91496
rect 105632 91447 106000 91456
rect 120752 91496 121120 91505
rect 120792 91456 120834 91496
rect 120874 91456 120916 91496
rect 120956 91456 120998 91496
rect 121038 91456 121080 91496
rect 120752 91447 121120 91456
rect 135872 91496 136240 91505
rect 135912 91456 135954 91496
rect 135994 91456 136036 91496
rect 136076 91456 136118 91496
rect 136158 91456 136200 91496
rect 135872 91447 136240 91456
rect 150992 91496 151360 91505
rect 151032 91456 151074 91496
rect 151114 91456 151156 91496
rect 151196 91456 151238 91496
rect 151278 91456 151320 91496
rect 150992 91447 151360 91456
rect 104392 90740 104760 90749
rect 104432 90700 104474 90740
rect 104514 90700 104556 90740
rect 104596 90700 104638 90740
rect 104678 90700 104720 90740
rect 104392 90691 104760 90700
rect 119512 90740 119880 90749
rect 119552 90700 119594 90740
rect 119634 90700 119676 90740
rect 119716 90700 119758 90740
rect 119798 90700 119840 90740
rect 119512 90691 119880 90700
rect 134632 90740 135000 90749
rect 134672 90700 134714 90740
rect 134754 90700 134796 90740
rect 134836 90700 134878 90740
rect 134918 90700 134960 90740
rect 134632 90691 135000 90700
rect 149752 90740 150120 90749
rect 149792 90700 149834 90740
rect 149874 90700 149916 90740
rect 149956 90700 149998 90740
rect 150038 90700 150080 90740
rect 149752 90691 150120 90700
rect 105632 89984 106000 89993
rect 105672 89944 105714 89984
rect 105754 89944 105796 89984
rect 105836 89944 105878 89984
rect 105918 89944 105960 89984
rect 105632 89935 106000 89944
rect 120752 89984 121120 89993
rect 120792 89944 120834 89984
rect 120874 89944 120916 89984
rect 120956 89944 120998 89984
rect 121038 89944 121080 89984
rect 120752 89935 121120 89944
rect 135872 89984 136240 89993
rect 135912 89944 135954 89984
rect 135994 89944 136036 89984
rect 136076 89944 136118 89984
rect 136158 89944 136200 89984
rect 135872 89935 136240 89944
rect 150992 89984 151360 89993
rect 151032 89944 151074 89984
rect 151114 89944 151156 89984
rect 151196 89944 151238 89984
rect 151278 89944 151320 89984
rect 150992 89935 151360 89944
rect 104392 89228 104760 89237
rect 104432 89188 104474 89228
rect 104514 89188 104556 89228
rect 104596 89188 104638 89228
rect 104678 89188 104720 89228
rect 104392 89179 104760 89188
rect 119512 89228 119880 89237
rect 119552 89188 119594 89228
rect 119634 89188 119676 89228
rect 119716 89188 119758 89228
rect 119798 89188 119840 89228
rect 119512 89179 119880 89188
rect 134632 89228 135000 89237
rect 134672 89188 134714 89228
rect 134754 89188 134796 89228
rect 134836 89188 134878 89228
rect 134918 89188 134960 89228
rect 134632 89179 135000 89188
rect 149752 89228 150120 89237
rect 149792 89188 149834 89228
rect 149874 89188 149916 89228
rect 149956 89188 149998 89228
rect 150038 89188 150080 89228
rect 149752 89179 150120 89188
rect 105632 88472 106000 88481
rect 105672 88432 105714 88472
rect 105754 88432 105796 88472
rect 105836 88432 105878 88472
rect 105918 88432 105960 88472
rect 105632 88423 106000 88432
rect 120752 88472 121120 88481
rect 120792 88432 120834 88472
rect 120874 88432 120916 88472
rect 120956 88432 120998 88472
rect 121038 88432 121080 88472
rect 120752 88423 121120 88432
rect 135872 88472 136240 88481
rect 135912 88432 135954 88472
rect 135994 88432 136036 88472
rect 136076 88432 136118 88472
rect 136158 88432 136200 88472
rect 135872 88423 136240 88432
rect 150992 88472 151360 88481
rect 151032 88432 151074 88472
rect 151114 88432 151156 88472
rect 151196 88432 151238 88472
rect 151278 88432 151320 88472
rect 150992 88423 151360 88432
rect 104392 87716 104760 87725
rect 104432 87676 104474 87716
rect 104514 87676 104556 87716
rect 104596 87676 104638 87716
rect 104678 87676 104720 87716
rect 104392 87667 104760 87676
rect 119512 87716 119880 87725
rect 119552 87676 119594 87716
rect 119634 87676 119676 87716
rect 119716 87676 119758 87716
rect 119798 87676 119840 87716
rect 119512 87667 119880 87676
rect 134632 87716 135000 87725
rect 134672 87676 134714 87716
rect 134754 87676 134796 87716
rect 134836 87676 134878 87716
rect 134918 87676 134960 87716
rect 134632 87667 135000 87676
rect 149752 87716 150120 87725
rect 149792 87676 149834 87716
rect 149874 87676 149916 87716
rect 149956 87676 149998 87716
rect 150038 87676 150080 87716
rect 149752 87667 150120 87676
rect 105632 86960 106000 86969
rect 105672 86920 105714 86960
rect 105754 86920 105796 86960
rect 105836 86920 105878 86960
rect 105918 86920 105960 86960
rect 105632 86911 106000 86920
rect 120752 86960 121120 86969
rect 120792 86920 120834 86960
rect 120874 86920 120916 86960
rect 120956 86920 120998 86960
rect 121038 86920 121080 86960
rect 120752 86911 121120 86920
rect 135872 86960 136240 86969
rect 135912 86920 135954 86960
rect 135994 86920 136036 86960
rect 136076 86920 136118 86960
rect 136158 86920 136200 86960
rect 135872 86911 136240 86920
rect 150992 86960 151360 86969
rect 151032 86920 151074 86960
rect 151114 86920 151156 86960
rect 151196 86920 151238 86960
rect 151278 86920 151320 86960
rect 150992 86911 151360 86920
rect 104392 86204 104760 86213
rect 104432 86164 104474 86204
rect 104514 86164 104556 86204
rect 104596 86164 104638 86204
rect 104678 86164 104720 86204
rect 104392 86155 104760 86164
rect 119512 86204 119880 86213
rect 119552 86164 119594 86204
rect 119634 86164 119676 86204
rect 119716 86164 119758 86204
rect 119798 86164 119840 86204
rect 119512 86155 119880 86164
rect 134632 86204 135000 86213
rect 134672 86164 134714 86204
rect 134754 86164 134796 86204
rect 134836 86164 134878 86204
rect 134918 86164 134960 86204
rect 134632 86155 135000 86164
rect 149752 86204 150120 86213
rect 149792 86164 149834 86204
rect 149874 86164 149916 86204
rect 149956 86164 149998 86204
rect 150038 86164 150080 86204
rect 149752 86155 150120 86164
rect 105632 85448 106000 85457
rect 105672 85408 105714 85448
rect 105754 85408 105796 85448
rect 105836 85408 105878 85448
rect 105918 85408 105960 85448
rect 105632 85399 106000 85408
rect 120752 85448 121120 85457
rect 120792 85408 120834 85448
rect 120874 85408 120916 85448
rect 120956 85408 120998 85448
rect 121038 85408 121080 85448
rect 120752 85399 121120 85408
rect 135872 85448 136240 85457
rect 135912 85408 135954 85448
rect 135994 85408 136036 85448
rect 136076 85408 136118 85448
rect 136158 85408 136200 85448
rect 135872 85399 136240 85408
rect 150992 85448 151360 85457
rect 151032 85408 151074 85448
rect 151114 85408 151156 85448
rect 151196 85408 151238 85448
rect 151278 85408 151320 85448
rect 150992 85399 151360 85408
rect 104392 84692 104760 84701
rect 104432 84652 104474 84692
rect 104514 84652 104556 84692
rect 104596 84652 104638 84692
rect 104678 84652 104720 84692
rect 104392 84643 104760 84652
rect 119512 84692 119880 84701
rect 119552 84652 119594 84692
rect 119634 84652 119676 84692
rect 119716 84652 119758 84692
rect 119798 84652 119840 84692
rect 119512 84643 119880 84652
rect 134632 84692 135000 84701
rect 134672 84652 134714 84692
rect 134754 84652 134796 84692
rect 134836 84652 134878 84692
rect 134918 84652 134960 84692
rect 134632 84643 135000 84652
rect 149752 84692 150120 84701
rect 149792 84652 149834 84692
rect 149874 84652 149916 84692
rect 149956 84652 149998 84692
rect 150038 84652 150080 84692
rect 149752 84643 150120 84652
rect 105632 83936 106000 83945
rect 105672 83896 105714 83936
rect 105754 83896 105796 83936
rect 105836 83896 105878 83936
rect 105918 83896 105960 83936
rect 105632 83887 106000 83896
rect 120752 83936 121120 83945
rect 120792 83896 120834 83936
rect 120874 83896 120916 83936
rect 120956 83896 120998 83936
rect 121038 83896 121080 83936
rect 120752 83887 121120 83896
rect 135872 83936 136240 83945
rect 135912 83896 135954 83936
rect 135994 83896 136036 83936
rect 136076 83896 136118 83936
rect 136158 83896 136200 83936
rect 135872 83887 136240 83896
rect 150992 83936 151360 83945
rect 151032 83896 151074 83936
rect 151114 83896 151156 83936
rect 151196 83896 151238 83936
rect 151278 83896 151320 83936
rect 150992 83887 151360 83896
rect 104392 83180 104760 83189
rect 104432 83140 104474 83180
rect 104514 83140 104556 83180
rect 104596 83140 104638 83180
rect 104678 83140 104720 83180
rect 104392 83131 104760 83140
rect 119512 83180 119880 83189
rect 119552 83140 119594 83180
rect 119634 83140 119676 83180
rect 119716 83140 119758 83180
rect 119798 83140 119840 83180
rect 119512 83131 119880 83140
rect 134632 83180 135000 83189
rect 134672 83140 134714 83180
rect 134754 83140 134796 83180
rect 134836 83140 134878 83180
rect 134918 83140 134960 83180
rect 134632 83131 135000 83140
rect 149752 83180 150120 83189
rect 149792 83140 149834 83180
rect 149874 83140 149916 83180
rect 149956 83140 149998 83180
rect 150038 83140 150080 83180
rect 149752 83131 150120 83140
rect 105632 82424 106000 82433
rect 105672 82384 105714 82424
rect 105754 82384 105796 82424
rect 105836 82384 105878 82424
rect 105918 82384 105960 82424
rect 105632 82375 106000 82384
rect 120752 82424 121120 82433
rect 120792 82384 120834 82424
rect 120874 82384 120916 82424
rect 120956 82384 120998 82424
rect 121038 82384 121080 82424
rect 120752 82375 121120 82384
rect 135872 82424 136240 82433
rect 135912 82384 135954 82424
rect 135994 82384 136036 82424
rect 136076 82384 136118 82424
rect 136158 82384 136200 82424
rect 135872 82375 136240 82384
rect 150992 82424 151360 82433
rect 151032 82384 151074 82424
rect 151114 82384 151156 82424
rect 151196 82384 151238 82424
rect 151278 82384 151320 82424
rect 150992 82375 151360 82384
rect 104392 81668 104760 81677
rect 104432 81628 104474 81668
rect 104514 81628 104556 81668
rect 104596 81628 104638 81668
rect 104678 81628 104720 81668
rect 104392 81619 104760 81628
rect 119512 81668 119880 81677
rect 119552 81628 119594 81668
rect 119634 81628 119676 81668
rect 119716 81628 119758 81668
rect 119798 81628 119840 81668
rect 119512 81619 119880 81628
rect 134632 81668 135000 81677
rect 134672 81628 134714 81668
rect 134754 81628 134796 81668
rect 134836 81628 134878 81668
rect 134918 81628 134960 81668
rect 134632 81619 135000 81628
rect 149752 81668 150120 81677
rect 149792 81628 149834 81668
rect 149874 81628 149916 81668
rect 149956 81628 149998 81668
rect 150038 81628 150080 81668
rect 149752 81619 150120 81628
rect 105632 80912 106000 80921
rect 105672 80872 105714 80912
rect 105754 80872 105796 80912
rect 105836 80872 105878 80912
rect 105918 80872 105960 80912
rect 105632 80863 106000 80872
rect 120752 80912 121120 80921
rect 120792 80872 120834 80912
rect 120874 80872 120916 80912
rect 120956 80872 120998 80912
rect 121038 80872 121080 80912
rect 120752 80863 121120 80872
rect 135872 80912 136240 80921
rect 135912 80872 135954 80912
rect 135994 80872 136036 80912
rect 136076 80872 136118 80912
rect 136158 80872 136200 80912
rect 135872 80863 136240 80872
rect 150992 80912 151360 80921
rect 151032 80872 151074 80912
rect 151114 80872 151156 80912
rect 151196 80872 151238 80912
rect 151278 80872 151320 80912
rect 150992 80863 151360 80872
rect 104392 80156 104760 80165
rect 104432 80116 104474 80156
rect 104514 80116 104556 80156
rect 104596 80116 104638 80156
rect 104678 80116 104720 80156
rect 104392 80107 104760 80116
rect 119512 80156 119880 80165
rect 119552 80116 119594 80156
rect 119634 80116 119676 80156
rect 119716 80116 119758 80156
rect 119798 80116 119840 80156
rect 119512 80107 119880 80116
rect 134632 80156 135000 80165
rect 134672 80116 134714 80156
rect 134754 80116 134796 80156
rect 134836 80116 134878 80156
rect 134918 80116 134960 80156
rect 134632 80107 135000 80116
rect 149752 80156 150120 80165
rect 149792 80116 149834 80156
rect 149874 80116 149916 80156
rect 149956 80116 149998 80156
rect 150038 80116 150080 80156
rect 149752 80107 150120 80116
rect 105632 79400 106000 79409
rect 105672 79360 105714 79400
rect 105754 79360 105796 79400
rect 105836 79360 105878 79400
rect 105918 79360 105960 79400
rect 105632 79351 106000 79360
rect 120752 79400 121120 79409
rect 120792 79360 120834 79400
rect 120874 79360 120916 79400
rect 120956 79360 120998 79400
rect 121038 79360 121080 79400
rect 120752 79351 121120 79360
rect 135872 79400 136240 79409
rect 135912 79360 135954 79400
rect 135994 79360 136036 79400
rect 136076 79360 136118 79400
rect 136158 79360 136200 79400
rect 135872 79351 136240 79360
rect 150992 79400 151360 79409
rect 151032 79360 151074 79400
rect 151114 79360 151156 79400
rect 151196 79360 151238 79400
rect 151278 79360 151320 79400
rect 150992 79351 151360 79360
rect 104392 78644 104760 78653
rect 104432 78604 104474 78644
rect 104514 78604 104556 78644
rect 104596 78604 104638 78644
rect 104678 78604 104720 78644
rect 104392 78595 104760 78604
rect 119512 78644 119880 78653
rect 119552 78604 119594 78644
rect 119634 78604 119676 78644
rect 119716 78604 119758 78644
rect 119798 78604 119840 78644
rect 119512 78595 119880 78604
rect 134632 78644 135000 78653
rect 134672 78604 134714 78644
rect 134754 78604 134796 78644
rect 134836 78604 134878 78644
rect 134918 78604 134960 78644
rect 134632 78595 135000 78604
rect 149752 78644 150120 78653
rect 149792 78604 149834 78644
rect 149874 78604 149916 78644
rect 149956 78604 149998 78644
rect 150038 78604 150080 78644
rect 149752 78595 150120 78604
rect 105632 77888 106000 77897
rect 105672 77848 105714 77888
rect 105754 77848 105796 77888
rect 105836 77848 105878 77888
rect 105918 77848 105960 77888
rect 105632 77839 106000 77848
rect 120752 77888 121120 77897
rect 120792 77848 120834 77888
rect 120874 77848 120916 77888
rect 120956 77848 120998 77888
rect 121038 77848 121080 77888
rect 120752 77839 121120 77848
rect 135872 77888 136240 77897
rect 135912 77848 135954 77888
rect 135994 77848 136036 77888
rect 136076 77848 136118 77888
rect 136158 77848 136200 77888
rect 135872 77839 136240 77848
rect 150992 77888 151360 77897
rect 151032 77848 151074 77888
rect 151114 77848 151156 77888
rect 151196 77848 151238 77888
rect 151278 77848 151320 77888
rect 150992 77839 151360 77848
rect 104392 77132 104760 77141
rect 104432 77092 104474 77132
rect 104514 77092 104556 77132
rect 104596 77092 104638 77132
rect 104678 77092 104720 77132
rect 104392 77083 104760 77092
rect 119512 77132 119880 77141
rect 119552 77092 119594 77132
rect 119634 77092 119676 77132
rect 119716 77092 119758 77132
rect 119798 77092 119840 77132
rect 119512 77083 119880 77092
rect 134632 77132 135000 77141
rect 134672 77092 134714 77132
rect 134754 77092 134796 77132
rect 134836 77092 134878 77132
rect 134918 77092 134960 77132
rect 134632 77083 135000 77092
rect 149752 77132 150120 77141
rect 149792 77092 149834 77132
rect 149874 77092 149916 77132
rect 149956 77092 149998 77132
rect 150038 77092 150080 77132
rect 149752 77083 150120 77092
rect 105632 76376 106000 76385
rect 105672 76336 105714 76376
rect 105754 76336 105796 76376
rect 105836 76336 105878 76376
rect 105918 76336 105960 76376
rect 105632 76327 106000 76336
rect 120752 76376 121120 76385
rect 120792 76336 120834 76376
rect 120874 76336 120916 76376
rect 120956 76336 120998 76376
rect 121038 76336 121080 76376
rect 120752 76327 121120 76336
rect 135872 76376 136240 76385
rect 135912 76336 135954 76376
rect 135994 76336 136036 76376
rect 136076 76336 136118 76376
rect 136158 76336 136200 76376
rect 135872 76327 136240 76336
rect 150992 76376 151360 76385
rect 151032 76336 151074 76376
rect 151114 76336 151156 76376
rect 151196 76336 151238 76376
rect 151278 76336 151320 76376
rect 150992 76327 151360 76336
rect 104392 75620 104760 75629
rect 104432 75580 104474 75620
rect 104514 75580 104556 75620
rect 104596 75580 104638 75620
rect 104678 75580 104720 75620
rect 104392 75571 104760 75580
rect 119512 75620 119880 75629
rect 119552 75580 119594 75620
rect 119634 75580 119676 75620
rect 119716 75580 119758 75620
rect 119798 75580 119840 75620
rect 119512 75571 119880 75580
rect 134632 75620 135000 75629
rect 134672 75580 134714 75620
rect 134754 75580 134796 75620
rect 134836 75580 134878 75620
rect 134918 75580 134960 75620
rect 134632 75571 135000 75580
rect 149752 75620 150120 75629
rect 149792 75580 149834 75620
rect 149874 75580 149916 75620
rect 149956 75580 149998 75620
rect 150038 75580 150080 75620
rect 149752 75571 150120 75580
rect 105632 74864 106000 74873
rect 105672 74824 105714 74864
rect 105754 74824 105796 74864
rect 105836 74824 105878 74864
rect 105918 74824 105960 74864
rect 105632 74815 106000 74824
rect 120752 74864 121120 74873
rect 120792 74824 120834 74864
rect 120874 74824 120916 74864
rect 120956 74824 120998 74864
rect 121038 74824 121080 74864
rect 120752 74815 121120 74824
rect 135872 74864 136240 74873
rect 135912 74824 135954 74864
rect 135994 74824 136036 74864
rect 136076 74824 136118 74864
rect 136158 74824 136200 74864
rect 135872 74815 136240 74824
rect 150992 74864 151360 74873
rect 151032 74824 151074 74864
rect 151114 74824 151156 74864
rect 151196 74824 151238 74864
rect 151278 74824 151320 74864
rect 150992 74815 151360 74824
rect 104392 74108 104760 74117
rect 104432 74068 104474 74108
rect 104514 74068 104556 74108
rect 104596 74068 104638 74108
rect 104678 74068 104720 74108
rect 104392 74059 104760 74068
rect 119512 74108 119880 74117
rect 119552 74068 119594 74108
rect 119634 74068 119676 74108
rect 119716 74068 119758 74108
rect 119798 74068 119840 74108
rect 119512 74059 119880 74068
rect 134632 74108 135000 74117
rect 134672 74068 134714 74108
rect 134754 74068 134796 74108
rect 134836 74068 134878 74108
rect 134918 74068 134960 74108
rect 134632 74059 135000 74068
rect 149752 74108 150120 74117
rect 149792 74068 149834 74108
rect 149874 74068 149916 74108
rect 149956 74068 149998 74108
rect 150038 74068 150080 74108
rect 149752 74059 150120 74068
rect 105632 73352 106000 73361
rect 105672 73312 105714 73352
rect 105754 73312 105796 73352
rect 105836 73312 105878 73352
rect 105918 73312 105960 73352
rect 105632 73303 106000 73312
rect 120752 73352 121120 73361
rect 120792 73312 120834 73352
rect 120874 73312 120916 73352
rect 120956 73312 120998 73352
rect 121038 73312 121080 73352
rect 120752 73303 121120 73312
rect 135872 73352 136240 73361
rect 135912 73312 135954 73352
rect 135994 73312 136036 73352
rect 136076 73312 136118 73352
rect 136158 73312 136200 73352
rect 135872 73303 136240 73312
rect 150992 73352 151360 73361
rect 151032 73312 151074 73352
rect 151114 73312 151156 73352
rect 151196 73312 151238 73352
rect 151278 73312 151320 73352
rect 150992 73303 151360 73312
rect 104392 72596 104760 72605
rect 104432 72556 104474 72596
rect 104514 72556 104556 72596
rect 104596 72556 104638 72596
rect 104678 72556 104720 72596
rect 104392 72547 104760 72556
rect 119512 72596 119880 72605
rect 119552 72556 119594 72596
rect 119634 72556 119676 72596
rect 119716 72556 119758 72596
rect 119798 72556 119840 72596
rect 119512 72547 119880 72556
rect 134632 72596 135000 72605
rect 134672 72556 134714 72596
rect 134754 72556 134796 72596
rect 134836 72556 134878 72596
rect 134918 72556 134960 72596
rect 134632 72547 135000 72556
rect 149752 72596 150120 72605
rect 149792 72556 149834 72596
rect 149874 72556 149916 72596
rect 149956 72556 149998 72596
rect 150038 72556 150080 72596
rect 149752 72547 150120 72556
rect 105632 71840 106000 71849
rect 105672 71800 105714 71840
rect 105754 71800 105796 71840
rect 105836 71800 105878 71840
rect 105918 71800 105960 71840
rect 105632 71791 106000 71800
rect 120752 71840 121120 71849
rect 120792 71800 120834 71840
rect 120874 71800 120916 71840
rect 120956 71800 120998 71840
rect 121038 71800 121080 71840
rect 120752 71791 121120 71800
rect 135872 71840 136240 71849
rect 135912 71800 135954 71840
rect 135994 71800 136036 71840
rect 136076 71800 136118 71840
rect 136158 71800 136200 71840
rect 135872 71791 136240 71800
rect 150992 71840 151360 71849
rect 151032 71800 151074 71840
rect 151114 71800 151156 71840
rect 151196 71800 151238 71840
rect 151278 71800 151320 71840
rect 150992 71791 151360 71800
rect 71975 64324 72020 64364
rect 87975 64324 88052 64364
rect 103975 64324 104084 64364
rect 71975 63966 72015 64324
rect 87975 63966 88015 64324
rect 103975 63966 104015 64324
rect 151564 64205 151604 158740
rect 151563 64196 151605 64205
rect 151563 64156 151564 64196
rect 151604 64156 151605 64196
rect 151563 64147 151605 64156
<< via2 >>
rect 71980 159412 72020 159452
rect 103660 159412 103700 159452
rect 104044 159412 104084 159452
rect 64108 152020 64148 152060
rect 64108 135976 64148 136016
rect 64108 120016 64148 120056
rect 64108 103972 64148 104012
rect 64108 88012 64148 88052
rect 64108 71968 64148 72008
rect 88012 159328 88052 159368
rect 75392 151936 75432 151976
rect 75474 151936 75514 151976
rect 75556 151936 75596 151976
rect 75638 151936 75678 151976
rect 75720 151936 75760 151976
rect 74152 151180 74192 151220
rect 74234 151180 74274 151220
rect 74316 151180 74356 151220
rect 74398 151180 74438 151220
rect 74480 151180 74520 151220
rect 75392 150424 75432 150464
rect 75474 150424 75514 150464
rect 75556 150424 75596 150464
rect 75638 150424 75678 150464
rect 75720 150424 75760 150464
rect 74152 149668 74192 149708
rect 74234 149668 74274 149708
rect 74316 149668 74356 149708
rect 74398 149668 74438 149708
rect 74480 149668 74520 149708
rect 75392 148912 75432 148952
rect 75474 148912 75514 148952
rect 75556 148912 75596 148952
rect 75638 148912 75678 148952
rect 75720 148912 75760 148952
rect 74152 148156 74192 148196
rect 74234 148156 74274 148196
rect 74316 148156 74356 148196
rect 74398 148156 74438 148196
rect 74480 148156 74520 148196
rect 75392 147400 75432 147440
rect 75474 147400 75514 147440
rect 75556 147400 75596 147440
rect 75638 147400 75678 147440
rect 75720 147400 75760 147440
rect 74152 146644 74192 146684
rect 74234 146644 74274 146684
rect 74316 146644 74356 146684
rect 74398 146644 74438 146684
rect 74480 146644 74520 146684
rect 75392 145888 75432 145928
rect 75474 145888 75514 145928
rect 75556 145888 75596 145928
rect 75638 145888 75678 145928
rect 75720 145888 75760 145928
rect 74152 145132 74192 145172
rect 74234 145132 74274 145172
rect 74316 145132 74356 145172
rect 74398 145132 74438 145172
rect 74480 145132 74520 145172
rect 75392 144376 75432 144416
rect 75474 144376 75514 144416
rect 75556 144376 75596 144416
rect 75638 144376 75678 144416
rect 75720 144376 75760 144416
rect 74152 143620 74192 143660
rect 74234 143620 74274 143660
rect 74316 143620 74356 143660
rect 74398 143620 74438 143660
rect 74480 143620 74520 143660
rect 75392 142864 75432 142904
rect 75474 142864 75514 142904
rect 75556 142864 75596 142904
rect 75638 142864 75678 142904
rect 75720 142864 75760 142904
rect 74152 142108 74192 142148
rect 74234 142108 74274 142148
rect 74316 142108 74356 142148
rect 74398 142108 74438 142148
rect 74480 142108 74520 142148
rect 75392 141352 75432 141392
rect 75474 141352 75514 141392
rect 75556 141352 75596 141392
rect 75638 141352 75678 141392
rect 75720 141352 75760 141392
rect 74152 140596 74192 140636
rect 74234 140596 74274 140636
rect 74316 140596 74356 140636
rect 74398 140596 74438 140636
rect 74480 140596 74520 140636
rect 75392 139840 75432 139880
rect 75474 139840 75514 139880
rect 75556 139840 75596 139880
rect 75638 139840 75678 139880
rect 75720 139840 75760 139880
rect 74152 139084 74192 139124
rect 74234 139084 74274 139124
rect 74316 139084 74356 139124
rect 74398 139084 74438 139124
rect 74480 139084 74520 139124
rect 75392 138328 75432 138368
rect 75474 138328 75514 138368
rect 75556 138328 75596 138368
rect 75638 138328 75678 138368
rect 75720 138328 75760 138368
rect 74152 137572 74192 137612
rect 74234 137572 74274 137612
rect 74316 137572 74356 137612
rect 74398 137572 74438 137612
rect 74480 137572 74520 137612
rect 75392 136816 75432 136856
rect 75474 136816 75514 136856
rect 75556 136816 75596 136856
rect 75638 136816 75678 136856
rect 75720 136816 75760 136856
rect 74152 136060 74192 136100
rect 74234 136060 74274 136100
rect 74316 136060 74356 136100
rect 74398 136060 74438 136100
rect 74480 136060 74520 136100
rect 75392 135304 75432 135344
rect 75474 135304 75514 135344
rect 75556 135304 75596 135344
rect 75638 135304 75678 135344
rect 75720 135304 75760 135344
rect 74152 134548 74192 134588
rect 74234 134548 74274 134588
rect 74316 134548 74356 134588
rect 74398 134548 74438 134588
rect 74480 134548 74520 134588
rect 75392 133792 75432 133832
rect 75474 133792 75514 133832
rect 75556 133792 75596 133832
rect 75638 133792 75678 133832
rect 75720 133792 75760 133832
rect 74152 133036 74192 133076
rect 74234 133036 74274 133076
rect 74316 133036 74356 133076
rect 74398 133036 74438 133076
rect 74480 133036 74520 133076
rect 75392 132280 75432 132320
rect 75474 132280 75514 132320
rect 75556 132280 75596 132320
rect 75638 132280 75678 132320
rect 75720 132280 75760 132320
rect 74152 131524 74192 131564
rect 74234 131524 74274 131564
rect 74316 131524 74356 131564
rect 74398 131524 74438 131564
rect 74480 131524 74520 131564
rect 75392 130768 75432 130808
rect 75474 130768 75514 130808
rect 75556 130768 75596 130808
rect 75638 130768 75678 130808
rect 75720 130768 75760 130808
rect 74152 130012 74192 130052
rect 74234 130012 74274 130052
rect 74316 130012 74356 130052
rect 74398 130012 74438 130052
rect 74480 130012 74520 130052
rect 75392 129256 75432 129296
rect 75474 129256 75514 129296
rect 75556 129256 75596 129296
rect 75638 129256 75678 129296
rect 75720 129256 75760 129296
rect 74152 128500 74192 128540
rect 74234 128500 74274 128540
rect 74316 128500 74356 128540
rect 74398 128500 74438 128540
rect 74480 128500 74520 128540
rect 75392 127744 75432 127784
rect 75474 127744 75514 127784
rect 75556 127744 75596 127784
rect 75638 127744 75678 127784
rect 75720 127744 75760 127784
rect 74152 126988 74192 127028
rect 74234 126988 74274 127028
rect 74316 126988 74356 127028
rect 74398 126988 74438 127028
rect 74480 126988 74520 127028
rect 75392 126232 75432 126272
rect 75474 126232 75514 126272
rect 75556 126232 75596 126272
rect 75638 126232 75678 126272
rect 75720 126232 75760 126272
rect 74152 125476 74192 125516
rect 74234 125476 74274 125516
rect 74316 125476 74356 125516
rect 74398 125476 74438 125516
rect 74480 125476 74520 125516
rect 75392 124720 75432 124760
rect 75474 124720 75514 124760
rect 75556 124720 75596 124760
rect 75638 124720 75678 124760
rect 75720 124720 75760 124760
rect 74152 123964 74192 124004
rect 74234 123964 74274 124004
rect 74316 123964 74356 124004
rect 74398 123964 74438 124004
rect 74480 123964 74520 124004
rect 75392 123208 75432 123248
rect 75474 123208 75514 123248
rect 75556 123208 75596 123248
rect 75638 123208 75678 123248
rect 75720 123208 75760 123248
rect 74152 122452 74192 122492
rect 74234 122452 74274 122492
rect 74316 122452 74356 122492
rect 74398 122452 74438 122492
rect 74480 122452 74520 122492
rect 75392 121696 75432 121736
rect 75474 121696 75514 121736
rect 75556 121696 75596 121736
rect 75638 121696 75678 121736
rect 75720 121696 75760 121736
rect 74152 120940 74192 120980
rect 74234 120940 74274 120980
rect 74316 120940 74356 120980
rect 74398 120940 74438 120980
rect 74480 120940 74520 120980
rect 75392 120184 75432 120224
rect 75474 120184 75514 120224
rect 75556 120184 75596 120224
rect 75638 120184 75678 120224
rect 75720 120184 75760 120224
rect 74152 119428 74192 119468
rect 74234 119428 74274 119468
rect 74316 119428 74356 119468
rect 74398 119428 74438 119468
rect 74480 119428 74520 119468
rect 75392 118672 75432 118712
rect 75474 118672 75514 118712
rect 75556 118672 75596 118712
rect 75638 118672 75678 118712
rect 75720 118672 75760 118712
rect 74152 117916 74192 117956
rect 74234 117916 74274 117956
rect 74316 117916 74356 117956
rect 74398 117916 74438 117956
rect 74480 117916 74520 117956
rect 75392 117160 75432 117200
rect 75474 117160 75514 117200
rect 75556 117160 75596 117200
rect 75638 117160 75678 117200
rect 75720 117160 75760 117200
rect 74152 116404 74192 116444
rect 74234 116404 74274 116444
rect 74316 116404 74356 116444
rect 74398 116404 74438 116444
rect 74480 116404 74520 116444
rect 75392 115648 75432 115688
rect 75474 115648 75514 115688
rect 75556 115648 75596 115688
rect 75638 115648 75678 115688
rect 75720 115648 75760 115688
rect 74152 114892 74192 114932
rect 74234 114892 74274 114932
rect 74316 114892 74356 114932
rect 74398 114892 74438 114932
rect 74480 114892 74520 114932
rect 75392 114136 75432 114176
rect 75474 114136 75514 114176
rect 75556 114136 75596 114176
rect 75638 114136 75678 114176
rect 75720 114136 75760 114176
rect 74152 113380 74192 113420
rect 74234 113380 74274 113420
rect 74316 113380 74356 113420
rect 74398 113380 74438 113420
rect 74480 113380 74520 113420
rect 75392 112624 75432 112664
rect 75474 112624 75514 112664
rect 75556 112624 75596 112664
rect 75638 112624 75678 112664
rect 75720 112624 75760 112664
rect 74152 111868 74192 111908
rect 74234 111868 74274 111908
rect 74316 111868 74356 111908
rect 74398 111868 74438 111908
rect 74480 111868 74520 111908
rect 75392 111112 75432 111152
rect 75474 111112 75514 111152
rect 75556 111112 75596 111152
rect 75638 111112 75678 111152
rect 75720 111112 75760 111152
rect 74152 110356 74192 110396
rect 74234 110356 74274 110396
rect 74316 110356 74356 110396
rect 74398 110356 74438 110396
rect 74480 110356 74520 110396
rect 75392 109600 75432 109640
rect 75474 109600 75514 109640
rect 75556 109600 75596 109640
rect 75638 109600 75678 109640
rect 75720 109600 75760 109640
rect 74152 108844 74192 108884
rect 74234 108844 74274 108884
rect 74316 108844 74356 108884
rect 74398 108844 74438 108884
rect 74480 108844 74520 108884
rect 75392 108088 75432 108128
rect 75474 108088 75514 108128
rect 75556 108088 75596 108128
rect 75638 108088 75678 108128
rect 75720 108088 75760 108128
rect 74152 107332 74192 107372
rect 74234 107332 74274 107372
rect 74316 107332 74356 107372
rect 74398 107332 74438 107372
rect 74480 107332 74520 107372
rect 75392 106576 75432 106616
rect 75474 106576 75514 106616
rect 75556 106576 75596 106616
rect 75638 106576 75678 106616
rect 75720 106576 75760 106616
rect 74152 105820 74192 105860
rect 74234 105820 74274 105860
rect 74316 105820 74356 105860
rect 74398 105820 74438 105860
rect 74480 105820 74520 105860
rect 75392 105064 75432 105104
rect 75474 105064 75514 105104
rect 75556 105064 75596 105104
rect 75638 105064 75678 105104
rect 75720 105064 75760 105104
rect 74152 104308 74192 104348
rect 74234 104308 74274 104348
rect 74316 104308 74356 104348
rect 74398 104308 74438 104348
rect 74480 104308 74520 104348
rect 75392 103552 75432 103592
rect 75474 103552 75514 103592
rect 75556 103552 75596 103592
rect 75638 103552 75678 103592
rect 75720 103552 75760 103592
rect 74152 102796 74192 102836
rect 74234 102796 74274 102836
rect 74316 102796 74356 102836
rect 74398 102796 74438 102836
rect 74480 102796 74520 102836
rect 75392 102040 75432 102080
rect 75474 102040 75514 102080
rect 75556 102040 75596 102080
rect 75638 102040 75678 102080
rect 75720 102040 75760 102080
rect 74152 101284 74192 101324
rect 74234 101284 74274 101324
rect 74316 101284 74356 101324
rect 74398 101284 74438 101324
rect 74480 101284 74520 101324
rect 75392 100528 75432 100568
rect 75474 100528 75514 100568
rect 75556 100528 75596 100568
rect 75638 100528 75678 100568
rect 75720 100528 75760 100568
rect 74152 99772 74192 99812
rect 74234 99772 74274 99812
rect 74316 99772 74356 99812
rect 74398 99772 74438 99812
rect 74480 99772 74520 99812
rect 75392 99016 75432 99056
rect 75474 99016 75514 99056
rect 75556 99016 75596 99056
rect 75638 99016 75678 99056
rect 75720 99016 75760 99056
rect 74152 98260 74192 98300
rect 74234 98260 74274 98300
rect 74316 98260 74356 98300
rect 74398 98260 74438 98300
rect 74480 98260 74520 98300
rect 75392 97504 75432 97544
rect 75474 97504 75514 97544
rect 75556 97504 75596 97544
rect 75638 97504 75678 97544
rect 75720 97504 75760 97544
rect 74152 96748 74192 96788
rect 74234 96748 74274 96788
rect 74316 96748 74356 96788
rect 74398 96748 74438 96788
rect 74480 96748 74520 96788
rect 75392 95992 75432 96032
rect 75474 95992 75514 96032
rect 75556 95992 75596 96032
rect 75638 95992 75678 96032
rect 75720 95992 75760 96032
rect 74152 95236 74192 95276
rect 74234 95236 74274 95276
rect 74316 95236 74356 95276
rect 74398 95236 74438 95276
rect 74480 95236 74520 95276
rect 75392 94480 75432 94520
rect 75474 94480 75514 94520
rect 75556 94480 75596 94520
rect 75638 94480 75678 94520
rect 75720 94480 75760 94520
rect 74152 93724 74192 93764
rect 74234 93724 74274 93764
rect 74316 93724 74356 93764
rect 74398 93724 74438 93764
rect 74480 93724 74520 93764
rect 75392 92968 75432 93008
rect 75474 92968 75514 93008
rect 75556 92968 75596 93008
rect 75638 92968 75678 93008
rect 75720 92968 75760 93008
rect 74152 92212 74192 92252
rect 74234 92212 74274 92252
rect 74316 92212 74356 92252
rect 74398 92212 74438 92252
rect 74480 92212 74520 92252
rect 75392 91456 75432 91496
rect 75474 91456 75514 91496
rect 75556 91456 75596 91496
rect 75638 91456 75678 91496
rect 75720 91456 75760 91496
rect 74152 90700 74192 90740
rect 74234 90700 74274 90740
rect 74316 90700 74356 90740
rect 74398 90700 74438 90740
rect 74480 90700 74520 90740
rect 75392 89944 75432 89984
rect 75474 89944 75514 89984
rect 75556 89944 75596 89984
rect 75638 89944 75678 89984
rect 75720 89944 75760 89984
rect 74152 89188 74192 89228
rect 74234 89188 74274 89228
rect 74316 89188 74356 89228
rect 74398 89188 74438 89228
rect 74480 89188 74520 89228
rect 75392 88432 75432 88472
rect 75474 88432 75514 88472
rect 75556 88432 75596 88472
rect 75638 88432 75678 88472
rect 75720 88432 75760 88472
rect 74152 87676 74192 87716
rect 74234 87676 74274 87716
rect 74316 87676 74356 87716
rect 74398 87676 74438 87716
rect 74480 87676 74520 87716
rect 75392 86920 75432 86960
rect 75474 86920 75514 86960
rect 75556 86920 75596 86960
rect 75638 86920 75678 86960
rect 75720 86920 75760 86960
rect 74152 86164 74192 86204
rect 74234 86164 74274 86204
rect 74316 86164 74356 86204
rect 74398 86164 74438 86204
rect 74480 86164 74520 86204
rect 75392 85408 75432 85448
rect 75474 85408 75514 85448
rect 75556 85408 75596 85448
rect 75638 85408 75678 85448
rect 75720 85408 75760 85448
rect 74152 84652 74192 84692
rect 74234 84652 74274 84692
rect 74316 84652 74356 84692
rect 74398 84652 74438 84692
rect 74480 84652 74520 84692
rect 75392 83896 75432 83936
rect 75474 83896 75514 83936
rect 75556 83896 75596 83936
rect 75638 83896 75678 83936
rect 75720 83896 75760 83936
rect 74152 83140 74192 83180
rect 74234 83140 74274 83180
rect 74316 83140 74356 83180
rect 74398 83140 74438 83180
rect 74480 83140 74520 83180
rect 75392 82384 75432 82424
rect 75474 82384 75514 82424
rect 75556 82384 75596 82424
rect 75638 82384 75678 82424
rect 75720 82384 75760 82424
rect 74152 81628 74192 81668
rect 74234 81628 74274 81668
rect 74316 81628 74356 81668
rect 74398 81628 74438 81668
rect 74480 81628 74520 81668
rect 75392 80872 75432 80912
rect 75474 80872 75514 80912
rect 75556 80872 75596 80912
rect 75638 80872 75678 80912
rect 75720 80872 75760 80912
rect 74152 80116 74192 80156
rect 74234 80116 74274 80156
rect 74316 80116 74356 80156
rect 74398 80116 74438 80156
rect 74480 80116 74520 80156
rect 75392 79360 75432 79400
rect 75474 79360 75514 79400
rect 75556 79360 75596 79400
rect 75638 79360 75678 79400
rect 75720 79360 75760 79400
rect 74152 78604 74192 78644
rect 74234 78604 74274 78644
rect 74316 78604 74356 78644
rect 74398 78604 74438 78644
rect 74480 78604 74520 78644
rect 75392 77848 75432 77888
rect 75474 77848 75514 77888
rect 75556 77848 75596 77888
rect 75638 77848 75678 77888
rect 75720 77848 75760 77888
rect 74152 77092 74192 77132
rect 74234 77092 74274 77132
rect 74316 77092 74356 77132
rect 74398 77092 74438 77132
rect 74480 77092 74520 77132
rect 75392 76336 75432 76376
rect 75474 76336 75514 76376
rect 75556 76336 75596 76376
rect 75638 76336 75678 76376
rect 75720 76336 75760 76376
rect 74152 75580 74192 75620
rect 74234 75580 74274 75620
rect 74316 75580 74356 75620
rect 74398 75580 74438 75620
rect 74480 75580 74520 75620
rect 75392 74824 75432 74864
rect 75474 74824 75514 74864
rect 75556 74824 75596 74864
rect 75638 74824 75678 74864
rect 75720 74824 75760 74864
rect 74152 74068 74192 74108
rect 74234 74068 74274 74108
rect 74316 74068 74356 74108
rect 74398 74068 74438 74108
rect 74480 74068 74520 74108
rect 75392 73312 75432 73352
rect 75474 73312 75514 73352
rect 75556 73312 75596 73352
rect 75638 73312 75678 73352
rect 75720 73312 75760 73352
rect 74152 72556 74192 72596
rect 74234 72556 74274 72596
rect 74316 72556 74356 72596
rect 74398 72556 74438 72596
rect 74480 72556 74520 72596
rect 75392 71800 75432 71840
rect 75474 71800 75514 71840
rect 75556 71800 75596 71840
rect 75638 71800 75678 71840
rect 75720 71800 75760 71840
rect 90512 151936 90552 151976
rect 90594 151936 90634 151976
rect 90676 151936 90716 151976
rect 90758 151936 90798 151976
rect 90840 151936 90880 151976
rect 89272 151180 89312 151220
rect 89354 151180 89394 151220
rect 89436 151180 89476 151220
rect 89518 151180 89558 151220
rect 89600 151180 89640 151220
rect 90512 150424 90552 150464
rect 90594 150424 90634 150464
rect 90676 150424 90716 150464
rect 90758 150424 90798 150464
rect 90840 150424 90880 150464
rect 89272 149668 89312 149708
rect 89354 149668 89394 149708
rect 89436 149668 89476 149708
rect 89518 149668 89558 149708
rect 89600 149668 89640 149708
rect 90512 148912 90552 148952
rect 90594 148912 90634 148952
rect 90676 148912 90716 148952
rect 90758 148912 90798 148952
rect 90840 148912 90880 148952
rect 89272 148156 89312 148196
rect 89354 148156 89394 148196
rect 89436 148156 89476 148196
rect 89518 148156 89558 148196
rect 89600 148156 89640 148196
rect 90512 147400 90552 147440
rect 90594 147400 90634 147440
rect 90676 147400 90716 147440
rect 90758 147400 90798 147440
rect 90840 147400 90880 147440
rect 89272 146644 89312 146684
rect 89354 146644 89394 146684
rect 89436 146644 89476 146684
rect 89518 146644 89558 146684
rect 89600 146644 89640 146684
rect 90512 145888 90552 145928
rect 90594 145888 90634 145928
rect 90676 145888 90716 145928
rect 90758 145888 90798 145928
rect 90840 145888 90880 145928
rect 89272 145132 89312 145172
rect 89354 145132 89394 145172
rect 89436 145132 89476 145172
rect 89518 145132 89558 145172
rect 89600 145132 89640 145172
rect 90512 144376 90552 144416
rect 90594 144376 90634 144416
rect 90676 144376 90716 144416
rect 90758 144376 90798 144416
rect 90840 144376 90880 144416
rect 89272 143620 89312 143660
rect 89354 143620 89394 143660
rect 89436 143620 89476 143660
rect 89518 143620 89558 143660
rect 89600 143620 89640 143660
rect 90512 142864 90552 142904
rect 90594 142864 90634 142904
rect 90676 142864 90716 142904
rect 90758 142864 90798 142904
rect 90840 142864 90880 142904
rect 89272 142108 89312 142148
rect 89354 142108 89394 142148
rect 89436 142108 89476 142148
rect 89518 142108 89558 142148
rect 89600 142108 89640 142148
rect 90512 141352 90552 141392
rect 90594 141352 90634 141392
rect 90676 141352 90716 141392
rect 90758 141352 90798 141392
rect 90840 141352 90880 141392
rect 89272 140596 89312 140636
rect 89354 140596 89394 140636
rect 89436 140596 89476 140636
rect 89518 140596 89558 140636
rect 89600 140596 89640 140636
rect 90512 139840 90552 139880
rect 90594 139840 90634 139880
rect 90676 139840 90716 139880
rect 90758 139840 90798 139880
rect 90840 139840 90880 139880
rect 89272 139084 89312 139124
rect 89354 139084 89394 139124
rect 89436 139084 89476 139124
rect 89518 139084 89558 139124
rect 89600 139084 89640 139124
rect 90512 138328 90552 138368
rect 90594 138328 90634 138368
rect 90676 138328 90716 138368
rect 90758 138328 90798 138368
rect 90840 138328 90880 138368
rect 89272 137572 89312 137612
rect 89354 137572 89394 137612
rect 89436 137572 89476 137612
rect 89518 137572 89558 137612
rect 89600 137572 89640 137612
rect 90512 136816 90552 136856
rect 90594 136816 90634 136856
rect 90676 136816 90716 136856
rect 90758 136816 90798 136856
rect 90840 136816 90880 136856
rect 89272 136060 89312 136100
rect 89354 136060 89394 136100
rect 89436 136060 89476 136100
rect 89518 136060 89558 136100
rect 89600 136060 89640 136100
rect 90512 135304 90552 135344
rect 90594 135304 90634 135344
rect 90676 135304 90716 135344
rect 90758 135304 90798 135344
rect 90840 135304 90880 135344
rect 89272 134548 89312 134588
rect 89354 134548 89394 134588
rect 89436 134548 89476 134588
rect 89518 134548 89558 134588
rect 89600 134548 89640 134588
rect 90512 133792 90552 133832
rect 90594 133792 90634 133832
rect 90676 133792 90716 133832
rect 90758 133792 90798 133832
rect 90840 133792 90880 133832
rect 89272 133036 89312 133076
rect 89354 133036 89394 133076
rect 89436 133036 89476 133076
rect 89518 133036 89558 133076
rect 89600 133036 89640 133076
rect 90512 132280 90552 132320
rect 90594 132280 90634 132320
rect 90676 132280 90716 132320
rect 90758 132280 90798 132320
rect 90840 132280 90880 132320
rect 89272 131524 89312 131564
rect 89354 131524 89394 131564
rect 89436 131524 89476 131564
rect 89518 131524 89558 131564
rect 89600 131524 89640 131564
rect 90512 130768 90552 130808
rect 90594 130768 90634 130808
rect 90676 130768 90716 130808
rect 90758 130768 90798 130808
rect 90840 130768 90880 130808
rect 89272 130012 89312 130052
rect 89354 130012 89394 130052
rect 89436 130012 89476 130052
rect 89518 130012 89558 130052
rect 89600 130012 89640 130052
rect 90512 129256 90552 129296
rect 90594 129256 90634 129296
rect 90676 129256 90716 129296
rect 90758 129256 90798 129296
rect 90840 129256 90880 129296
rect 89272 128500 89312 128540
rect 89354 128500 89394 128540
rect 89436 128500 89476 128540
rect 89518 128500 89558 128540
rect 89600 128500 89640 128540
rect 90512 127744 90552 127784
rect 90594 127744 90634 127784
rect 90676 127744 90716 127784
rect 90758 127744 90798 127784
rect 90840 127744 90880 127784
rect 89272 126988 89312 127028
rect 89354 126988 89394 127028
rect 89436 126988 89476 127028
rect 89518 126988 89558 127028
rect 89600 126988 89640 127028
rect 90512 126232 90552 126272
rect 90594 126232 90634 126272
rect 90676 126232 90716 126272
rect 90758 126232 90798 126272
rect 90840 126232 90880 126272
rect 89272 125476 89312 125516
rect 89354 125476 89394 125516
rect 89436 125476 89476 125516
rect 89518 125476 89558 125516
rect 89600 125476 89640 125516
rect 90512 124720 90552 124760
rect 90594 124720 90634 124760
rect 90676 124720 90716 124760
rect 90758 124720 90798 124760
rect 90840 124720 90880 124760
rect 89272 123964 89312 124004
rect 89354 123964 89394 124004
rect 89436 123964 89476 124004
rect 89518 123964 89558 124004
rect 89600 123964 89640 124004
rect 90512 123208 90552 123248
rect 90594 123208 90634 123248
rect 90676 123208 90716 123248
rect 90758 123208 90798 123248
rect 90840 123208 90880 123248
rect 89272 122452 89312 122492
rect 89354 122452 89394 122492
rect 89436 122452 89476 122492
rect 89518 122452 89558 122492
rect 89600 122452 89640 122492
rect 90512 121696 90552 121736
rect 90594 121696 90634 121736
rect 90676 121696 90716 121736
rect 90758 121696 90798 121736
rect 90840 121696 90880 121736
rect 89272 120940 89312 120980
rect 89354 120940 89394 120980
rect 89436 120940 89476 120980
rect 89518 120940 89558 120980
rect 89600 120940 89640 120980
rect 90512 120184 90552 120224
rect 90594 120184 90634 120224
rect 90676 120184 90716 120224
rect 90758 120184 90798 120224
rect 90840 120184 90880 120224
rect 89272 119428 89312 119468
rect 89354 119428 89394 119468
rect 89436 119428 89476 119468
rect 89518 119428 89558 119468
rect 89600 119428 89640 119468
rect 90512 118672 90552 118712
rect 90594 118672 90634 118712
rect 90676 118672 90716 118712
rect 90758 118672 90798 118712
rect 90840 118672 90880 118712
rect 89272 117916 89312 117956
rect 89354 117916 89394 117956
rect 89436 117916 89476 117956
rect 89518 117916 89558 117956
rect 89600 117916 89640 117956
rect 90512 117160 90552 117200
rect 90594 117160 90634 117200
rect 90676 117160 90716 117200
rect 90758 117160 90798 117200
rect 90840 117160 90880 117200
rect 89272 116404 89312 116444
rect 89354 116404 89394 116444
rect 89436 116404 89476 116444
rect 89518 116404 89558 116444
rect 89600 116404 89640 116444
rect 90512 115648 90552 115688
rect 90594 115648 90634 115688
rect 90676 115648 90716 115688
rect 90758 115648 90798 115688
rect 90840 115648 90880 115688
rect 89272 114892 89312 114932
rect 89354 114892 89394 114932
rect 89436 114892 89476 114932
rect 89518 114892 89558 114932
rect 89600 114892 89640 114932
rect 90512 114136 90552 114176
rect 90594 114136 90634 114176
rect 90676 114136 90716 114176
rect 90758 114136 90798 114176
rect 90840 114136 90880 114176
rect 89272 113380 89312 113420
rect 89354 113380 89394 113420
rect 89436 113380 89476 113420
rect 89518 113380 89558 113420
rect 89600 113380 89640 113420
rect 90512 112624 90552 112664
rect 90594 112624 90634 112664
rect 90676 112624 90716 112664
rect 90758 112624 90798 112664
rect 90840 112624 90880 112664
rect 89272 111868 89312 111908
rect 89354 111868 89394 111908
rect 89436 111868 89476 111908
rect 89518 111868 89558 111908
rect 89600 111868 89640 111908
rect 90512 111112 90552 111152
rect 90594 111112 90634 111152
rect 90676 111112 90716 111152
rect 90758 111112 90798 111152
rect 90840 111112 90880 111152
rect 89272 110356 89312 110396
rect 89354 110356 89394 110396
rect 89436 110356 89476 110396
rect 89518 110356 89558 110396
rect 89600 110356 89640 110396
rect 90512 109600 90552 109640
rect 90594 109600 90634 109640
rect 90676 109600 90716 109640
rect 90758 109600 90798 109640
rect 90840 109600 90880 109640
rect 89272 108844 89312 108884
rect 89354 108844 89394 108884
rect 89436 108844 89476 108884
rect 89518 108844 89558 108884
rect 89600 108844 89640 108884
rect 90512 108088 90552 108128
rect 90594 108088 90634 108128
rect 90676 108088 90716 108128
rect 90758 108088 90798 108128
rect 90840 108088 90880 108128
rect 89272 107332 89312 107372
rect 89354 107332 89394 107372
rect 89436 107332 89476 107372
rect 89518 107332 89558 107372
rect 89600 107332 89640 107372
rect 90512 106576 90552 106616
rect 90594 106576 90634 106616
rect 90676 106576 90716 106616
rect 90758 106576 90798 106616
rect 90840 106576 90880 106616
rect 89272 105820 89312 105860
rect 89354 105820 89394 105860
rect 89436 105820 89476 105860
rect 89518 105820 89558 105860
rect 89600 105820 89640 105860
rect 90512 105064 90552 105104
rect 90594 105064 90634 105104
rect 90676 105064 90716 105104
rect 90758 105064 90798 105104
rect 90840 105064 90880 105104
rect 89272 104308 89312 104348
rect 89354 104308 89394 104348
rect 89436 104308 89476 104348
rect 89518 104308 89558 104348
rect 89600 104308 89640 104348
rect 90512 103552 90552 103592
rect 90594 103552 90634 103592
rect 90676 103552 90716 103592
rect 90758 103552 90798 103592
rect 90840 103552 90880 103592
rect 89272 102796 89312 102836
rect 89354 102796 89394 102836
rect 89436 102796 89476 102836
rect 89518 102796 89558 102836
rect 89600 102796 89640 102836
rect 90512 102040 90552 102080
rect 90594 102040 90634 102080
rect 90676 102040 90716 102080
rect 90758 102040 90798 102080
rect 90840 102040 90880 102080
rect 89272 101284 89312 101324
rect 89354 101284 89394 101324
rect 89436 101284 89476 101324
rect 89518 101284 89558 101324
rect 89600 101284 89640 101324
rect 90512 100528 90552 100568
rect 90594 100528 90634 100568
rect 90676 100528 90716 100568
rect 90758 100528 90798 100568
rect 90840 100528 90880 100568
rect 89272 99772 89312 99812
rect 89354 99772 89394 99812
rect 89436 99772 89476 99812
rect 89518 99772 89558 99812
rect 89600 99772 89640 99812
rect 90512 99016 90552 99056
rect 90594 99016 90634 99056
rect 90676 99016 90716 99056
rect 90758 99016 90798 99056
rect 90840 99016 90880 99056
rect 89272 98260 89312 98300
rect 89354 98260 89394 98300
rect 89436 98260 89476 98300
rect 89518 98260 89558 98300
rect 89600 98260 89640 98300
rect 90512 97504 90552 97544
rect 90594 97504 90634 97544
rect 90676 97504 90716 97544
rect 90758 97504 90798 97544
rect 90840 97504 90880 97544
rect 89272 96748 89312 96788
rect 89354 96748 89394 96788
rect 89436 96748 89476 96788
rect 89518 96748 89558 96788
rect 89600 96748 89640 96788
rect 90512 95992 90552 96032
rect 90594 95992 90634 96032
rect 90676 95992 90716 96032
rect 90758 95992 90798 96032
rect 90840 95992 90880 96032
rect 89272 95236 89312 95276
rect 89354 95236 89394 95276
rect 89436 95236 89476 95276
rect 89518 95236 89558 95276
rect 89600 95236 89640 95276
rect 90512 94480 90552 94520
rect 90594 94480 90634 94520
rect 90676 94480 90716 94520
rect 90758 94480 90798 94520
rect 90840 94480 90880 94520
rect 89272 93724 89312 93764
rect 89354 93724 89394 93764
rect 89436 93724 89476 93764
rect 89518 93724 89558 93764
rect 89600 93724 89640 93764
rect 90512 92968 90552 93008
rect 90594 92968 90634 93008
rect 90676 92968 90716 93008
rect 90758 92968 90798 93008
rect 90840 92968 90880 93008
rect 89272 92212 89312 92252
rect 89354 92212 89394 92252
rect 89436 92212 89476 92252
rect 89518 92212 89558 92252
rect 89600 92212 89640 92252
rect 90512 91456 90552 91496
rect 90594 91456 90634 91496
rect 90676 91456 90716 91496
rect 90758 91456 90798 91496
rect 90840 91456 90880 91496
rect 89272 90700 89312 90740
rect 89354 90700 89394 90740
rect 89436 90700 89476 90740
rect 89518 90700 89558 90740
rect 89600 90700 89640 90740
rect 90512 89944 90552 89984
rect 90594 89944 90634 89984
rect 90676 89944 90716 89984
rect 90758 89944 90798 89984
rect 90840 89944 90880 89984
rect 89272 89188 89312 89228
rect 89354 89188 89394 89228
rect 89436 89188 89476 89228
rect 89518 89188 89558 89228
rect 89600 89188 89640 89228
rect 90512 88432 90552 88472
rect 90594 88432 90634 88472
rect 90676 88432 90716 88472
rect 90758 88432 90798 88472
rect 90840 88432 90880 88472
rect 89272 87676 89312 87716
rect 89354 87676 89394 87716
rect 89436 87676 89476 87716
rect 89518 87676 89558 87716
rect 89600 87676 89640 87716
rect 90512 86920 90552 86960
rect 90594 86920 90634 86960
rect 90676 86920 90716 86960
rect 90758 86920 90798 86960
rect 90840 86920 90880 86960
rect 89272 86164 89312 86204
rect 89354 86164 89394 86204
rect 89436 86164 89476 86204
rect 89518 86164 89558 86204
rect 89600 86164 89640 86204
rect 90512 85408 90552 85448
rect 90594 85408 90634 85448
rect 90676 85408 90716 85448
rect 90758 85408 90798 85448
rect 90840 85408 90880 85448
rect 89272 84652 89312 84692
rect 89354 84652 89394 84692
rect 89436 84652 89476 84692
rect 89518 84652 89558 84692
rect 89600 84652 89640 84692
rect 90512 83896 90552 83936
rect 90594 83896 90634 83936
rect 90676 83896 90716 83936
rect 90758 83896 90798 83936
rect 90840 83896 90880 83936
rect 89272 83140 89312 83180
rect 89354 83140 89394 83180
rect 89436 83140 89476 83180
rect 89518 83140 89558 83180
rect 89600 83140 89640 83180
rect 90512 82384 90552 82424
rect 90594 82384 90634 82424
rect 90676 82384 90716 82424
rect 90758 82384 90798 82424
rect 90840 82384 90880 82424
rect 89272 81628 89312 81668
rect 89354 81628 89394 81668
rect 89436 81628 89476 81668
rect 89518 81628 89558 81668
rect 89600 81628 89640 81668
rect 90512 80872 90552 80912
rect 90594 80872 90634 80912
rect 90676 80872 90716 80912
rect 90758 80872 90798 80912
rect 90840 80872 90880 80912
rect 89272 80116 89312 80156
rect 89354 80116 89394 80156
rect 89436 80116 89476 80156
rect 89518 80116 89558 80156
rect 89600 80116 89640 80156
rect 90512 79360 90552 79400
rect 90594 79360 90634 79400
rect 90676 79360 90716 79400
rect 90758 79360 90798 79400
rect 90840 79360 90880 79400
rect 89272 78604 89312 78644
rect 89354 78604 89394 78644
rect 89436 78604 89476 78644
rect 89518 78604 89558 78644
rect 89600 78604 89640 78644
rect 90512 77848 90552 77888
rect 90594 77848 90634 77888
rect 90676 77848 90716 77888
rect 90758 77848 90798 77888
rect 90840 77848 90880 77888
rect 89272 77092 89312 77132
rect 89354 77092 89394 77132
rect 89436 77092 89476 77132
rect 89518 77092 89558 77132
rect 89600 77092 89640 77132
rect 90512 76336 90552 76376
rect 90594 76336 90634 76376
rect 90676 76336 90716 76376
rect 90758 76336 90798 76376
rect 90840 76336 90880 76376
rect 89272 75580 89312 75620
rect 89354 75580 89394 75620
rect 89436 75580 89476 75620
rect 89518 75580 89558 75620
rect 89600 75580 89640 75620
rect 90512 74824 90552 74864
rect 90594 74824 90634 74864
rect 90676 74824 90716 74864
rect 90758 74824 90798 74864
rect 90840 74824 90880 74864
rect 89272 74068 89312 74108
rect 89354 74068 89394 74108
rect 89436 74068 89476 74108
rect 89518 74068 89558 74108
rect 89600 74068 89640 74108
rect 90512 73312 90552 73352
rect 90594 73312 90634 73352
rect 90676 73312 90716 73352
rect 90758 73312 90798 73352
rect 90840 73312 90880 73352
rect 89272 72556 89312 72596
rect 89354 72556 89394 72596
rect 89436 72556 89476 72596
rect 89518 72556 89558 72596
rect 89600 72556 89640 72596
rect 90512 71800 90552 71840
rect 90594 71800 90634 71840
rect 90676 71800 90716 71840
rect 90758 71800 90798 71840
rect 90840 71800 90880 71840
rect 135724 159412 135764 159452
rect 119692 159328 119732 159368
rect 105632 151936 105672 151976
rect 105714 151936 105754 151976
rect 105796 151936 105836 151976
rect 105878 151936 105918 151976
rect 105960 151936 106000 151976
rect 120752 151936 120792 151976
rect 120834 151936 120874 151976
rect 120916 151936 120956 151976
rect 120998 151936 121038 151976
rect 121080 151936 121120 151976
rect 135872 151936 135912 151976
rect 135954 151936 135994 151976
rect 136036 151936 136076 151976
rect 136118 151936 136158 151976
rect 136200 151936 136240 151976
rect 150992 151936 151032 151976
rect 151074 151936 151114 151976
rect 151156 151936 151196 151976
rect 151238 151936 151278 151976
rect 151320 151936 151360 151976
rect 104392 151180 104432 151220
rect 104474 151180 104514 151220
rect 104556 151180 104596 151220
rect 104638 151180 104678 151220
rect 104720 151180 104760 151220
rect 119512 151180 119552 151220
rect 119594 151180 119634 151220
rect 119676 151180 119716 151220
rect 119758 151180 119798 151220
rect 119840 151180 119880 151220
rect 134632 151180 134672 151220
rect 134714 151180 134754 151220
rect 134796 151180 134836 151220
rect 134878 151180 134918 151220
rect 134960 151180 135000 151220
rect 149752 151180 149792 151220
rect 149834 151180 149874 151220
rect 149916 151180 149956 151220
rect 149998 151180 150038 151220
rect 150080 151180 150120 151220
rect 105632 150424 105672 150464
rect 105714 150424 105754 150464
rect 105796 150424 105836 150464
rect 105878 150424 105918 150464
rect 105960 150424 106000 150464
rect 120752 150424 120792 150464
rect 120834 150424 120874 150464
rect 120916 150424 120956 150464
rect 120998 150424 121038 150464
rect 121080 150424 121120 150464
rect 135872 150424 135912 150464
rect 135954 150424 135994 150464
rect 136036 150424 136076 150464
rect 136118 150424 136158 150464
rect 136200 150424 136240 150464
rect 150992 150424 151032 150464
rect 151074 150424 151114 150464
rect 151156 150424 151196 150464
rect 151238 150424 151278 150464
rect 151320 150424 151360 150464
rect 104392 149668 104432 149708
rect 104474 149668 104514 149708
rect 104556 149668 104596 149708
rect 104638 149668 104678 149708
rect 104720 149668 104760 149708
rect 119512 149668 119552 149708
rect 119594 149668 119634 149708
rect 119676 149668 119716 149708
rect 119758 149668 119798 149708
rect 119840 149668 119880 149708
rect 134632 149668 134672 149708
rect 134714 149668 134754 149708
rect 134796 149668 134836 149708
rect 134878 149668 134918 149708
rect 134960 149668 135000 149708
rect 149752 149668 149792 149708
rect 149834 149668 149874 149708
rect 149916 149668 149956 149708
rect 149998 149668 150038 149708
rect 150080 149668 150120 149708
rect 105632 148912 105672 148952
rect 105714 148912 105754 148952
rect 105796 148912 105836 148952
rect 105878 148912 105918 148952
rect 105960 148912 106000 148952
rect 120752 148912 120792 148952
rect 120834 148912 120874 148952
rect 120916 148912 120956 148952
rect 120998 148912 121038 148952
rect 121080 148912 121120 148952
rect 135872 148912 135912 148952
rect 135954 148912 135994 148952
rect 136036 148912 136076 148952
rect 136118 148912 136158 148952
rect 136200 148912 136240 148952
rect 150992 148912 151032 148952
rect 151074 148912 151114 148952
rect 151156 148912 151196 148952
rect 151238 148912 151278 148952
rect 151320 148912 151360 148952
rect 104392 148156 104432 148196
rect 104474 148156 104514 148196
rect 104556 148156 104596 148196
rect 104638 148156 104678 148196
rect 104720 148156 104760 148196
rect 119512 148156 119552 148196
rect 119594 148156 119634 148196
rect 119676 148156 119716 148196
rect 119758 148156 119798 148196
rect 119840 148156 119880 148196
rect 134632 148156 134672 148196
rect 134714 148156 134754 148196
rect 134796 148156 134836 148196
rect 134878 148156 134918 148196
rect 134960 148156 135000 148196
rect 149752 148156 149792 148196
rect 149834 148156 149874 148196
rect 149916 148156 149956 148196
rect 149998 148156 150038 148196
rect 150080 148156 150120 148196
rect 105632 147400 105672 147440
rect 105714 147400 105754 147440
rect 105796 147400 105836 147440
rect 105878 147400 105918 147440
rect 105960 147400 106000 147440
rect 120752 147400 120792 147440
rect 120834 147400 120874 147440
rect 120916 147400 120956 147440
rect 120998 147400 121038 147440
rect 121080 147400 121120 147440
rect 135872 147400 135912 147440
rect 135954 147400 135994 147440
rect 136036 147400 136076 147440
rect 136118 147400 136158 147440
rect 136200 147400 136240 147440
rect 150992 147400 151032 147440
rect 151074 147400 151114 147440
rect 151156 147400 151196 147440
rect 151238 147400 151278 147440
rect 151320 147400 151360 147440
rect 104392 146644 104432 146684
rect 104474 146644 104514 146684
rect 104556 146644 104596 146684
rect 104638 146644 104678 146684
rect 104720 146644 104760 146684
rect 119512 146644 119552 146684
rect 119594 146644 119634 146684
rect 119676 146644 119716 146684
rect 119758 146644 119798 146684
rect 119840 146644 119880 146684
rect 134632 146644 134672 146684
rect 134714 146644 134754 146684
rect 134796 146644 134836 146684
rect 134878 146644 134918 146684
rect 134960 146644 135000 146684
rect 149752 146644 149792 146684
rect 149834 146644 149874 146684
rect 149916 146644 149956 146684
rect 149998 146644 150038 146684
rect 150080 146644 150120 146684
rect 105632 145888 105672 145928
rect 105714 145888 105754 145928
rect 105796 145888 105836 145928
rect 105878 145888 105918 145928
rect 105960 145888 106000 145928
rect 120752 145888 120792 145928
rect 120834 145888 120874 145928
rect 120916 145888 120956 145928
rect 120998 145888 121038 145928
rect 121080 145888 121120 145928
rect 135872 145888 135912 145928
rect 135954 145888 135994 145928
rect 136036 145888 136076 145928
rect 136118 145888 136158 145928
rect 136200 145888 136240 145928
rect 150992 145888 151032 145928
rect 151074 145888 151114 145928
rect 151156 145888 151196 145928
rect 151238 145888 151278 145928
rect 151320 145888 151360 145928
rect 104392 145132 104432 145172
rect 104474 145132 104514 145172
rect 104556 145132 104596 145172
rect 104638 145132 104678 145172
rect 104720 145132 104760 145172
rect 119512 145132 119552 145172
rect 119594 145132 119634 145172
rect 119676 145132 119716 145172
rect 119758 145132 119798 145172
rect 119840 145132 119880 145172
rect 134632 145132 134672 145172
rect 134714 145132 134754 145172
rect 134796 145132 134836 145172
rect 134878 145132 134918 145172
rect 134960 145132 135000 145172
rect 149752 145132 149792 145172
rect 149834 145132 149874 145172
rect 149916 145132 149956 145172
rect 149998 145132 150038 145172
rect 150080 145132 150120 145172
rect 105632 144376 105672 144416
rect 105714 144376 105754 144416
rect 105796 144376 105836 144416
rect 105878 144376 105918 144416
rect 105960 144376 106000 144416
rect 120752 144376 120792 144416
rect 120834 144376 120874 144416
rect 120916 144376 120956 144416
rect 120998 144376 121038 144416
rect 121080 144376 121120 144416
rect 135872 144376 135912 144416
rect 135954 144376 135994 144416
rect 136036 144376 136076 144416
rect 136118 144376 136158 144416
rect 136200 144376 136240 144416
rect 150992 144376 151032 144416
rect 151074 144376 151114 144416
rect 151156 144376 151196 144416
rect 151238 144376 151278 144416
rect 151320 144376 151360 144416
rect 104392 143620 104432 143660
rect 104474 143620 104514 143660
rect 104556 143620 104596 143660
rect 104638 143620 104678 143660
rect 104720 143620 104760 143660
rect 119512 143620 119552 143660
rect 119594 143620 119634 143660
rect 119676 143620 119716 143660
rect 119758 143620 119798 143660
rect 119840 143620 119880 143660
rect 134632 143620 134672 143660
rect 134714 143620 134754 143660
rect 134796 143620 134836 143660
rect 134878 143620 134918 143660
rect 134960 143620 135000 143660
rect 149752 143620 149792 143660
rect 149834 143620 149874 143660
rect 149916 143620 149956 143660
rect 149998 143620 150038 143660
rect 150080 143620 150120 143660
rect 105632 142864 105672 142904
rect 105714 142864 105754 142904
rect 105796 142864 105836 142904
rect 105878 142864 105918 142904
rect 105960 142864 106000 142904
rect 120752 142864 120792 142904
rect 120834 142864 120874 142904
rect 120916 142864 120956 142904
rect 120998 142864 121038 142904
rect 121080 142864 121120 142904
rect 135872 142864 135912 142904
rect 135954 142864 135994 142904
rect 136036 142864 136076 142904
rect 136118 142864 136158 142904
rect 136200 142864 136240 142904
rect 150992 142864 151032 142904
rect 151074 142864 151114 142904
rect 151156 142864 151196 142904
rect 151238 142864 151278 142904
rect 151320 142864 151360 142904
rect 104392 142108 104432 142148
rect 104474 142108 104514 142148
rect 104556 142108 104596 142148
rect 104638 142108 104678 142148
rect 104720 142108 104760 142148
rect 119512 142108 119552 142148
rect 119594 142108 119634 142148
rect 119676 142108 119716 142148
rect 119758 142108 119798 142148
rect 119840 142108 119880 142148
rect 134632 142108 134672 142148
rect 134714 142108 134754 142148
rect 134796 142108 134836 142148
rect 134878 142108 134918 142148
rect 134960 142108 135000 142148
rect 149752 142108 149792 142148
rect 149834 142108 149874 142148
rect 149916 142108 149956 142148
rect 149998 142108 150038 142148
rect 150080 142108 150120 142148
rect 105632 141352 105672 141392
rect 105714 141352 105754 141392
rect 105796 141352 105836 141392
rect 105878 141352 105918 141392
rect 105960 141352 106000 141392
rect 120752 141352 120792 141392
rect 120834 141352 120874 141392
rect 120916 141352 120956 141392
rect 120998 141352 121038 141392
rect 121080 141352 121120 141392
rect 135872 141352 135912 141392
rect 135954 141352 135994 141392
rect 136036 141352 136076 141392
rect 136118 141352 136158 141392
rect 136200 141352 136240 141392
rect 150992 141352 151032 141392
rect 151074 141352 151114 141392
rect 151156 141352 151196 141392
rect 151238 141352 151278 141392
rect 151320 141352 151360 141392
rect 104392 140596 104432 140636
rect 104474 140596 104514 140636
rect 104556 140596 104596 140636
rect 104638 140596 104678 140636
rect 104720 140596 104760 140636
rect 119512 140596 119552 140636
rect 119594 140596 119634 140636
rect 119676 140596 119716 140636
rect 119758 140596 119798 140636
rect 119840 140596 119880 140636
rect 134632 140596 134672 140636
rect 134714 140596 134754 140636
rect 134796 140596 134836 140636
rect 134878 140596 134918 140636
rect 134960 140596 135000 140636
rect 149752 140596 149792 140636
rect 149834 140596 149874 140636
rect 149916 140596 149956 140636
rect 149998 140596 150038 140636
rect 150080 140596 150120 140636
rect 105632 139840 105672 139880
rect 105714 139840 105754 139880
rect 105796 139840 105836 139880
rect 105878 139840 105918 139880
rect 105960 139840 106000 139880
rect 120752 139840 120792 139880
rect 120834 139840 120874 139880
rect 120916 139840 120956 139880
rect 120998 139840 121038 139880
rect 121080 139840 121120 139880
rect 135872 139840 135912 139880
rect 135954 139840 135994 139880
rect 136036 139840 136076 139880
rect 136118 139840 136158 139880
rect 136200 139840 136240 139880
rect 150992 139840 151032 139880
rect 151074 139840 151114 139880
rect 151156 139840 151196 139880
rect 151238 139840 151278 139880
rect 151320 139840 151360 139880
rect 104392 139084 104432 139124
rect 104474 139084 104514 139124
rect 104556 139084 104596 139124
rect 104638 139084 104678 139124
rect 104720 139084 104760 139124
rect 119512 139084 119552 139124
rect 119594 139084 119634 139124
rect 119676 139084 119716 139124
rect 119758 139084 119798 139124
rect 119840 139084 119880 139124
rect 134632 139084 134672 139124
rect 134714 139084 134754 139124
rect 134796 139084 134836 139124
rect 134878 139084 134918 139124
rect 134960 139084 135000 139124
rect 149752 139084 149792 139124
rect 149834 139084 149874 139124
rect 149916 139084 149956 139124
rect 149998 139084 150038 139124
rect 150080 139084 150120 139124
rect 105632 138328 105672 138368
rect 105714 138328 105754 138368
rect 105796 138328 105836 138368
rect 105878 138328 105918 138368
rect 105960 138328 106000 138368
rect 120752 138328 120792 138368
rect 120834 138328 120874 138368
rect 120916 138328 120956 138368
rect 120998 138328 121038 138368
rect 121080 138328 121120 138368
rect 135872 138328 135912 138368
rect 135954 138328 135994 138368
rect 136036 138328 136076 138368
rect 136118 138328 136158 138368
rect 136200 138328 136240 138368
rect 150992 138328 151032 138368
rect 151074 138328 151114 138368
rect 151156 138328 151196 138368
rect 151238 138328 151278 138368
rect 151320 138328 151360 138368
rect 104392 137572 104432 137612
rect 104474 137572 104514 137612
rect 104556 137572 104596 137612
rect 104638 137572 104678 137612
rect 104720 137572 104760 137612
rect 119512 137572 119552 137612
rect 119594 137572 119634 137612
rect 119676 137572 119716 137612
rect 119758 137572 119798 137612
rect 119840 137572 119880 137612
rect 134632 137572 134672 137612
rect 134714 137572 134754 137612
rect 134796 137572 134836 137612
rect 134878 137572 134918 137612
rect 134960 137572 135000 137612
rect 149752 137572 149792 137612
rect 149834 137572 149874 137612
rect 149916 137572 149956 137612
rect 149998 137572 150038 137612
rect 150080 137572 150120 137612
rect 105632 136816 105672 136856
rect 105714 136816 105754 136856
rect 105796 136816 105836 136856
rect 105878 136816 105918 136856
rect 105960 136816 106000 136856
rect 120752 136816 120792 136856
rect 120834 136816 120874 136856
rect 120916 136816 120956 136856
rect 120998 136816 121038 136856
rect 121080 136816 121120 136856
rect 135872 136816 135912 136856
rect 135954 136816 135994 136856
rect 136036 136816 136076 136856
rect 136118 136816 136158 136856
rect 136200 136816 136240 136856
rect 150992 136816 151032 136856
rect 151074 136816 151114 136856
rect 151156 136816 151196 136856
rect 151238 136816 151278 136856
rect 151320 136816 151360 136856
rect 104392 136060 104432 136100
rect 104474 136060 104514 136100
rect 104556 136060 104596 136100
rect 104638 136060 104678 136100
rect 104720 136060 104760 136100
rect 119512 136060 119552 136100
rect 119594 136060 119634 136100
rect 119676 136060 119716 136100
rect 119758 136060 119798 136100
rect 119840 136060 119880 136100
rect 134632 136060 134672 136100
rect 134714 136060 134754 136100
rect 134796 136060 134836 136100
rect 134878 136060 134918 136100
rect 134960 136060 135000 136100
rect 149752 136060 149792 136100
rect 149834 136060 149874 136100
rect 149916 136060 149956 136100
rect 149998 136060 150038 136100
rect 150080 136060 150120 136100
rect 105632 135304 105672 135344
rect 105714 135304 105754 135344
rect 105796 135304 105836 135344
rect 105878 135304 105918 135344
rect 105960 135304 106000 135344
rect 120752 135304 120792 135344
rect 120834 135304 120874 135344
rect 120916 135304 120956 135344
rect 120998 135304 121038 135344
rect 121080 135304 121120 135344
rect 135872 135304 135912 135344
rect 135954 135304 135994 135344
rect 136036 135304 136076 135344
rect 136118 135304 136158 135344
rect 136200 135304 136240 135344
rect 150992 135304 151032 135344
rect 151074 135304 151114 135344
rect 151156 135304 151196 135344
rect 151238 135304 151278 135344
rect 151320 135304 151360 135344
rect 104392 134548 104432 134588
rect 104474 134548 104514 134588
rect 104556 134548 104596 134588
rect 104638 134548 104678 134588
rect 104720 134548 104760 134588
rect 119512 134548 119552 134588
rect 119594 134548 119634 134588
rect 119676 134548 119716 134588
rect 119758 134548 119798 134588
rect 119840 134548 119880 134588
rect 134632 134548 134672 134588
rect 134714 134548 134754 134588
rect 134796 134548 134836 134588
rect 134878 134548 134918 134588
rect 134960 134548 135000 134588
rect 149752 134548 149792 134588
rect 149834 134548 149874 134588
rect 149916 134548 149956 134588
rect 149998 134548 150038 134588
rect 150080 134548 150120 134588
rect 105632 133792 105672 133832
rect 105714 133792 105754 133832
rect 105796 133792 105836 133832
rect 105878 133792 105918 133832
rect 105960 133792 106000 133832
rect 120752 133792 120792 133832
rect 120834 133792 120874 133832
rect 120916 133792 120956 133832
rect 120998 133792 121038 133832
rect 121080 133792 121120 133832
rect 135872 133792 135912 133832
rect 135954 133792 135994 133832
rect 136036 133792 136076 133832
rect 136118 133792 136158 133832
rect 136200 133792 136240 133832
rect 150992 133792 151032 133832
rect 151074 133792 151114 133832
rect 151156 133792 151196 133832
rect 151238 133792 151278 133832
rect 151320 133792 151360 133832
rect 104392 133036 104432 133076
rect 104474 133036 104514 133076
rect 104556 133036 104596 133076
rect 104638 133036 104678 133076
rect 104720 133036 104760 133076
rect 119512 133036 119552 133076
rect 119594 133036 119634 133076
rect 119676 133036 119716 133076
rect 119758 133036 119798 133076
rect 119840 133036 119880 133076
rect 134632 133036 134672 133076
rect 134714 133036 134754 133076
rect 134796 133036 134836 133076
rect 134878 133036 134918 133076
rect 134960 133036 135000 133076
rect 149752 133036 149792 133076
rect 149834 133036 149874 133076
rect 149916 133036 149956 133076
rect 149998 133036 150038 133076
rect 150080 133036 150120 133076
rect 105632 132280 105672 132320
rect 105714 132280 105754 132320
rect 105796 132280 105836 132320
rect 105878 132280 105918 132320
rect 105960 132280 106000 132320
rect 120752 132280 120792 132320
rect 120834 132280 120874 132320
rect 120916 132280 120956 132320
rect 120998 132280 121038 132320
rect 121080 132280 121120 132320
rect 135872 132280 135912 132320
rect 135954 132280 135994 132320
rect 136036 132280 136076 132320
rect 136118 132280 136158 132320
rect 136200 132280 136240 132320
rect 150992 132280 151032 132320
rect 151074 132280 151114 132320
rect 151156 132280 151196 132320
rect 151238 132280 151278 132320
rect 151320 132280 151360 132320
rect 104392 131524 104432 131564
rect 104474 131524 104514 131564
rect 104556 131524 104596 131564
rect 104638 131524 104678 131564
rect 104720 131524 104760 131564
rect 119512 131524 119552 131564
rect 119594 131524 119634 131564
rect 119676 131524 119716 131564
rect 119758 131524 119798 131564
rect 119840 131524 119880 131564
rect 134632 131524 134672 131564
rect 134714 131524 134754 131564
rect 134796 131524 134836 131564
rect 134878 131524 134918 131564
rect 134960 131524 135000 131564
rect 149752 131524 149792 131564
rect 149834 131524 149874 131564
rect 149916 131524 149956 131564
rect 149998 131524 150038 131564
rect 150080 131524 150120 131564
rect 105632 130768 105672 130808
rect 105714 130768 105754 130808
rect 105796 130768 105836 130808
rect 105878 130768 105918 130808
rect 105960 130768 106000 130808
rect 120752 130768 120792 130808
rect 120834 130768 120874 130808
rect 120916 130768 120956 130808
rect 120998 130768 121038 130808
rect 121080 130768 121120 130808
rect 135872 130768 135912 130808
rect 135954 130768 135994 130808
rect 136036 130768 136076 130808
rect 136118 130768 136158 130808
rect 136200 130768 136240 130808
rect 150992 130768 151032 130808
rect 151074 130768 151114 130808
rect 151156 130768 151196 130808
rect 151238 130768 151278 130808
rect 151320 130768 151360 130808
rect 104392 130012 104432 130052
rect 104474 130012 104514 130052
rect 104556 130012 104596 130052
rect 104638 130012 104678 130052
rect 104720 130012 104760 130052
rect 119512 130012 119552 130052
rect 119594 130012 119634 130052
rect 119676 130012 119716 130052
rect 119758 130012 119798 130052
rect 119840 130012 119880 130052
rect 134632 130012 134672 130052
rect 134714 130012 134754 130052
rect 134796 130012 134836 130052
rect 134878 130012 134918 130052
rect 134960 130012 135000 130052
rect 149752 130012 149792 130052
rect 149834 130012 149874 130052
rect 149916 130012 149956 130052
rect 149998 130012 150038 130052
rect 150080 130012 150120 130052
rect 105632 129256 105672 129296
rect 105714 129256 105754 129296
rect 105796 129256 105836 129296
rect 105878 129256 105918 129296
rect 105960 129256 106000 129296
rect 120752 129256 120792 129296
rect 120834 129256 120874 129296
rect 120916 129256 120956 129296
rect 120998 129256 121038 129296
rect 121080 129256 121120 129296
rect 135872 129256 135912 129296
rect 135954 129256 135994 129296
rect 136036 129256 136076 129296
rect 136118 129256 136158 129296
rect 136200 129256 136240 129296
rect 150992 129256 151032 129296
rect 151074 129256 151114 129296
rect 151156 129256 151196 129296
rect 151238 129256 151278 129296
rect 151320 129256 151360 129296
rect 104392 128500 104432 128540
rect 104474 128500 104514 128540
rect 104556 128500 104596 128540
rect 104638 128500 104678 128540
rect 104720 128500 104760 128540
rect 119512 128500 119552 128540
rect 119594 128500 119634 128540
rect 119676 128500 119716 128540
rect 119758 128500 119798 128540
rect 119840 128500 119880 128540
rect 134632 128500 134672 128540
rect 134714 128500 134754 128540
rect 134796 128500 134836 128540
rect 134878 128500 134918 128540
rect 134960 128500 135000 128540
rect 149752 128500 149792 128540
rect 149834 128500 149874 128540
rect 149916 128500 149956 128540
rect 149998 128500 150038 128540
rect 150080 128500 150120 128540
rect 105632 127744 105672 127784
rect 105714 127744 105754 127784
rect 105796 127744 105836 127784
rect 105878 127744 105918 127784
rect 105960 127744 106000 127784
rect 120752 127744 120792 127784
rect 120834 127744 120874 127784
rect 120916 127744 120956 127784
rect 120998 127744 121038 127784
rect 121080 127744 121120 127784
rect 135872 127744 135912 127784
rect 135954 127744 135994 127784
rect 136036 127744 136076 127784
rect 136118 127744 136158 127784
rect 136200 127744 136240 127784
rect 150992 127744 151032 127784
rect 151074 127744 151114 127784
rect 151156 127744 151196 127784
rect 151238 127744 151278 127784
rect 151320 127744 151360 127784
rect 104392 126988 104432 127028
rect 104474 126988 104514 127028
rect 104556 126988 104596 127028
rect 104638 126988 104678 127028
rect 104720 126988 104760 127028
rect 119512 126988 119552 127028
rect 119594 126988 119634 127028
rect 119676 126988 119716 127028
rect 119758 126988 119798 127028
rect 119840 126988 119880 127028
rect 134632 126988 134672 127028
rect 134714 126988 134754 127028
rect 134796 126988 134836 127028
rect 134878 126988 134918 127028
rect 134960 126988 135000 127028
rect 149752 126988 149792 127028
rect 149834 126988 149874 127028
rect 149916 126988 149956 127028
rect 149998 126988 150038 127028
rect 150080 126988 150120 127028
rect 105632 126232 105672 126272
rect 105714 126232 105754 126272
rect 105796 126232 105836 126272
rect 105878 126232 105918 126272
rect 105960 126232 106000 126272
rect 120752 126232 120792 126272
rect 120834 126232 120874 126272
rect 120916 126232 120956 126272
rect 120998 126232 121038 126272
rect 121080 126232 121120 126272
rect 135872 126232 135912 126272
rect 135954 126232 135994 126272
rect 136036 126232 136076 126272
rect 136118 126232 136158 126272
rect 136200 126232 136240 126272
rect 150992 126232 151032 126272
rect 151074 126232 151114 126272
rect 151156 126232 151196 126272
rect 151238 126232 151278 126272
rect 151320 126232 151360 126272
rect 104392 125476 104432 125516
rect 104474 125476 104514 125516
rect 104556 125476 104596 125516
rect 104638 125476 104678 125516
rect 104720 125476 104760 125516
rect 119512 125476 119552 125516
rect 119594 125476 119634 125516
rect 119676 125476 119716 125516
rect 119758 125476 119798 125516
rect 119840 125476 119880 125516
rect 134632 125476 134672 125516
rect 134714 125476 134754 125516
rect 134796 125476 134836 125516
rect 134878 125476 134918 125516
rect 134960 125476 135000 125516
rect 149752 125476 149792 125516
rect 149834 125476 149874 125516
rect 149916 125476 149956 125516
rect 149998 125476 150038 125516
rect 150080 125476 150120 125516
rect 105632 124720 105672 124760
rect 105714 124720 105754 124760
rect 105796 124720 105836 124760
rect 105878 124720 105918 124760
rect 105960 124720 106000 124760
rect 120752 124720 120792 124760
rect 120834 124720 120874 124760
rect 120916 124720 120956 124760
rect 120998 124720 121038 124760
rect 121080 124720 121120 124760
rect 135872 124720 135912 124760
rect 135954 124720 135994 124760
rect 136036 124720 136076 124760
rect 136118 124720 136158 124760
rect 136200 124720 136240 124760
rect 150992 124720 151032 124760
rect 151074 124720 151114 124760
rect 151156 124720 151196 124760
rect 151238 124720 151278 124760
rect 151320 124720 151360 124760
rect 104392 123964 104432 124004
rect 104474 123964 104514 124004
rect 104556 123964 104596 124004
rect 104638 123964 104678 124004
rect 104720 123964 104760 124004
rect 119512 123964 119552 124004
rect 119594 123964 119634 124004
rect 119676 123964 119716 124004
rect 119758 123964 119798 124004
rect 119840 123964 119880 124004
rect 134632 123964 134672 124004
rect 134714 123964 134754 124004
rect 134796 123964 134836 124004
rect 134878 123964 134918 124004
rect 134960 123964 135000 124004
rect 149752 123964 149792 124004
rect 149834 123964 149874 124004
rect 149916 123964 149956 124004
rect 149998 123964 150038 124004
rect 150080 123964 150120 124004
rect 105632 123208 105672 123248
rect 105714 123208 105754 123248
rect 105796 123208 105836 123248
rect 105878 123208 105918 123248
rect 105960 123208 106000 123248
rect 120752 123208 120792 123248
rect 120834 123208 120874 123248
rect 120916 123208 120956 123248
rect 120998 123208 121038 123248
rect 121080 123208 121120 123248
rect 135872 123208 135912 123248
rect 135954 123208 135994 123248
rect 136036 123208 136076 123248
rect 136118 123208 136158 123248
rect 136200 123208 136240 123248
rect 150992 123208 151032 123248
rect 151074 123208 151114 123248
rect 151156 123208 151196 123248
rect 151238 123208 151278 123248
rect 151320 123208 151360 123248
rect 104392 122452 104432 122492
rect 104474 122452 104514 122492
rect 104556 122452 104596 122492
rect 104638 122452 104678 122492
rect 104720 122452 104760 122492
rect 119512 122452 119552 122492
rect 119594 122452 119634 122492
rect 119676 122452 119716 122492
rect 119758 122452 119798 122492
rect 119840 122452 119880 122492
rect 134632 122452 134672 122492
rect 134714 122452 134754 122492
rect 134796 122452 134836 122492
rect 134878 122452 134918 122492
rect 134960 122452 135000 122492
rect 149752 122452 149792 122492
rect 149834 122452 149874 122492
rect 149916 122452 149956 122492
rect 149998 122452 150038 122492
rect 150080 122452 150120 122492
rect 105632 121696 105672 121736
rect 105714 121696 105754 121736
rect 105796 121696 105836 121736
rect 105878 121696 105918 121736
rect 105960 121696 106000 121736
rect 120752 121696 120792 121736
rect 120834 121696 120874 121736
rect 120916 121696 120956 121736
rect 120998 121696 121038 121736
rect 121080 121696 121120 121736
rect 135872 121696 135912 121736
rect 135954 121696 135994 121736
rect 136036 121696 136076 121736
rect 136118 121696 136158 121736
rect 136200 121696 136240 121736
rect 150992 121696 151032 121736
rect 151074 121696 151114 121736
rect 151156 121696 151196 121736
rect 151238 121696 151278 121736
rect 151320 121696 151360 121736
rect 104392 120940 104432 120980
rect 104474 120940 104514 120980
rect 104556 120940 104596 120980
rect 104638 120940 104678 120980
rect 104720 120940 104760 120980
rect 119512 120940 119552 120980
rect 119594 120940 119634 120980
rect 119676 120940 119716 120980
rect 119758 120940 119798 120980
rect 119840 120940 119880 120980
rect 134632 120940 134672 120980
rect 134714 120940 134754 120980
rect 134796 120940 134836 120980
rect 134878 120940 134918 120980
rect 134960 120940 135000 120980
rect 149752 120940 149792 120980
rect 149834 120940 149874 120980
rect 149916 120940 149956 120980
rect 149998 120940 150038 120980
rect 150080 120940 150120 120980
rect 105632 120184 105672 120224
rect 105714 120184 105754 120224
rect 105796 120184 105836 120224
rect 105878 120184 105918 120224
rect 105960 120184 106000 120224
rect 120752 120184 120792 120224
rect 120834 120184 120874 120224
rect 120916 120184 120956 120224
rect 120998 120184 121038 120224
rect 121080 120184 121120 120224
rect 135872 120184 135912 120224
rect 135954 120184 135994 120224
rect 136036 120184 136076 120224
rect 136118 120184 136158 120224
rect 136200 120184 136240 120224
rect 150992 120184 151032 120224
rect 151074 120184 151114 120224
rect 151156 120184 151196 120224
rect 151238 120184 151278 120224
rect 151320 120184 151360 120224
rect 104392 119428 104432 119468
rect 104474 119428 104514 119468
rect 104556 119428 104596 119468
rect 104638 119428 104678 119468
rect 104720 119428 104760 119468
rect 119512 119428 119552 119468
rect 119594 119428 119634 119468
rect 119676 119428 119716 119468
rect 119758 119428 119798 119468
rect 119840 119428 119880 119468
rect 134632 119428 134672 119468
rect 134714 119428 134754 119468
rect 134796 119428 134836 119468
rect 134878 119428 134918 119468
rect 134960 119428 135000 119468
rect 149752 119428 149792 119468
rect 149834 119428 149874 119468
rect 149916 119428 149956 119468
rect 149998 119428 150038 119468
rect 150080 119428 150120 119468
rect 105632 118672 105672 118712
rect 105714 118672 105754 118712
rect 105796 118672 105836 118712
rect 105878 118672 105918 118712
rect 105960 118672 106000 118712
rect 120752 118672 120792 118712
rect 120834 118672 120874 118712
rect 120916 118672 120956 118712
rect 120998 118672 121038 118712
rect 121080 118672 121120 118712
rect 135872 118672 135912 118712
rect 135954 118672 135994 118712
rect 136036 118672 136076 118712
rect 136118 118672 136158 118712
rect 136200 118672 136240 118712
rect 150992 118672 151032 118712
rect 151074 118672 151114 118712
rect 151156 118672 151196 118712
rect 151238 118672 151278 118712
rect 151320 118672 151360 118712
rect 104392 117916 104432 117956
rect 104474 117916 104514 117956
rect 104556 117916 104596 117956
rect 104638 117916 104678 117956
rect 104720 117916 104760 117956
rect 119512 117916 119552 117956
rect 119594 117916 119634 117956
rect 119676 117916 119716 117956
rect 119758 117916 119798 117956
rect 119840 117916 119880 117956
rect 134632 117916 134672 117956
rect 134714 117916 134754 117956
rect 134796 117916 134836 117956
rect 134878 117916 134918 117956
rect 134960 117916 135000 117956
rect 149752 117916 149792 117956
rect 149834 117916 149874 117956
rect 149916 117916 149956 117956
rect 149998 117916 150038 117956
rect 150080 117916 150120 117956
rect 105632 117160 105672 117200
rect 105714 117160 105754 117200
rect 105796 117160 105836 117200
rect 105878 117160 105918 117200
rect 105960 117160 106000 117200
rect 120752 117160 120792 117200
rect 120834 117160 120874 117200
rect 120916 117160 120956 117200
rect 120998 117160 121038 117200
rect 121080 117160 121120 117200
rect 135872 117160 135912 117200
rect 135954 117160 135994 117200
rect 136036 117160 136076 117200
rect 136118 117160 136158 117200
rect 136200 117160 136240 117200
rect 150992 117160 151032 117200
rect 151074 117160 151114 117200
rect 151156 117160 151196 117200
rect 151238 117160 151278 117200
rect 151320 117160 151360 117200
rect 104392 116404 104432 116444
rect 104474 116404 104514 116444
rect 104556 116404 104596 116444
rect 104638 116404 104678 116444
rect 104720 116404 104760 116444
rect 119512 116404 119552 116444
rect 119594 116404 119634 116444
rect 119676 116404 119716 116444
rect 119758 116404 119798 116444
rect 119840 116404 119880 116444
rect 134632 116404 134672 116444
rect 134714 116404 134754 116444
rect 134796 116404 134836 116444
rect 134878 116404 134918 116444
rect 134960 116404 135000 116444
rect 149752 116404 149792 116444
rect 149834 116404 149874 116444
rect 149916 116404 149956 116444
rect 149998 116404 150038 116444
rect 150080 116404 150120 116444
rect 105632 115648 105672 115688
rect 105714 115648 105754 115688
rect 105796 115648 105836 115688
rect 105878 115648 105918 115688
rect 105960 115648 106000 115688
rect 120752 115648 120792 115688
rect 120834 115648 120874 115688
rect 120916 115648 120956 115688
rect 120998 115648 121038 115688
rect 121080 115648 121120 115688
rect 135872 115648 135912 115688
rect 135954 115648 135994 115688
rect 136036 115648 136076 115688
rect 136118 115648 136158 115688
rect 136200 115648 136240 115688
rect 150992 115648 151032 115688
rect 151074 115648 151114 115688
rect 151156 115648 151196 115688
rect 151238 115648 151278 115688
rect 151320 115648 151360 115688
rect 104392 114892 104432 114932
rect 104474 114892 104514 114932
rect 104556 114892 104596 114932
rect 104638 114892 104678 114932
rect 104720 114892 104760 114932
rect 119512 114892 119552 114932
rect 119594 114892 119634 114932
rect 119676 114892 119716 114932
rect 119758 114892 119798 114932
rect 119840 114892 119880 114932
rect 134632 114892 134672 114932
rect 134714 114892 134754 114932
rect 134796 114892 134836 114932
rect 134878 114892 134918 114932
rect 134960 114892 135000 114932
rect 149752 114892 149792 114932
rect 149834 114892 149874 114932
rect 149916 114892 149956 114932
rect 149998 114892 150038 114932
rect 150080 114892 150120 114932
rect 105632 114136 105672 114176
rect 105714 114136 105754 114176
rect 105796 114136 105836 114176
rect 105878 114136 105918 114176
rect 105960 114136 106000 114176
rect 120752 114136 120792 114176
rect 120834 114136 120874 114176
rect 120916 114136 120956 114176
rect 120998 114136 121038 114176
rect 121080 114136 121120 114176
rect 135872 114136 135912 114176
rect 135954 114136 135994 114176
rect 136036 114136 136076 114176
rect 136118 114136 136158 114176
rect 136200 114136 136240 114176
rect 150992 114136 151032 114176
rect 151074 114136 151114 114176
rect 151156 114136 151196 114176
rect 151238 114136 151278 114176
rect 151320 114136 151360 114176
rect 104392 113380 104432 113420
rect 104474 113380 104514 113420
rect 104556 113380 104596 113420
rect 104638 113380 104678 113420
rect 104720 113380 104760 113420
rect 119512 113380 119552 113420
rect 119594 113380 119634 113420
rect 119676 113380 119716 113420
rect 119758 113380 119798 113420
rect 119840 113380 119880 113420
rect 134632 113380 134672 113420
rect 134714 113380 134754 113420
rect 134796 113380 134836 113420
rect 134878 113380 134918 113420
rect 134960 113380 135000 113420
rect 149752 113380 149792 113420
rect 149834 113380 149874 113420
rect 149916 113380 149956 113420
rect 149998 113380 150038 113420
rect 150080 113380 150120 113420
rect 105632 112624 105672 112664
rect 105714 112624 105754 112664
rect 105796 112624 105836 112664
rect 105878 112624 105918 112664
rect 105960 112624 106000 112664
rect 120752 112624 120792 112664
rect 120834 112624 120874 112664
rect 120916 112624 120956 112664
rect 120998 112624 121038 112664
rect 121080 112624 121120 112664
rect 135872 112624 135912 112664
rect 135954 112624 135994 112664
rect 136036 112624 136076 112664
rect 136118 112624 136158 112664
rect 136200 112624 136240 112664
rect 150992 112624 151032 112664
rect 151074 112624 151114 112664
rect 151156 112624 151196 112664
rect 151238 112624 151278 112664
rect 151320 112624 151360 112664
rect 104392 111868 104432 111908
rect 104474 111868 104514 111908
rect 104556 111868 104596 111908
rect 104638 111868 104678 111908
rect 104720 111868 104760 111908
rect 119512 111868 119552 111908
rect 119594 111868 119634 111908
rect 119676 111868 119716 111908
rect 119758 111868 119798 111908
rect 119840 111868 119880 111908
rect 134632 111868 134672 111908
rect 134714 111868 134754 111908
rect 134796 111868 134836 111908
rect 134878 111868 134918 111908
rect 134960 111868 135000 111908
rect 149752 111868 149792 111908
rect 149834 111868 149874 111908
rect 149916 111868 149956 111908
rect 149998 111868 150038 111908
rect 150080 111868 150120 111908
rect 105632 111112 105672 111152
rect 105714 111112 105754 111152
rect 105796 111112 105836 111152
rect 105878 111112 105918 111152
rect 105960 111112 106000 111152
rect 120752 111112 120792 111152
rect 120834 111112 120874 111152
rect 120916 111112 120956 111152
rect 120998 111112 121038 111152
rect 121080 111112 121120 111152
rect 135872 111112 135912 111152
rect 135954 111112 135994 111152
rect 136036 111112 136076 111152
rect 136118 111112 136158 111152
rect 136200 111112 136240 111152
rect 150992 111112 151032 111152
rect 151074 111112 151114 111152
rect 151156 111112 151196 111152
rect 151238 111112 151278 111152
rect 151320 111112 151360 111152
rect 104392 110356 104432 110396
rect 104474 110356 104514 110396
rect 104556 110356 104596 110396
rect 104638 110356 104678 110396
rect 104720 110356 104760 110396
rect 119512 110356 119552 110396
rect 119594 110356 119634 110396
rect 119676 110356 119716 110396
rect 119758 110356 119798 110396
rect 119840 110356 119880 110396
rect 134632 110356 134672 110396
rect 134714 110356 134754 110396
rect 134796 110356 134836 110396
rect 134878 110356 134918 110396
rect 134960 110356 135000 110396
rect 149752 110356 149792 110396
rect 149834 110356 149874 110396
rect 149916 110356 149956 110396
rect 149998 110356 150038 110396
rect 150080 110356 150120 110396
rect 105632 109600 105672 109640
rect 105714 109600 105754 109640
rect 105796 109600 105836 109640
rect 105878 109600 105918 109640
rect 105960 109600 106000 109640
rect 120752 109600 120792 109640
rect 120834 109600 120874 109640
rect 120916 109600 120956 109640
rect 120998 109600 121038 109640
rect 121080 109600 121120 109640
rect 135872 109600 135912 109640
rect 135954 109600 135994 109640
rect 136036 109600 136076 109640
rect 136118 109600 136158 109640
rect 136200 109600 136240 109640
rect 150992 109600 151032 109640
rect 151074 109600 151114 109640
rect 151156 109600 151196 109640
rect 151238 109600 151278 109640
rect 151320 109600 151360 109640
rect 104392 108844 104432 108884
rect 104474 108844 104514 108884
rect 104556 108844 104596 108884
rect 104638 108844 104678 108884
rect 104720 108844 104760 108884
rect 119512 108844 119552 108884
rect 119594 108844 119634 108884
rect 119676 108844 119716 108884
rect 119758 108844 119798 108884
rect 119840 108844 119880 108884
rect 134632 108844 134672 108884
rect 134714 108844 134754 108884
rect 134796 108844 134836 108884
rect 134878 108844 134918 108884
rect 134960 108844 135000 108884
rect 149752 108844 149792 108884
rect 149834 108844 149874 108884
rect 149916 108844 149956 108884
rect 149998 108844 150038 108884
rect 150080 108844 150120 108884
rect 105632 108088 105672 108128
rect 105714 108088 105754 108128
rect 105796 108088 105836 108128
rect 105878 108088 105918 108128
rect 105960 108088 106000 108128
rect 120752 108088 120792 108128
rect 120834 108088 120874 108128
rect 120916 108088 120956 108128
rect 120998 108088 121038 108128
rect 121080 108088 121120 108128
rect 135872 108088 135912 108128
rect 135954 108088 135994 108128
rect 136036 108088 136076 108128
rect 136118 108088 136158 108128
rect 136200 108088 136240 108128
rect 150992 108088 151032 108128
rect 151074 108088 151114 108128
rect 151156 108088 151196 108128
rect 151238 108088 151278 108128
rect 151320 108088 151360 108128
rect 104392 107332 104432 107372
rect 104474 107332 104514 107372
rect 104556 107332 104596 107372
rect 104638 107332 104678 107372
rect 104720 107332 104760 107372
rect 119512 107332 119552 107372
rect 119594 107332 119634 107372
rect 119676 107332 119716 107372
rect 119758 107332 119798 107372
rect 119840 107332 119880 107372
rect 134632 107332 134672 107372
rect 134714 107332 134754 107372
rect 134796 107332 134836 107372
rect 134878 107332 134918 107372
rect 134960 107332 135000 107372
rect 149752 107332 149792 107372
rect 149834 107332 149874 107372
rect 149916 107332 149956 107372
rect 149998 107332 150038 107372
rect 150080 107332 150120 107372
rect 105632 106576 105672 106616
rect 105714 106576 105754 106616
rect 105796 106576 105836 106616
rect 105878 106576 105918 106616
rect 105960 106576 106000 106616
rect 120752 106576 120792 106616
rect 120834 106576 120874 106616
rect 120916 106576 120956 106616
rect 120998 106576 121038 106616
rect 121080 106576 121120 106616
rect 135872 106576 135912 106616
rect 135954 106576 135994 106616
rect 136036 106576 136076 106616
rect 136118 106576 136158 106616
rect 136200 106576 136240 106616
rect 150992 106576 151032 106616
rect 151074 106576 151114 106616
rect 151156 106576 151196 106616
rect 151238 106576 151278 106616
rect 151320 106576 151360 106616
rect 104392 105820 104432 105860
rect 104474 105820 104514 105860
rect 104556 105820 104596 105860
rect 104638 105820 104678 105860
rect 104720 105820 104760 105860
rect 119512 105820 119552 105860
rect 119594 105820 119634 105860
rect 119676 105820 119716 105860
rect 119758 105820 119798 105860
rect 119840 105820 119880 105860
rect 134632 105820 134672 105860
rect 134714 105820 134754 105860
rect 134796 105820 134836 105860
rect 134878 105820 134918 105860
rect 134960 105820 135000 105860
rect 149752 105820 149792 105860
rect 149834 105820 149874 105860
rect 149916 105820 149956 105860
rect 149998 105820 150038 105860
rect 150080 105820 150120 105860
rect 105632 105064 105672 105104
rect 105714 105064 105754 105104
rect 105796 105064 105836 105104
rect 105878 105064 105918 105104
rect 105960 105064 106000 105104
rect 120752 105064 120792 105104
rect 120834 105064 120874 105104
rect 120916 105064 120956 105104
rect 120998 105064 121038 105104
rect 121080 105064 121120 105104
rect 135872 105064 135912 105104
rect 135954 105064 135994 105104
rect 136036 105064 136076 105104
rect 136118 105064 136158 105104
rect 136200 105064 136240 105104
rect 150992 105064 151032 105104
rect 151074 105064 151114 105104
rect 151156 105064 151196 105104
rect 151238 105064 151278 105104
rect 151320 105064 151360 105104
rect 104392 104308 104432 104348
rect 104474 104308 104514 104348
rect 104556 104308 104596 104348
rect 104638 104308 104678 104348
rect 104720 104308 104760 104348
rect 119512 104308 119552 104348
rect 119594 104308 119634 104348
rect 119676 104308 119716 104348
rect 119758 104308 119798 104348
rect 119840 104308 119880 104348
rect 134632 104308 134672 104348
rect 134714 104308 134754 104348
rect 134796 104308 134836 104348
rect 134878 104308 134918 104348
rect 134960 104308 135000 104348
rect 149752 104308 149792 104348
rect 149834 104308 149874 104348
rect 149916 104308 149956 104348
rect 149998 104308 150038 104348
rect 150080 104308 150120 104348
rect 105632 103552 105672 103592
rect 105714 103552 105754 103592
rect 105796 103552 105836 103592
rect 105878 103552 105918 103592
rect 105960 103552 106000 103592
rect 120752 103552 120792 103592
rect 120834 103552 120874 103592
rect 120916 103552 120956 103592
rect 120998 103552 121038 103592
rect 121080 103552 121120 103592
rect 135872 103552 135912 103592
rect 135954 103552 135994 103592
rect 136036 103552 136076 103592
rect 136118 103552 136158 103592
rect 136200 103552 136240 103592
rect 150992 103552 151032 103592
rect 151074 103552 151114 103592
rect 151156 103552 151196 103592
rect 151238 103552 151278 103592
rect 151320 103552 151360 103592
rect 104392 102796 104432 102836
rect 104474 102796 104514 102836
rect 104556 102796 104596 102836
rect 104638 102796 104678 102836
rect 104720 102796 104760 102836
rect 119512 102796 119552 102836
rect 119594 102796 119634 102836
rect 119676 102796 119716 102836
rect 119758 102796 119798 102836
rect 119840 102796 119880 102836
rect 134632 102796 134672 102836
rect 134714 102796 134754 102836
rect 134796 102796 134836 102836
rect 134878 102796 134918 102836
rect 134960 102796 135000 102836
rect 149752 102796 149792 102836
rect 149834 102796 149874 102836
rect 149916 102796 149956 102836
rect 149998 102796 150038 102836
rect 150080 102796 150120 102836
rect 105632 102040 105672 102080
rect 105714 102040 105754 102080
rect 105796 102040 105836 102080
rect 105878 102040 105918 102080
rect 105960 102040 106000 102080
rect 120752 102040 120792 102080
rect 120834 102040 120874 102080
rect 120916 102040 120956 102080
rect 120998 102040 121038 102080
rect 121080 102040 121120 102080
rect 135872 102040 135912 102080
rect 135954 102040 135994 102080
rect 136036 102040 136076 102080
rect 136118 102040 136158 102080
rect 136200 102040 136240 102080
rect 150992 102040 151032 102080
rect 151074 102040 151114 102080
rect 151156 102040 151196 102080
rect 151238 102040 151278 102080
rect 151320 102040 151360 102080
rect 104392 101284 104432 101324
rect 104474 101284 104514 101324
rect 104556 101284 104596 101324
rect 104638 101284 104678 101324
rect 104720 101284 104760 101324
rect 119512 101284 119552 101324
rect 119594 101284 119634 101324
rect 119676 101284 119716 101324
rect 119758 101284 119798 101324
rect 119840 101284 119880 101324
rect 134632 101284 134672 101324
rect 134714 101284 134754 101324
rect 134796 101284 134836 101324
rect 134878 101284 134918 101324
rect 134960 101284 135000 101324
rect 149752 101284 149792 101324
rect 149834 101284 149874 101324
rect 149916 101284 149956 101324
rect 149998 101284 150038 101324
rect 150080 101284 150120 101324
rect 105632 100528 105672 100568
rect 105714 100528 105754 100568
rect 105796 100528 105836 100568
rect 105878 100528 105918 100568
rect 105960 100528 106000 100568
rect 120752 100528 120792 100568
rect 120834 100528 120874 100568
rect 120916 100528 120956 100568
rect 120998 100528 121038 100568
rect 121080 100528 121120 100568
rect 135872 100528 135912 100568
rect 135954 100528 135994 100568
rect 136036 100528 136076 100568
rect 136118 100528 136158 100568
rect 136200 100528 136240 100568
rect 150992 100528 151032 100568
rect 151074 100528 151114 100568
rect 151156 100528 151196 100568
rect 151238 100528 151278 100568
rect 151320 100528 151360 100568
rect 104392 99772 104432 99812
rect 104474 99772 104514 99812
rect 104556 99772 104596 99812
rect 104638 99772 104678 99812
rect 104720 99772 104760 99812
rect 119512 99772 119552 99812
rect 119594 99772 119634 99812
rect 119676 99772 119716 99812
rect 119758 99772 119798 99812
rect 119840 99772 119880 99812
rect 134632 99772 134672 99812
rect 134714 99772 134754 99812
rect 134796 99772 134836 99812
rect 134878 99772 134918 99812
rect 134960 99772 135000 99812
rect 149752 99772 149792 99812
rect 149834 99772 149874 99812
rect 149916 99772 149956 99812
rect 149998 99772 150038 99812
rect 150080 99772 150120 99812
rect 105632 99016 105672 99056
rect 105714 99016 105754 99056
rect 105796 99016 105836 99056
rect 105878 99016 105918 99056
rect 105960 99016 106000 99056
rect 120752 99016 120792 99056
rect 120834 99016 120874 99056
rect 120916 99016 120956 99056
rect 120998 99016 121038 99056
rect 121080 99016 121120 99056
rect 135872 99016 135912 99056
rect 135954 99016 135994 99056
rect 136036 99016 136076 99056
rect 136118 99016 136158 99056
rect 136200 99016 136240 99056
rect 150992 99016 151032 99056
rect 151074 99016 151114 99056
rect 151156 99016 151196 99056
rect 151238 99016 151278 99056
rect 151320 99016 151360 99056
rect 104392 98260 104432 98300
rect 104474 98260 104514 98300
rect 104556 98260 104596 98300
rect 104638 98260 104678 98300
rect 104720 98260 104760 98300
rect 119512 98260 119552 98300
rect 119594 98260 119634 98300
rect 119676 98260 119716 98300
rect 119758 98260 119798 98300
rect 119840 98260 119880 98300
rect 134632 98260 134672 98300
rect 134714 98260 134754 98300
rect 134796 98260 134836 98300
rect 134878 98260 134918 98300
rect 134960 98260 135000 98300
rect 149752 98260 149792 98300
rect 149834 98260 149874 98300
rect 149916 98260 149956 98300
rect 149998 98260 150038 98300
rect 150080 98260 150120 98300
rect 105632 97504 105672 97544
rect 105714 97504 105754 97544
rect 105796 97504 105836 97544
rect 105878 97504 105918 97544
rect 105960 97504 106000 97544
rect 120752 97504 120792 97544
rect 120834 97504 120874 97544
rect 120916 97504 120956 97544
rect 120998 97504 121038 97544
rect 121080 97504 121120 97544
rect 135872 97504 135912 97544
rect 135954 97504 135994 97544
rect 136036 97504 136076 97544
rect 136118 97504 136158 97544
rect 136200 97504 136240 97544
rect 150992 97504 151032 97544
rect 151074 97504 151114 97544
rect 151156 97504 151196 97544
rect 151238 97504 151278 97544
rect 151320 97504 151360 97544
rect 104392 96748 104432 96788
rect 104474 96748 104514 96788
rect 104556 96748 104596 96788
rect 104638 96748 104678 96788
rect 104720 96748 104760 96788
rect 119512 96748 119552 96788
rect 119594 96748 119634 96788
rect 119676 96748 119716 96788
rect 119758 96748 119798 96788
rect 119840 96748 119880 96788
rect 134632 96748 134672 96788
rect 134714 96748 134754 96788
rect 134796 96748 134836 96788
rect 134878 96748 134918 96788
rect 134960 96748 135000 96788
rect 149752 96748 149792 96788
rect 149834 96748 149874 96788
rect 149916 96748 149956 96788
rect 149998 96748 150038 96788
rect 150080 96748 150120 96788
rect 105632 95992 105672 96032
rect 105714 95992 105754 96032
rect 105796 95992 105836 96032
rect 105878 95992 105918 96032
rect 105960 95992 106000 96032
rect 120752 95992 120792 96032
rect 120834 95992 120874 96032
rect 120916 95992 120956 96032
rect 120998 95992 121038 96032
rect 121080 95992 121120 96032
rect 135872 95992 135912 96032
rect 135954 95992 135994 96032
rect 136036 95992 136076 96032
rect 136118 95992 136158 96032
rect 136200 95992 136240 96032
rect 150992 95992 151032 96032
rect 151074 95992 151114 96032
rect 151156 95992 151196 96032
rect 151238 95992 151278 96032
rect 151320 95992 151360 96032
rect 104392 95236 104432 95276
rect 104474 95236 104514 95276
rect 104556 95236 104596 95276
rect 104638 95236 104678 95276
rect 104720 95236 104760 95276
rect 119512 95236 119552 95276
rect 119594 95236 119634 95276
rect 119676 95236 119716 95276
rect 119758 95236 119798 95276
rect 119840 95236 119880 95276
rect 134632 95236 134672 95276
rect 134714 95236 134754 95276
rect 134796 95236 134836 95276
rect 134878 95236 134918 95276
rect 134960 95236 135000 95276
rect 149752 95236 149792 95276
rect 149834 95236 149874 95276
rect 149916 95236 149956 95276
rect 149998 95236 150038 95276
rect 150080 95236 150120 95276
rect 105632 94480 105672 94520
rect 105714 94480 105754 94520
rect 105796 94480 105836 94520
rect 105878 94480 105918 94520
rect 105960 94480 106000 94520
rect 120752 94480 120792 94520
rect 120834 94480 120874 94520
rect 120916 94480 120956 94520
rect 120998 94480 121038 94520
rect 121080 94480 121120 94520
rect 135872 94480 135912 94520
rect 135954 94480 135994 94520
rect 136036 94480 136076 94520
rect 136118 94480 136158 94520
rect 136200 94480 136240 94520
rect 150992 94480 151032 94520
rect 151074 94480 151114 94520
rect 151156 94480 151196 94520
rect 151238 94480 151278 94520
rect 151320 94480 151360 94520
rect 104392 93724 104432 93764
rect 104474 93724 104514 93764
rect 104556 93724 104596 93764
rect 104638 93724 104678 93764
rect 104720 93724 104760 93764
rect 119512 93724 119552 93764
rect 119594 93724 119634 93764
rect 119676 93724 119716 93764
rect 119758 93724 119798 93764
rect 119840 93724 119880 93764
rect 134632 93724 134672 93764
rect 134714 93724 134754 93764
rect 134796 93724 134836 93764
rect 134878 93724 134918 93764
rect 134960 93724 135000 93764
rect 149752 93724 149792 93764
rect 149834 93724 149874 93764
rect 149916 93724 149956 93764
rect 149998 93724 150038 93764
rect 150080 93724 150120 93764
rect 105632 92968 105672 93008
rect 105714 92968 105754 93008
rect 105796 92968 105836 93008
rect 105878 92968 105918 93008
rect 105960 92968 106000 93008
rect 120752 92968 120792 93008
rect 120834 92968 120874 93008
rect 120916 92968 120956 93008
rect 120998 92968 121038 93008
rect 121080 92968 121120 93008
rect 135872 92968 135912 93008
rect 135954 92968 135994 93008
rect 136036 92968 136076 93008
rect 136118 92968 136158 93008
rect 136200 92968 136240 93008
rect 150992 92968 151032 93008
rect 151074 92968 151114 93008
rect 151156 92968 151196 93008
rect 151238 92968 151278 93008
rect 151320 92968 151360 93008
rect 104392 92212 104432 92252
rect 104474 92212 104514 92252
rect 104556 92212 104596 92252
rect 104638 92212 104678 92252
rect 104720 92212 104760 92252
rect 119512 92212 119552 92252
rect 119594 92212 119634 92252
rect 119676 92212 119716 92252
rect 119758 92212 119798 92252
rect 119840 92212 119880 92252
rect 134632 92212 134672 92252
rect 134714 92212 134754 92252
rect 134796 92212 134836 92252
rect 134878 92212 134918 92252
rect 134960 92212 135000 92252
rect 149752 92212 149792 92252
rect 149834 92212 149874 92252
rect 149916 92212 149956 92252
rect 149998 92212 150038 92252
rect 150080 92212 150120 92252
rect 105632 91456 105672 91496
rect 105714 91456 105754 91496
rect 105796 91456 105836 91496
rect 105878 91456 105918 91496
rect 105960 91456 106000 91496
rect 120752 91456 120792 91496
rect 120834 91456 120874 91496
rect 120916 91456 120956 91496
rect 120998 91456 121038 91496
rect 121080 91456 121120 91496
rect 135872 91456 135912 91496
rect 135954 91456 135994 91496
rect 136036 91456 136076 91496
rect 136118 91456 136158 91496
rect 136200 91456 136240 91496
rect 150992 91456 151032 91496
rect 151074 91456 151114 91496
rect 151156 91456 151196 91496
rect 151238 91456 151278 91496
rect 151320 91456 151360 91496
rect 104392 90700 104432 90740
rect 104474 90700 104514 90740
rect 104556 90700 104596 90740
rect 104638 90700 104678 90740
rect 104720 90700 104760 90740
rect 119512 90700 119552 90740
rect 119594 90700 119634 90740
rect 119676 90700 119716 90740
rect 119758 90700 119798 90740
rect 119840 90700 119880 90740
rect 134632 90700 134672 90740
rect 134714 90700 134754 90740
rect 134796 90700 134836 90740
rect 134878 90700 134918 90740
rect 134960 90700 135000 90740
rect 149752 90700 149792 90740
rect 149834 90700 149874 90740
rect 149916 90700 149956 90740
rect 149998 90700 150038 90740
rect 150080 90700 150120 90740
rect 105632 89944 105672 89984
rect 105714 89944 105754 89984
rect 105796 89944 105836 89984
rect 105878 89944 105918 89984
rect 105960 89944 106000 89984
rect 120752 89944 120792 89984
rect 120834 89944 120874 89984
rect 120916 89944 120956 89984
rect 120998 89944 121038 89984
rect 121080 89944 121120 89984
rect 135872 89944 135912 89984
rect 135954 89944 135994 89984
rect 136036 89944 136076 89984
rect 136118 89944 136158 89984
rect 136200 89944 136240 89984
rect 150992 89944 151032 89984
rect 151074 89944 151114 89984
rect 151156 89944 151196 89984
rect 151238 89944 151278 89984
rect 151320 89944 151360 89984
rect 104392 89188 104432 89228
rect 104474 89188 104514 89228
rect 104556 89188 104596 89228
rect 104638 89188 104678 89228
rect 104720 89188 104760 89228
rect 119512 89188 119552 89228
rect 119594 89188 119634 89228
rect 119676 89188 119716 89228
rect 119758 89188 119798 89228
rect 119840 89188 119880 89228
rect 134632 89188 134672 89228
rect 134714 89188 134754 89228
rect 134796 89188 134836 89228
rect 134878 89188 134918 89228
rect 134960 89188 135000 89228
rect 149752 89188 149792 89228
rect 149834 89188 149874 89228
rect 149916 89188 149956 89228
rect 149998 89188 150038 89228
rect 150080 89188 150120 89228
rect 105632 88432 105672 88472
rect 105714 88432 105754 88472
rect 105796 88432 105836 88472
rect 105878 88432 105918 88472
rect 105960 88432 106000 88472
rect 120752 88432 120792 88472
rect 120834 88432 120874 88472
rect 120916 88432 120956 88472
rect 120998 88432 121038 88472
rect 121080 88432 121120 88472
rect 135872 88432 135912 88472
rect 135954 88432 135994 88472
rect 136036 88432 136076 88472
rect 136118 88432 136158 88472
rect 136200 88432 136240 88472
rect 150992 88432 151032 88472
rect 151074 88432 151114 88472
rect 151156 88432 151196 88472
rect 151238 88432 151278 88472
rect 151320 88432 151360 88472
rect 104392 87676 104432 87716
rect 104474 87676 104514 87716
rect 104556 87676 104596 87716
rect 104638 87676 104678 87716
rect 104720 87676 104760 87716
rect 119512 87676 119552 87716
rect 119594 87676 119634 87716
rect 119676 87676 119716 87716
rect 119758 87676 119798 87716
rect 119840 87676 119880 87716
rect 134632 87676 134672 87716
rect 134714 87676 134754 87716
rect 134796 87676 134836 87716
rect 134878 87676 134918 87716
rect 134960 87676 135000 87716
rect 149752 87676 149792 87716
rect 149834 87676 149874 87716
rect 149916 87676 149956 87716
rect 149998 87676 150038 87716
rect 150080 87676 150120 87716
rect 105632 86920 105672 86960
rect 105714 86920 105754 86960
rect 105796 86920 105836 86960
rect 105878 86920 105918 86960
rect 105960 86920 106000 86960
rect 120752 86920 120792 86960
rect 120834 86920 120874 86960
rect 120916 86920 120956 86960
rect 120998 86920 121038 86960
rect 121080 86920 121120 86960
rect 135872 86920 135912 86960
rect 135954 86920 135994 86960
rect 136036 86920 136076 86960
rect 136118 86920 136158 86960
rect 136200 86920 136240 86960
rect 150992 86920 151032 86960
rect 151074 86920 151114 86960
rect 151156 86920 151196 86960
rect 151238 86920 151278 86960
rect 151320 86920 151360 86960
rect 104392 86164 104432 86204
rect 104474 86164 104514 86204
rect 104556 86164 104596 86204
rect 104638 86164 104678 86204
rect 104720 86164 104760 86204
rect 119512 86164 119552 86204
rect 119594 86164 119634 86204
rect 119676 86164 119716 86204
rect 119758 86164 119798 86204
rect 119840 86164 119880 86204
rect 134632 86164 134672 86204
rect 134714 86164 134754 86204
rect 134796 86164 134836 86204
rect 134878 86164 134918 86204
rect 134960 86164 135000 86204
rect 149752 86164 149792 86204
rect 149834 86164 149874 86204
rect 149916 86164 149956 86204
rect 149998 86164 150038 86204
rect 150080 86164 150120 86204
rect 105632 85408 105672 85448
rect 105714 85408 105754 85448
rect 105796 85408 105836 85448
rect 105878 85408 105918 85448
rect 105960 85408 106000 85448
rect 120752 85408 120792 85448
rect 120834 85408 120874 85448
rect 120916 85408 120956 85448
rect 120998 85408 121038 85448
rect 121080 85408 121120 85448
rect 135872 85408 135912 85448
rect 135954 85408 135994 85448
rect 136036 85408 136076 85448
rect 136118 85408 136158 85448
rect 136200 85408 136240 85448
rect 150992 85408 151032 85448
rect 151074 85408 151114 85448
rect 151156 85408 151196 85448
rect 151238 85408 151278 85448
rect 151320 85408 151360 85448
rect 104392 84652 104432 84692
rect 104474 84652 104514 84692
rect 104556 84652 104596 84692
rect 104638 84652 104678 84692
rect 104720 84652 104760 84692
rect 119512 84652 119552 84692
rect 119594 84652 119634 84692
rect 119676 84652 119716 84692
rect 119758 84652 119798 84692
rect 119840 84652 119880 84692
rect 134632 84652 134672 84692
rect 134714 84652 134754 84692
rect 134796 84652 134836 84692
rect 134878 84652 134918 84692
rect 134960 84652 135000 84692
rect 149752 84652 149792 84692
rect 149834 84652 149874 84692
rect 149916 84652 149956 84692
rect 149998 84652 150038 84692
rect 150080 84652 150120 84692
rect 105632 83896 105672 83936
rect 105714 83896 105754 83936
rect 105796 83896 105836 83936
rect 105878 83896 105918 83936
rect 105960 83896 106000 83936
rect 120752 83896 120792 83936
rect 120834 83896 120874 83936
rect 120916 83896 120956 83936
rect 120998 83896 121038 83936
rect 121080 83896 121120 83936
rect 135872 83896 135912 83936
rect 135954 83896 135994 83936
rect 136036 83896 136076 83936
rect 136118 83896 136158 83936
rect 136200 83896 136240 83936
rect 150992 83896 151032 83936
rect 151074 83896 151114 83936
rect 151156 83896 151196 83936
rect 151238 83896 151278 83936
rect 151320 83896 151360 83936
rect 104392 83140 104432 83180
rect 104474 83140 104514 83180
rect 104556 83140 104596 83180
rect 104638 83140 104678 83180
rect 104720 83140 104760 83180
rect 119512 83140 119552 83180
rect 119594 83140 119634 83180
rect 119676 83140 119716 83180
rect 119758 83140 119798 83180
rect 119840 83140 119880 83180
rect 134632 83140 134672 83180
rect 134714 83140 134754 83180
rect 134796 83140 134836 83180
rect 134878 83140 134918 83180
rect 134960 83140 135000 83180
rect 149752 83140 149792 83180
rect 149834 83140 149874 83180
rect 149916 83140 149956 83180
rect 149998 83140 150038 83180
rect 150080 83140 150120 83180
rect 105632 82384 105672 82424
rect 105714 82384 105754 82424
rect 105796 82384 105836 82424
rect 105878 82384 105918 82424
rect 105960 82384 106000 82424
rect 120752 82384 120792 82424
rect 120834 82384 120874 82424
rect 120916 82384 120956 82424
rect 120998 82384 121038 82424
rect 121080 82384 121120 82424
rect 135872 82384 135912 82424
rect 135954 82384 135994 82424
rect 136036 82384 136076 82424
rect 136118 82384 136158 82424
rect 136200 82384 136240 82424
rect 150992 82384 151032 82424
rect 151074 82384 151114 82424
rect 151156 82384 151196 82424
rect 151238 82384 151278 82424
rect 151320 82384 151360 82424
rect 104392 81628 104432 81668
rect 104474 81628 104514 81668
rect 104556 81628 104596 81668
rect 104638 81628 104678 81668
rect 104720 81628 104760 81668
rect 119512 81628 119552 81668
rect 119594 81628 119634 81668
rect 119676 81628 119716 81668
rect 119758 81628 119798 81668
rect 119840 81628 119880 81668
rect 134632 81628 134672 81668
rect 134714 81628 134754 81668
rect 134796 81628 134836 81668
rect 134878 81628 134918 81668
rect 134960 81628 135000 81668
rect 149752 81628 149792 81668
rect 149834 81628 149874 81668
rect 149916 81628 149956 81668
rect 149998 81628 150038 81668
rect 150080 81628 150120 81668
rect 105632 80872 105672 80912
rect 105714 80872 105754 80912
rect 105796 80872 105836 80912
rect 105878 80872 105918 80912
rect 105960 80872 106000 80912
rect 120752 80872 120792 80912
rect 120834 80872 120874 80912
rect 120916 80872 120956 80912
rect 120998 80872 121038 80912
rect 121080 80872 121120 80912
rect 135872 80872 135912 80912
rect 135954 80872 135994 80912
rect 136036 80872 136076 80912
rect 136118 80872 136158 80912
rect 136200 80872 136240 80912
rect 150992 80872 151032 80912
rect 151074 80872 151114 80912
rect 151156 80872 151196 80912
rect 151238 80872 151278 80912
rect 151320 80872 151360 80912
rect 104392 80116 104432 80156
rect 104474 80116 104514 80156
rect 104556 80116 104596 80156
rect 104638 80116 104678 80156
rect 104720 80116 104760 80156
rect 119512 80116 119552 80156
rect 119594 80116 119634 80156
rect 119676 80116 119716 80156
rect 119758 80116 119798 80156
rect 119840 80116 119880 80156
rect 134632 80116 134672 80156
rect 134714 80116 134754 80156
rect 134796 80116 134836 80156
rect 134878 80116 134918 80156
rect 134960 80116 135000 80156
rect 149752 80116 149792 80156
rect 149834 80116 149874 80156
rect 149916 80116 149956 80156
rect 149998 80116 150038 80156
rect 150080 80116 150120 80156
rect 105632 79360 105672 79400
rect 105714 79360 105754 79400
rect 105796 79360 105836 79400
rect 105878 79360 105918 79400
rect 105960 79360 106000 79400
rect 120752 79360 120792 79400
rect 120834 79360 120874 79400
rect 120916 79360 120956 79400
rect 120998 79360 121038 79400
rect 121080 79360 121120 79400
rect 135872 79360 135912 79400
rect 135954 79360 135994 79400
rect 136036 79360 136076 79400
rect 136118 79360 136158 79400
rect 136200 79360 136240 79400
rect 150992 79360 151032 79400
rect 151074 79360 151114 79400
rect 151156 79360 151196 79400
rect 151238 79360 151278 79400
rect 151320 79360 151360 79400
rect 104392 78604 104432 78644
rect 104474 78604 104514 78644
rect 104556 78604 104596 78644
rect 104638 78604 104678 78644
rect 104720 78604 104760 78644
rect 119512 78604 119552 78644
rect 119594 78604 119634 78644
rect 119676 78604 119716 78644
rect 119758 78604 119798 78644
rect 119840 78604 119880 78644
rect 134632 78604 134672 78644
rect 134714 78604 134754 78644
rect 134796 78604 134836 78644
rect 134878 78604 134918 78644
rect 134960 78604 135000 78644
rect 149752 78604 149792 78644
rect 149834 78604 149874 78644
rect 149916 78604 149956 78644
rect 149998 78604 150038 78644
rect 150080 78604 150120 78644
rect 105632 77848 105672 77888
rect 105714 77848 105754 77888
rect 105796 77848 105836 77888
rect 105878 77848 105918 77888
rect 105960 77848 106000 77888
rect 120752 77848 120792 77888
rect 120834 77848 120874 77888
rect 120916 77848 120956 77888
rect 120998 77848 121038 77888
rect 121080 77848 121120 77888
rect 135872 77848 135912 77888
rect 135954 77848 135994 77888
rect 136036 77848 136076 77888
rect 136118 77848 136158 77888
rect 136200 77848 136240 77888
rect 150992 77848 151032 77888
rect 151074 77848 151114 77888
rect 151156 77848 151196 77888
rect 151238 77848 151278 77888
rect 151320 77848 151360 77888
rect 104392 77092 104432 77132
rect 104474 77092 104514 77132
rect 104556 77092 104596 77132
rect 104638 77092 104678 77132
rect 104720 77092 104760 77132
rect 119512 77092 119552 77132
rect 119594 77092 119634 77132
rect 119676 77092 119716 77132
rect 119758 77092 119798 77132
rect 119840 77092 119880 77132
rect 134632 77092 134672 77132
rect 134714 77092 134754 77132
rect 134796 77092 134836 77132
rect 134878 77092 134918 77132
rect 134960 77092 135000 77132
rect 149752 77092 149792 77132
rect 149834 77092 149874 77132
rect 149916 77092 149956 77132
rect 149998 77092 150038 77132
rect 150080 77092 150120 77132
rect 105632 76336 105672 76376
rect 105714 76336 105754 76376
rect 105796 76336 105836 76376
rect 105878 76336 105918 76376
rect 105960 76336 106000 76376
rect 120752 76336 120792 76376
rect 120834 76336 120874 76376
rect 120916 76336 120956 76376
rect 120998 76336 121038 76376
rect 121080 76336 121120 76376
rect 135872 76336 135912 76376
rect 135954 76336 135994 76376
rect 136036 76336 136076 76376
rect 136118 76336 136158 76376
rect 136200 76336 136240 76376
rect 150992 76336 151032 76376
rect 151074 76336 151114 76376
rect 151156 76336 151196 76376
rect 151238 76336 151278 76376
rect 151320 76336 151360 76376
rect 104392 75580 104432 75620
rect 104474 75580 104514 75620
rect 104556 75580 104596 75620
rect 104638 75580 104678 75620
rect 104720 75580 104760 75620
rect 119512 75580 119552 75620
rect 119594 75580 119634 75620
rect 119676 75580 119716 75620
rect 119758 75580 119798 75620
rect 119840 75580 119880 75620
rect 134632 75580 134672 75620
rect 134714 75580 134754 75620
rect 134796 75580 134836 75620
rect 134878 75580 134918 75620
rect 134960 75580 135000 75620
rect 149752 75580 149792 75620
rect 149834 75580 149874 75620
rect 149916 75580 149956 75620
rect 149998 75580 150038 75620
rect 150080 75580 150120 75620
rect 105632 74824 105672 74864
rect 105714 74824 105754 74864
rect 105796 74824 105836 74864
rect 105878 74824 105918 74864
rect 105960 74824 106000 74864
rect 120752 74824 120792 74864
rect 120834 74824 120874 74864
rect 120916 74824 120956 74864
rect 120998 74824 121038 74864
rect 121080 74824 121120 74864
rect 135872 74824 135912 74864
rect 135954 74824 135994 74864
rect 136036 74824 136076 74864
rect 136118 74824 136158 74864
rect 136200 74824 136240 74864
rect 150992 74824 151032 74864
rect 151074 74824 151114 74864
rect 151156 74824 151196 74864
rect 151238 74824 151278 74864
rect 151320 74824 151360 74864
rect 104392 74068 104432 74108
rect 104474 74068 104514 74108
rect 104556 74068 104596 74108
rect 104638 74068 104678 74108
rect 104720 74068 104760 74108
rect 119512 74068 119552 74108
rect 119594 74068 119634 74108
rect 119676 74068 119716 74108
rect 119758 74068 119798 74108
rect 119840 74068 119880 74108
rect 134632 74068 134672 74108
rect 134714 74068 134754 74108
rect 134796 74068 134836 74108
rect 134878 74068 134918 74108
rect 134960 74068 135000 74108
rect 149752 74068 149792 74108
rect 149834 74068 149874 74108
rect 149916 74068 149956 74108
rect 149998 74068 150038 74108
rect 150080 74068 150120 74108
rect 105632 73312 105672 73352
rect 105714 73312 105754 73352
rect 105796 73312 105836 73352
rect 105878 73312 105918 73352
rect 105960 73312 106000 73352
rect 120752 73312 120792 73352
rect 120834 73312 120874 73352
rect 120916 73312 120956 73352
rect 120998 73312 121038 73352
rect 121080 73312 121120 73352
rect 135872 73312 135912 73352
rect 135954 73312 135994 73352
rect 136036 73312 136076 73352
rect 136118 73312 136158 73352
rect 136200 73312 136240 73352
rect 150992 73312 151032 73352
rect 151074 73312 151114 73352
rect 151156 73312 151196 73352
rect 151238 73312 151278 73352
rect 151320 73312 151360 73352
rect 104392 72556 104432 72596
rect 104474 72556 104514 72596
rect 104556 72556 104596 72596
rect 104638 72556 104678 72596
rect 104720 72556 104760 72596
rect 119512 72556 119552 72596
rect 119594 72556 119634 72596
rect 119676 72556 119716 72596
rect 119758 72556 119798 72596
rect 119840 72556 119880 72596
rect 134632 72556 134672 72596
rect 134714 72556 134754 72596
rect 134796 72556 134836 72596
rect 134878 72556 134918 72596
rect 134960 72556 135000 72596
rect 149752 72556 149792 72596
rect 149834 72556 149874 72596
rect 149916 72556 149956 72596
rect 149998 72556 150038 72596
rect 150080 72556 150120 72596
rect 105632 71800 105672 71840
rect 105714 71800 105754 71840
rect 105796 71800 105836 71840
rect 105878 71800 105918 71840
rect 105960 71800 106000 71840
rect 120752 71800 120792 71840
rect 120834 71800 120874 71840
rect 120916 71800 120956 71840
rect 120998 71800 121038 71840
rect 121080 71800 121120 71840
rect 135872 71800 135912 71840
rect 135954 71800 135994 71840
rect 136036 71800 136076 71840
rect 136118 71800 136158 71840
rect 136200 71800 136240 71840
rect 150992 71800 151032 71840
rect 151074 71800 151114 71840
rect 151156 71800 151196 71840
rect 151238 71800 151278 71840
rect 151320 71800 151360 71840
rect 151564 64156 151604 64196
<< metal3 >>
rect 71971 159412 71980 159452
rect 72020 159412 103660 159452
rect 103700 159412 103709 159452
rect 104035 159412 104044 159452
rect 104084 159412 135724 159452
rect 135764 159412 135773 159452
rect 88003 159328 88012 159368
rect 88052 159328 119692 159368
rect 119732 159328 119741 159368
rect 64099 152020 64108 152060
rect 64148 152020 160032 152060
rect 75383 151936 75392 151976
rect 75432 151936 75474 151976
rect 75514 151936 75556 151976
rect 75596 151936 75638 151976
rect 75678 151936 75720 151976
rect 75760 151936 75769 151976
rect 90503 151936 90512 151976
rect 90552 151936 90594 151976
rect 90634 151936 90676 151976
rect 90716 151936 90758 151976
rect 90798 151936 90840 151976
rect 90880 151936 90889 151976
rect 105623 151936 105632 151976
rect 105672 151936 105714 151976
rect 105754 151936 105796 151976
rect 105836 151936 105878 151976
rect 105918 151936 105960 151976
rect 106000 151936 106009 151976
rect 120743 151936 120752 151976
rect 120792 151936 120834 151976
rect 120874 151936 120916 151976
rect 120956 151936 120998 151976
rect 121038 151936 121080 151976
rect 121120 151936 121129 151976
rect 135863 151936 135872 151976
rect 135912 151936 135954 151976
rect 135994 151936 136036 151976
rect 136076 151936 136118 151976
rect 136158 151936 136200 151976
rect 136240 151936 136249 151976
rect 150983 151936 150992 151976
rect 151032 151936 151074 151976
rect 151114 151936 151156 151976
rect 151196 151936 151238 151976
rect 151278 151936 151320 151976
rect 151360 151936 151369 151976
rect 74143 151180 74152 151220
rect 74192 151180 74234 151220
rect 74274 151180 74316 151220
rect 74356 151180 74398 151220
rect 74438 151180 74480 151220
rect 74520 151180 74529 151220
rect 89263 151180 89272 151220
rect 89312 151180 89354 151220
rect 89394 151180 89436 151220
rect 89476 151180 89518 151220
rect 89558 151180 89600 151220
rect 89640 151180 89649 151220
rect 104383 151180 104392 151220
rect 104432 151180 104474 151220
rect 104514 151180 104556 151220
rect 104596 151180 104638 151220
rect 104678 151180 104720 151220
rect 104760 151180 104769 151220
rect 119503 151180 119512 151220
rect 119552 151180 119594 151220
rect 119634 151180 119676 151220
rect 119716 151180 119758 151220
rect 119798 151180 119840 151220
rect 119880 151180 119889 151220
rect 134623 151180 134632 151220
rect 134672 151180 134714 151220
rect 134754 151180 134796 151220
rect 134836 151180 134878 151220
rect 134918 151180 134960 151220
rect 135000 151180 135009 151220
rect 149743 151180 149752 151220
rect 149792 151180 149834 151220
rect 149874 151180 149916 151220
rect 149956 151180 149998 151220
rect 150038 151180 150080 151220
rect 150120 151180 150129 151220
rect 75383 150424 75392 150464
rect 75432 150424 75474 150464
rect 75514 150424 75556 150464
rect 75596 150424 75638 150464
rect 75678 150424 75720 150464
rect 75760 150424 75769 150464
rect 90503 150424 90512 150464
rect 90552 150424 90594 150464
rect 90634 150424 90676 150464
rect 90716 150424 90758 150464
rect 90798 150424 90840 150464
rect 90880 150424 90889 150464
rect 105623 150424 105632 150464
rect 105672 150424 105714 150464
rect 105754 150424 105796 150464
rect 105836 150424 105878 150464
rect 105918 150424 105960 150464
rect 106000 150424 106009 150464
rect 120743 150424 120752 150464
rect 120792 150424 120834 150464
rect 120874 150424 120916 150464
rect 120956 150424 120998 150464
rect 121038 150424 121080 150464
rect 121120 150424 121129 150464
rect 135863 150424 135872 150464
rect 135912 150424 135954 150464
rect 135994 150424 136036 150464
rect 136076 150424 136118 150464
rect 136158 150424 136200 150464
rect 136240 150424 136249 150464
rect 150983 150424 150992 150464
rect 151032 150424 151074 150464
rect 151114 150424 151156 150464
rect 151196 150424 151238 150464
rect 151278 150424 151320 150464
rect 151360 150424 151369 150464
rect 74143 149668 74152 149708
rect 74192 149668 74234 149708
rect 74274 149668 74316 149708
rect 74356 149668 74398 149708
rect 74438 149668 74480 149708
rect 74520 149668 74529 149708
rect 89263 149668 89272 149708
rect 89312 149668 89354 149708
rect 89394 149668 89436 149708
rect 89476 149668 89518 149708
rect 89558 149668 89600 149708
rect 89640 149668 89649 149708
rect 104383 149668 104392 149708
rect 104432 149668 104474 149708
rect 104514 149668 104556 149708
rect 104596 149668 104638 149708
rect 104678 149668 104720 149708
rect 104760 149668 104769 149708
rect 119503 149668 119512 149708
rect 119552 149668 119594 149708
rect 119634 149668 119676 149708
rect 119716 149668 119758 149708
rect 119798 149668 119840 149708
rect 119880 149668 119889 149708
rect 134623 149668 134632 149708
rect 134672 149668 134714 149708
rect 134754 149668 134796 149708
rect 134836 149668 134878 149708
rect 134918 149668 134960 149708
rect 135000 149668 135009 149708
rect 149743 149668 149752 149708
rect 149792 149668 149834 149708
rect 149874 149668 149916 149708
rect 149956 149668 149998 149708
rect 150038 149668 150080 149708
rect 150120 149668 150129 149708
rect 75383 148912 75392 148952
rect 75432 148912 75474 148952
rect 75514 148912 75556 148952
rect 75596 148912 75638 148952
rect 75678 148912 75720 148952
rect 75760 148912 75769 148952
rect 90503 148912 90512 148952
rect 90552 148912 90594 148952
rect 90634 148912 90676 148952
rect 90716 148912 90758 148952
rect 90798 148912 90840 148952
rect 90880 148912 90889 148952
rect 105623 148912 105632 148952
rect 105672 148912 105714 148952
rect 105754 148912 105796 148952
rect 105836 148912 105878 148952
rect 105918 148912 105960 148952
rect 106000 148912 106009 148952
rect 120743 148912 120752 148952
rect 120792 148912 120834 148952
rect 120874 148912 120916 148952
rect 120956 148912 120998 148952
rect 121038 148912 121080 148952
rect 121120 148912 121129 148952
rect 135863 148912 135872 148952
rect 135912 148912 135954 148952
rect 135994 148912 136036 148952
rect 136076 148912 136118 148952
rect 136158 148912 136200 148952
rect 136240 148912 136249 148952
rect 150983 148912 150992 148952
rect 151032 148912 151074 148952
rect 151114 148912 151156 148952
rect 151196 148912 151238 148952
rect 151278 148912 151320 148952
rect 151360 148912 151369 148952
rect 74143 148156 74152 148196
rect 74192 148156 74234 148196
rect 74274 148156 74316 148196
rect 74356 148156 74398 148196
rect 74438 148156 74480 148196
rect 74520 148156 74529 148196
rect 89263 148156 89272 148196
rect 89312 148156 89354 148196
rect 89394 148156 89436 148196
rect 89476 148156 89518 148196
rect 89558 148156 89600 148196
rect 89640 148156 89649 148196
rect 104383 148156 104392 148196
rect 104432 148156 104474 148196
rect 104514 148156 104556 148196
rect 104596 148156 104638 148196
rect 104678 148156 104720 148196
rect 104760 148156 104769 148196
rect 119503 148156 119512 148196
rect 119552 148156 119594 148196
rect 119634 148156 119676 148196
rect 119716 148156 119758 148196
rect 119798 148156 119840 148196
rect 119880 148156 119889 148196
rect 134623 148156 134632 148196
rect 134672 148156 134714 148196
rect 134754 148156 134796 148196
rect 134836 148156 134878 148196
rect 134918 148156 134960 148196
rect 135000 148156 135009 148196
rect 149743 148156 149752 148196
rect 149792 148156 149834 148196
rect 149874 148156 149916 148196
rect 149956 148156 149998 148196
rect 150038 148156 150080 148196
rect 150120 148156 150129 148196
rect 75383 147400 75392 147440
rect 75432 147400 75474 147440
rect 75514 147400 75556 147440
rect 75596 147400 75638 147440
rect 75678 147400 75720 147440
rect 75760 147400 75769 147440
rect 90503 147400 90512 147440
rect 90552 147400 90594 147440
rect 90634 147400 90676 147440
rect 90716 147400 90758 147440
rect 90798 147400 90840 147440
rect 90880 147400 90889 147440
rect 105623 147400 105632 147440
rect 105672 147400 105714 147440
rect 105754 147400 105796 147440
rect 105836 147400 105878 147440
rect 105918 147400 105960 147440
rect 106000 147400 106009 147440
rect 120743 147400 120752 147440
rect 120792 147400 120834 147440
rect 120874 147400 120916 147440
rect 120956 147400 120998 147440
rect 121038 147400 121080 147440
rect 121120 147400 121129 147440
rect 135863 147400 135872 147440
rect 135912 147400 135954 147440
rect 135994 147400 136036 147440
rect 136076 147400 136118 147440
rect 136158 147400 136200 147440
rect 136240 147400 136249 147440
rect 150983 147400 150992 147440
rect 151032 147400 151074 147440
rect 151114 147400 151156 147440
rect 151196 147400 151238 147440
rect 151278 147400 151320 147440
rect 151360 147400 151369 147440
rect 74143 146644 74152 146684
rect 74192 146644 74234 146684
rect 74274 146644 74316 146684
rect 74356 146644 74398 146684
rect 74438 146644 74480 146684
rect 74520 146644 74529 146684
rect 89263 146644 89272 146684
rect 89312 146644 89354 146684
rect 89394 146644 89436 146684
rect 89476 146644 89518 146684
rect 89558 146644 89600 146684
rect 89640 146644 89649 146684
rect 104383 146644 104392 146684
rect 104432 146644 104474 146684
rect 104514 146644 104556 146684
rect 104596 146644 104638 146684
rect 104678 146644 104720 146684
rect 104760 146644 104769 146684
rect 119503 146644 119512 146684
rect 119552 146644 119594 146684
rect 119634 146644 119676 146684
rect 119716 146644 119758 146684
rect 119798 146644 119840 146684
rect 119880 146644 119889 146684
rect 134623 146644 134632 146684
rect 134672 146644 134714 146684
rect 134754 146644 134796 146684
rect 134836 146644 134878 146684
rect 134918 146644 134960 146684
rect 135000 146644 135009 146684
rect 149743 146644 149752 146684
rect 149792 146644 149834 146684
rect 149874 146644 149916 146684
rect 149956 146644 149998 146684
rect 150038 146644 150080 146684
rect 150120 146644 150129 146684
rect 75383 145888 75392 145928
rect 75432 145888 75474 145928
rect 75514 145888 75556 145928
rect 75596 145888 75638 145928
rect 75678 145888 75720 145928
rect 75760 145888 75769 145928
rect 90503 145888 90512 145928
rect 90552 145888 90594 145928
rect 90634 145888 90676 145928
rect 90716 145888 90758 145928
rect 90798 145888 90840 145928
rect 90880 145888 90889 145928
rect 105623 145888 105632 145928
rect 105672 145888 105714 145928
rect 105754 145888 105796 145928
rect 105836 145888 105878 145928
rect 105918 145888 105960 145928
rect 106000 145888 106009 145928
rect 120743 145888 120752 145928
rect 120792 145888 120834 145928
rect 120874 145888 120916 145928
rect 120956 145888 120998 145928
rect 121038 145888 121080 145928
rect 121120 145888 121129 145928
rect 135863 145888 135872 145928
rect 135912 145888 135954 145928
rect 135994 145888 136036 145928
rect 136076 145888 136118 145928
rect 136158 145888 136200 145928
rect 136240 145888 136249 145928
rect 150983 145888 150992 145928
rect 151032 145888 151074 145928
rect 151114 145888 151156 145928
rect 151196 145888 151238 145928
rect 151278 145888 151320 145928
rect 151360 145888 151369 145928
rect 74143 145132 74152 145172
rect 74192 145132 74234 145172
rect 74274 145132 74316 145172
rect 74356 145132 74398 145172
rect 74438 145132 74480 145172
rect 74520 145132 74529 145172
rect 89263 145132 89272 145172
rect 89312 145132 89354 145172
rect 89394 145132 89436 145172
rect 89476 145132 89518 145172
rect 89558 145132 89600 145172
rect 89640 145132 89649 145172
rect 104383 145132 104392 145172
rect 104432 145132 104474 145172
rect 104514 145132 104556 145172
rect 104596 145132 104638 145172
rect 104678 145132 104720 145172
rect 104760 145132 104769 145172
rect 119503 145132 119512 145172
rect 119552 145132 119594 145172
rect 119634 145132 119676 145172
rect 119716 145132 119758 145172
rect 119798 145132 119840 145172
rect 119880 145132 119889 145172
rect 134623 145132 134632 145172
rect 134672 145132 134714 145172
rect 134754 145132 134796 145172
rect 134836 145132 134878 145172
rect 134918 145132 134960 145172
rect 135000 145132 135009 145172
rect 149743 145132 149752 145172
rect 149792 145132 149834 145172
rect 149874 145132 149916 145172
rect 149956 145132 149998 145172
rect 150038 145132 150080 145172
rect 150120 145132 150129 145172
rect 75383 144376 75392 144416
rect 75432 144376 75474 144416
rect 75514 144376 75556 144416
rect 75596 144376 75638 144416
rect 75678 144376 75720 144416
rect 75760 144376 75769 144416
rect 90503 144376 90512 144416
rect 90552 144376 90594 144416
rect 90634 144376 90676 144416
rect 90716 144376 90758 144416
rect 90798 144376 90840 144416
rect 90880 144376 90889 144416
rect 105623 144376 105632 144416
rect 105672 144376 105714 144416
rect 105754 144376 105796 144416
rect 105836 144376 105878 144416
rect 105918 144376 105960 144416
rect 106000 144376 106009 144416
rect 120743 144376 120752 144416
rect 120792 144376 120834 144416
rect 120874 144376 120916 144416
rect 120956 144376 120998 144416
rect 121038 144376 121080 144416
rect 121120 144376 121129 144416
rect 135863 144376 135872 144416
rect 135912 144376 135954 144416
rect 135994 144376 136036 144416
rect 136076 144376 136118 144416
rect 136158 144376 136200 144416
rect 136240 144376 136249 144416
rect 150983 144376 150992 144416
rect 151032 144376 151074 144416
rect 151114 144376 151156 144416
rect 151196 144376 151238 144416
rect 151278 144376 151320 144416
rect 151360 144376 151369 144416
rect 74143 143620 74152 143660
rect 74192 143620 74234 143660
rect 74274 143620 74316 143660
rect 74356 143620 74398 143660
rect 74438 143620 74480 143660
rect 74520 143620 74529 143660
rect 89263 143620 89272 143660
rect 89312 143620 89354 143660
rect 89394 143620 89436 143660
rect 89476 143620 89518 143660
rect 89558 143620 89600 143660
rect 89640 143620 89649 143660
rect 104383 143620 104392 143660
rect 104432 143620 104474 143660
rect 104514 143620 104556 143660
rect 104596 143620 104638 143660
rect 104678 143620 104720 143660
rect 104760 143620 104769 143660
rect 119503 143620 119512 143660
rect 119552 143620 119594 143660
rect 119634 143620 119676 143660
rect 119716 143620 119758 143660
rect 119798 143620 119840 143660
rect 119880 143620 119889 143660
rect 134623 143620 134632 143660
rect 134672 143620 134714 143660
rect 134754 143620 134796 143660
rect 134836 143620 134878 143660
rect 134918 143620 134960 143660
rect 135000 143620 135009 143660
rect 149743 143620 149752 143660
rect 149792 143620 149834 143660
rect 149874 143620 149916 143660
rect 149956 143620 149998 143660
rect 150038 143620 150080 143660
rect 150120 143620 150129 143660
rect 75383 142864 75392 142904
rect 75432 142864 75474 142904
rect 75514 142864 75556 142904
rect 75596 142864 75638 142904
rect 75678 142864 75720 142904
rect 75760 142864 75769 142904
rect 90503 142864 90512 142904
rect 90552 142864 90594 142904
rect 90634 142864 90676 142904
rect 90716 142864 90758 142904
rect 90798 142864 90840 142904
rect 90880 142864 90889 142904
rect 105623 142864 105632 142904
rect 105672 142864 105714 142904
rect 105754 142864 105796 142904
rect 105836 142864 105878 142904
rect 105918 142864 105960 142904
rect 106000 142864 106009 142904
rect 120743 142864 120752 142904
rect 120792 142864 120834 142904
rect 120874 142864 120916 142904
rect 120956 142864 120998 142904
rect 121038 142864 121080 142904
rect 121120 142864 121129 142904
rect 135863 142864 135872 142904
rect 135912 142864 135954 142904
rect 135994 142864 136036 142904
rect 136076 142864 136118 142904
rect 136158 142864 136200 142904
rect 136240 142864 136249 142904
rect 150983 142864 150992 142904
rect 151032 142864 151074 142904
rect 151114 142864 151156 142904
rect 151196 142864 151238 142904
rect 151278 142864 151320 142904
rect 151360 142864 151369 142904
rect 74143 142108 74152 142148
rect 74192 142108 74234 142148
rect 74274 142108 74316 142148
rect 74356 142108 74398 142148
rect 74438 142108 74480 142148
rect 74520 142108 74529 142148
rect 89263 142108 89272 142148
rect 89312 142108 89354 142148
rect 89394 142108 89436 142148
rect 89476 142108 89518 142148
rect 89558 142108 89600 142148
rect 89640 142108 89649 142148
rect 104383 142108 104392 142148
rect 104432 142108 104474 142148
rect 104514 142108 104556 142148
rect 104596 142108 104638 142148
rect 104678 142108 104720 142148
rect 104760 142108 104769 142148
rect 119503 142108 119512 142148
rect 119552 142108 119594 142148
rect 119634 142108 119676 142148
rect 119716 142108 119758 142148
rect 119798 142108 119840 142148
rect 119880 142108 119889 142148
rect 134623 142108 134632 142148
rect 134672 142108 134714 142148
rect 134754 142108 134796 142148
rect 134836 142108 134878 142148
rect 134918 142108 134960 142148
rect 135000 142108 135009 142148
rect 149743 142108 149752 142148
rect 149792 142108 149834 142148
rect 149874 142108 149916 142148
rect 149956 142108 149998 142148
rect 150038 142108 150080 142148
rect 150120 142108 150129 142148
rect 75383 141352 75392 141392
rect 75432 141352 75474 141392
rect 75514 141352 75556 141392
rect 75596 141352 75638 141392
rect 75678 141352 75720 141392
rect 75760 141352 75769 141392
rect 90503 141352 90512 141392
rect 90552 141352 90594 141392
rect 90634 141352 90676 141392
rect 90716 141352 90758 141392
rect 90798 141352 90840 141392
rect 90880 141352 90889 141392
rect 105623 141352 105632 141392
rect 105672 141352 105714 141392
rect 105754 141352 105796 141392
rect 105836 141352 105878 141392
rect 105918 141352 105960 141392
rect 106000 141352 106009 141392
rect 120743 141352 120752 141392
rect 120792 141352 120834 141392
rect 120874 141352 120916 141392
rect 120956 141352 120998 141392
rect 121038 141352 121080 141392
rect 121120 141352 121129 141392
rect 135863 141352 135872 141392
rect 135912 141352 135954 141392
rect 135994 141352 136036 141392
rect 136076 141352 136118 141392
rect 136158 141352 136200 141392
rect 136240 141352 136249 141392
rect 150983 141352 150992 141392
rect 151032 141352 151074 141392
rect 151114 141352 151156 141392
rect 151196 141352 151238 141392
rect 151278 141352 151320 141392
rect 151360 141352 151369 141392
rect 74143 140596 74152 140636
rect 74192 140596 74234 140636
rect 74274 140596 74316 140636
rect 74356 140596 74398 140636
rect 74438 140596 74480 140636
rect 74520 140596 74529 140636
rect 89263 140596 89272 140636
rect 89312 140596 89354 140636
rect 89394 140596 89436 140636
rect 89476 140596 89518 140636
rect 89558 140596 89600 140636
rect 89640 140596 89649 140636
rect 104383 140596 104392 140636
rect 104432 140596 104474 140636
rect 104514 140596 104556 140636
rect 104596 140596 104638 140636
rect 104678 140596 104720 140636
rect 104760 140596 104769 140636
rect 119503 140596 119512 140636
rect 119552 140596 119594 140636
rect 119634 140596 119676 140636
rect 119716 140596 119758 140636
rect 119798 140596 119840 140636
rect 119880 140596 119889 140636
rect 134623 140596 134632 140636
rect 134672 140596 134714 140636
rect 134754 140596 134796 140636
rect 134836 140596 134878 140636
rect 134918 140596 134960 140636
rect 135000 140596 135009 140636
rect 149743 140596 149752 140636
rect 149792 140596 149834 140636
rect 149874 140596 149916 140636
rect 149956 140596 149998 140636
rect 150038 140596 150080 140636
rect 150120 140596 150129 140636
rect 75383 139840 75392 139880
rect 75432 139840 75474 139880
rect 75514 139840 75556 139880
rect 75596 139840 75638 139880
rect 75678 139840 75720 139880
rect 75760 139840 75769 139880
rect 90503 139840 90512 139880
rect 90552 139840 90594 139880
rect 90634 139840 90676 139880
rect 90716 139840 90758 139880
rect 90798 139840 90840 139880
rect 90880 139840 90889 139880
rect 105623 139840 105632 139880
rect 105672 139840 105714 139880
rect 105754 139840 105796 139880
rect 105836 139840 105878 139880
rect 105918 139840 105960 139880
rect 106000 139840 106009 139880
rect 120743 139840 120752 139880
rect 120792 139840 120834 139880
rect 120874 139840 120916 139880
rect 120956 139840 120998 139880
rect 121038 139840 121080 139880
rect 121120 139840 121129 139880
rect 135863 139840 135872 139880
rect 135912 139840 135954 139880
rect 135994 139840 136036 139880
rect 136076 139840 136118 139880
rect 136158 139840 136200 139880
rect 136240 139840 136249 139880
rect 150983 139840 150992 139880
rect 151032 139840 151074 139880
rect 151114 139840 151156 139880
rect 151196 139840 151238 139880
rect 151278 139840 151320 139880
rect 151360 139840 151369 139880
rect 74143 139084 74152 139124
rect 74192 139084 74234 139124
rect 74274 139084 74316 139124
rect 74356 139084 74398 139124
rect 74438 139084 74480 139124
rect 74520 139084 74529 139124
rect 89263 139084 89272 139124
rect 89312 139084 89354 139124
rect 89394 139084 89436 139124
rect 89476 139084 89518 139124
rect 89558 139084 89600 139124
rect 89640 139084 89649 139124
rect 104383 139084 104392 139124
rect 104432 139084 104474 139124
rect 104514 139084 104556 139124
rect 104596 139084 104638 139124
rect 104678 139084 104720 139124
rect 104760 139084 104769 139124
rect 119503 139084 119512 139124
rect 119552 139084 119594 139124
rect 119634 139084 119676 139124
rect 119716 139084 119758 139124
rect 119798 139084 119840 139124
rect 119880 139084 119889 139124
rect 134623 139084 134632 139124
rect 134672 139084 134714 139124
rect 134754 139084 134796 139124
rect 134836 139084 134878 139124
rect 134918 139084 134960 139124
rect 135000 139084 135009 139124
rect 149743 139084 149752 139124
rect 149792 139084 149834 139124
rect 149874 139084 149916 139124
rect 149956 139084 149998 139124
rect 150038 139084 150080 139124
rect 150120 139084 150129 139124
rect 75383 138328 75392 138368
rect 75432 138328 75474 138368
rect 75514 138328 75556 138368
rect 75596 138328 75638 138368
rect 75678 138328 75720 138368
rect 75760 138328 75769 138368
rect 90503 138328 90512 138368
rect 90552 138328 90594 138368
rect 90634 138328 90676 138368
rect 90716 138328 90758 138368
rect 90798 138328 90840 138368
rect 90880 138328 90889 138368
rect 105623 138328 105632 138368
rect 105672 138328 105714 138368
rect 105754 138328 105796 138368
rect 105836 138328 105878 138368
rect 105918 138328 105960 138368
rect 106000 138328 106009 138368
rect 120743 138328 120752 138368
rect 120792 138328 120834 138368
rect 120874 138328 120916 138368
rect 120956 138328 120998 138368
rect 121038 138328 121080 138368
rect 121120 138328 121129 138368
rect 135863 138328 135872 138368
rect 135912 138328 135954 138368
rect 135994 138328 136036 138368
rect 136076 138328 136118 138368
rect 136158 138328 136200 138368
rect 136240 138328 136249 138368
rect 150983 138328 150992 138368
rect 151032 138328 151074 138368
rect 151114 138328 151156 138368
rect 151196 138328 151238 138368
rect 151278 138328 151320 138368
rect 151360 138328 151369 138368
rect 74143 137572 74152 137612
rect 74192 137572 74234 137612
rect 74274 137572 74316 137612
rect 74356 137572 74398 137612
rect 74438 137572 74480 137612
rect 74520 137572 74529 137612
rect 89263 137572 89272 137612
rect 89312 137572 89354 137612
rect 89394 137572 89436 137612
rect 89476 137572 89518 137612
rect 89558 137572 89600 137612
rect 89640 137572 89649 137612
rect 104383 137572 104392 137612
rect 104432 137572 104474 137612
rect 104514 137572 104556 137612
rect 104596 137572 104638 137612
rect 104678 137572 104720 137612
rect 104760 137572 104769 137612
rect 119503 137572 119512 137612
rect 119552 137572 119594 137612
rect 119634 137572 119676 137612
rect 119716 137572 119758 137612
rect 119798 137572 119840 137612
rect 119880 137572 119889 137612
rect 134623 137572 134632 137612
rect 134672 137572 134714 137612
rect 134754 137572 134796 137612
rect 134836 137572 134878 137612
rect 134918 137572 134960 137612
rect 135000 137572 135009 137612
rect 149743 137572 149752 137612
rect 149792 137572 149834 137612
rect 149874 137572 149916 137612
rect 149956 137572 149998 137612
rect 150038 137572 150080 137612
rect 150120 137572 150129 137612
rect 75383 136816 75392 136856
rect 75432 136816 75474 136856
rect 75514 136816 75556 136856
rect 75596 136816 75638 136856
rect 75678 136816 75720 136856
rect 75760 136816 75769 136856
rect 90503 136816 90512 136856
rect 90552 136816 90594 136856
rect 90634 136816 90676 136856
rect 90716 136816 90758 136856
rect 90798 136816 90840 136856
rect 90880 136816 90889 136856
rect 105623 136816 105632 136856
rect 105672 136816 105714 136856
rect 105754 136816 105796 136856
rect 105836 136816 105878 136856
rect 105918 136816 105960 136856
rect 106000 136816 106009 136856
rect 120743 136816 120752 136856
rect 120792 136816 120834 136856
rect 120874 136816 120916 136856
rect 120956 136816 120998 136856
rect 121038 136816 121080 136856
rect 121120 136816 121129 136856
rect 135863 136816 135872 136856
rect 135912 136816 135954 136856
rect 135994 136816 136036 136856
rect 136076 136816 136118 136856
rect 136158 136816 136200 136856
rect 136240 136816 136249 136856
rect 150983 136816 150992 136856
rect 151032 136816 151074 136856
rect 151114 136816 151156 136856
rect 151196 136816 151238 136856
rect 151278 136816 151320 136856
rect 151360 136816 151369 136856
rect 74143 136060 74152 136100
rect 74192 136060 74234 136100
rect 74274 136060 74316 136100
rect 74356 136060 74398 136100
rect 74438 136060 74480 136100
rect 74520 136060 74529 136100
rect 89263 136060 89272 136100
rect 89312 136060 89354 136100
rect 89394 136060 89436 136100
rect 89476 136060 89518 136100
rect 89558 136060 89600 136100
rect 89640 136060 89649 136100
rect 104383 136060 104392 136100
rect 104432 136060 104474 136100
rect 104514 136060 104556 136100
rect 104596 136060 104638 136100
rect 104678 136060 104720 136100
rect 104760 136060 104769 136100
rect 119503 136060 119512 136100
rect 119552 136060 119594 136100
rect 119634 136060 119676 136100
rect 119716 136060 119758 136100
rect 119798 136060 119840 136100
rect 119880 136060 119889 136100
rect 134623 136060 134632 136100
rect 134672 136060 134714 136100
rect 134754 136060 134796 136100
rect 134836 136060 134878 136100
rect 134918 136060 134960 136100
rect 135000 136060 135009 136100
rect 149743 136060 149752 136100
rect 149792 136060 149834 136100
rect 149874 136060 149916 136100
rect 149956 136060 149998 136100
rect 150038 136060 150080 136100
rect 150120 136060 150129 136100
rect 64099 135976 64108 136016
rect 64148 135976 160032 136016
rect 75383 135304 75392 135344
rect 75432 135304 75474 135344
rect 75514 135304 75556 135344
rect 75596 135304 75638 135344
rect 75678 135304 75720 135344
rect 75760 135304 75769 135344
rect 90503 135304 90512 135344
rect 90552 135304 90594 135344
rect 90634 135304 90676 135344
rect 90716 135304 90758 135344
rect 90798 135304 90840 135344
rect 90880 135304 90889 135344
rect 105623 135304 105632 135344
rect 105672 135304 105714 135344
rect 105754 135304 105796 135344
rect 105836 135304 105878 135344
rect 105918 135304 105960 135344
rect 106000 135304 106009 135344
rect 120743 135304 120752 135344
rect 120792 135304 120834 135344
rect 120874 135304 120916 135344
rect 120956 135304 120998 135344
rect 121038 135304 121080 135344
rect 121120 135304 121129 135344
rect 135863 135304 135872 135344
rect 135912 135304 135954 135344
rect 135994 135304 136036 135344
rect 136076 135304 136118 135344
rect 136158 135304 136200 135344
rect 136240 135304 136249 135344
rect 150983 135304 150992 135344
rect 151032 135304 151074 135344
rect 151114 135304 151156 135344
rect 151196 135304 151238 135344
rect 151278 135304 151320 135344
rect 151360 135304 151369 135344
rect 74143 134548 74152 134588
rect 74192 134548 74234 134588
rect 74274 134548 74316 134588
rect 74356 134548 74398 134588
rect 74438 134548 74480 134588
rect 74520 134548 74529 134588
rect 89263 134548 89272 134588
rect 89312 134548 89354 134588
rect 89394 134548 89436 134588
rect 89476 134548 89518 134588
rect 89558 134548 89600 134588
rect 89640 134548 89649 134588
rect 104383 134548 104392 134588
rect 104432 134548 104474 134588
rect 104514 134548 104556 134588
rect 104596 134548 104638 134588
rect 104678 134548 104720 134588
rect 104760 134548 104769 134588
rect 119503 134548 119512 134588
rect 119552 134548 119594 134588
rect 119634 134548 119676 134588
rect 119716 134548 119758 134588
rect 119798 134548 119840 134588
rect 119880 134548 119889 134588
rect 134623 134548 134632 134588
rect 134672 134548 134714 134588
rect 134754 134548 134796 134588
rect 134836 134548 134878 134588
rect 134918 134548 134960 134588
rect 135000 134548 135009 134588
rect 149743 134548 149752 134588
rect 149792 134548 149834 134588
rect 149874 134548 149916 134588
rect 149956 134548 149998 134588
rect 150038 134548 150080 134588
rect 150120 134548 150129 134588
rect 75383 133792 75392 133832
rect 75432 133792 75474 133832
rect 75514 133792 75556 133832
rect 75596 133792 75638 133832
rect 75678 133792 75720 133832
rect 75760 133792 75769 133832
rect 90503 133792 90512 133832
rect 90552 133792 90594 133832
rect 90634 133792 90676 133832
rect 90716 133792 90758 133832
rect 90798 133792 90840 133832
rect 90880 133792 90889 133832
rect 105623 133792 105632 133832
rect 105672 133792 105714 133832
rect 105754 133792 105796 133832
rect 105836 133792 105878 133832
rect 105918 133792 105960 133832
rect 106000 133792 106009 133832
rect 120743 133792 120752 133832
rect 120792 133792 120834 133832
rect 120874 133792 120916 133832
rect 120956 133792 120998 133832
rect 121038 133792 121080 133832
rect 121120 133792 121129 133832
rect 135863 133792 135872 133832
rect 135912 133792 135954 133832
rect 135994 133792 136036 133832
rect 136076 133792 136118 133832
rect 136158 133792 136200 133832
rect 136240 133792 136249 133832
rect 150983 133792 150992 133832
rect 151032 133792 151074 133832
rect 151114 133792 151156 133832
rect 151196 133792 151238 133832
rect 151278 133792 151320 133832
rect 151360 133792 151369 133832
rect 74143 133036 74152 133076
rect 74192 133036 74234 133076
rect 74274 133036 74316 133076
rect 74356 133036 74398 133076
rect 74438 133036 74480 133076
rect 74520 133036 74529 133076
rect 89263 133036 89272 133076
rect 89312 133036 89354 133076
rect 89394 133036 89436 133076
rect 89476 133036 89518 133076
rect 89558 133036 89600 133076
rect 89640 133036 89649 133076
rect 104383 133036 104392 133076
rect 104432 133036 104474 133076
rect 104514 133036 104556 133076
rect 104596 133036 104638 133076
rect 104678 133036 104720 133076
rect 104760 133036 104769 133076
rect 119503 133036 119512 133076
rect 119552 133036 119594 133076
rect 119634 133036 119676 133076
rect 119716 133036 119758 133076
rect 119798 133036 119840 133076
rect 119880 133036 119889 133076
rect 134623 133036 134632 133076
rect 134672 133036 134714 133076
rect 134754 133036 134796 133076
rect 134836 133036 134878 133076
rect 134918 133036 134960 133076
rect 135000 133036 135009 133076
rect 149743 133036 149752 133076
rect 149792 133036 149834 133076
rect 149874 133036 149916 133076
rect 149956 133036 149998 133076
rect 150038 133036 150080 133076
rect 150120 133036 150129 133076
rect 75383 132280 75392 132320
rect 75432 132280 75474 132320
rect 75514 132280 75556 132320
rect 75596 132280 75638 132320
rect 75678 132280 75720 132320
rect 75760 132280 75769 132320
rect 90503 132280 90512 132320
rect 90552 132280 90594 132320
rect 90634 132280 90676 132320
rect 90716 132280 90758 132320
rect 90798 132280 90840 132320
rect 90880 132280 90889 132320
rect 105623 132280 105632 132320
rect 105672 132280 105714 132320
rect 105754 132280 105796 132320
rect 105836 132280 105878 132320
rect 105918 132280 105960 132320
rect 106000 132280 106009 132320
rect 120743 132280 120752 132320
rect 120792 132280 120834 132320
rect 120874 132280 120916 132320
rect 120956 132280 120998 132320
rect 121038 132280 121080 132320
rect 121120 132280 121129 132320
rect 135863 132280 135872 132320
rect 135912 132280 135954 132320
rect 135994 132280 136036 132320
rect 136076 132280 136118 132320
rect 136158 132280 136200 132320
rect 136240 132280 136249 132320
rect 150983 132280 150992 132320
rect 151032 132280 151074 132320
rect 151114 132280 151156 132320
rect 151196 132280 151238 132320
rect 151278 132280 151320 132320
rect 151360 132280 151369 132320
rect 74143 131524 74152 131564
rect 74192 131524 74234 131564
rect 74274 131524 74316 131564
rect 74356 131524 74398 131564
rect 74438 131524 74480 131564
rect 74520 131524 74529 131564
rect 89263 131524 89272 131564
rect 89312 131524 89354 131564
rect 89394 131524 89436 131564
rect 89476 131524 89518 131564
rect 89558 131524 89600 131564
rect 89640 131524 89649 131564
rect 104383 131524 104392 131564
rect 104432 131524 104474 131564
rect 104514 131524 104556 131564
rect 104596 131524 104638 131564
rect 104678 131524 104720 131564
rect 104760 131524 104769 131564
rect 119503 131524 119512 131564
rect 119552 131524 119594 131564
rect 119634 131524 119676 131564
rect 119716 131524 119758 131564
rect 119798 131524 119840 131564
rect 119880 131524 119889 131564
rect 134623 131524 134632 131564
rect 134672 131524 134714 131564
rect 134754 131524 134796 131564
rect 134836 131524 134878 131564
rect 134918 131524 134960 131564
rect 135000 131524 135009 131564
rect 149743 131524 149752 131564
rect 149792 131524 149834 131564
rect 149874 131524 149916 131564
rect 149956 131524 149998 131564
rect 150038 131524 150080 131564
rect 150120 131524 150129 131564
rect 75383 130768 75392 130808
rect 75432 130768 75474 130808
rect 75514 130768 75556 130808
rect 75596 130768 75638 130808
rect 75678 130768 75720 130808
rect 75760 130768 75769 130808
rect 90503 130768 90512 130808
rect 90552 130768 90594 130808
rect 90634 130768 90676 130808
rect 90716 130768 90758 130808
rect 90798 130768 90840 130808
rect 90880 130768 90889 130808
rect 105623 130768 105632 130808
rect 105672 130768 105714 130808
rect 105754 130768 105796 130808
rect 105836 130768 105878 130808
rect 105918 130768 105960 130808
rect 106000 130768 106009 130808
rect 120743 130768 120752 130808
rect 120792 130768 120834 130808
rect 120874 130768 120916 130808
rect 120956 130768 120998 130808
rect 121038 130768 121080 130808
rect 121120 130768 121129 130808
rect 135863 130768 135872 130808
rect 135912 130768 135954 130808
rect 135994 130768 136036 130808
rect 136076 130768 136118 130808
rect 136158 130768 136200 130808
rect 136240 130768 136249 130808
rect 150983 130768 150992 130808
rect 151032 130768 151074 130808
rect 151114 130768 151156 130808
rect 151196 130768 151238 130808
rect 151278 130768 151320 130808
rect 151360 130768 151369 130808
rect 74143 130012 74152 130052
rect 74192 130012 74234 130052
rect 74274 130012 74316 130052
rect 74356 130012 74398 130052
rect 74438 130012 74480 130052
rect 74520 130012 74529 130052
rect 89263 130012 89272 130052
rect 89312 130012 89354 130052
rect 89394 130012 89436 130052
rect 89476 130012 89518 130052
rect 89558 130012 89600 130052
rect 89640 130012 89649 130052
rect 104383 130012 104392 130052
rect 104432 130012 104474 130052
rect 104514 130012 104556 130052
rect 104596 130012 104638 130052
rect 104678 130012 104720 130052
rect 104760 130012 104769 130052
rect 119503 130012 119512 130052
rect 119552 130012 119594 130052
rect 119634 130012 119676 130052
rect 119716 130012 119758 130052
rect 119798 130012 119840 130052
rect 119880 130012 119889 130052
rect 134623 130012 134632 130052
rect 134672 130012 134714 130052
rect 134754 130012 134796 130052
rect 134836 130012 134878 130052
rect 134918 130012 134960 130052
rect 135000 130012 135009 130052
rect 149743 130012 149752 130052
rect 149792 130012 149834 130052
rect 149874 130012 149916 130052
rect 149956 130012 149998 130052
rect 150038 130012 150080 130052
rect 150120 130012 150129 130052
rect 75383 129256 75392 129296
rect 75432 129256 75474 129296
rect 75514 129256 75556 129296
rect 75596 129256 75638 129296
rect 75678 129256 75720 129296
rect 75760 129256 75769 129296
rect 90503 129256 90512 129296
rect 90552 129256 90594 129296
rect 90634 129256 90676 129296
rect 90716 129256 90758 129296
rect 90798 129256 90840 129296
rect 90880 129256 90889 129296
rect 105623 129256 105632 129296
rect 105672 129256 105714 129296
rect 105754 129256 105796 129296
rect 105836 129256 105878 129296
rect 105918 129256 105960 129296
rect 106000 129256 106009 129296
rect 120743 129256 120752 129296
rect 120792 129256 120834 129296
rect 120874 129256 120916 129296
rect 120956 129256 120998 129296
rect 121038 129256 121080 129296
rect 121120 129256 121129 129296
rect 135863 129256 135872 129296
rect 135912 129256 135954 129296
rect 135994 129256 136036 129296
rect 136076 129256 136118 129296
rect 136158 129256 136200 129296
rect 136240 129256 136249 129296
rect 150983 129256 150992 129296
rect 151032 129256 151074 129296
rect 151114 129256 151156 129296
rect 151196 129256 151238 129296
rect 151278 129256 151320 129296
rect 151360 129256 151369 129296
rect 74143 128500 74152 128540
rect 74192 128500 74234 128540
rect 74274 128500 74316 128540
rect 74356 128500 74398 128540
rect 74438 128500 74480 128540
rect 74520 128500 74529 128540
rect 89263 128500 89272 128540
rect 89312 128500 89354 128540
rect 89394 128500 89436 128540
rect 89476 128500 89518 128540
rect 89558 128500 89600 128540
rect 89640 128500 89649 128540
rect 104383 128500 104392 128540
rect 104432 128500 104474 128540
rect 104514 128500 104556 128540
rect 104596 128500 104638 128540
rect 104678 128500 104720 128540
rect 104760 128500 104769 128540
rect 119503 128500 119512 128540
rect 119552 128500 119594 128540
rect 119634 128500 119676 128540
rect 119716 128500 119758 128540
rect 119798 128500 119840 128540
rect 119880 128500 119889 128540
rect 134623 128500 134632 128540
rect 134672 128500 134714 128540
rect 134754 128500 134796 128540
rect 134836 128500 134878 128540
rect 134918 128500 134960 128540
rect 135000 128500 135009 128540
rect 149743 128500 149752 128540
rect 149792 128500 149834 128540
rect 149874 128500 149916 128540
rect 149956 128500 149998 128540
rect 150038 128500 150080 128540
rect 150120 128500 150129 128540
rect 75383 127744 75392 127784
rect 75432 127744 75474 127784
rect 75514 127744 75556 127784
rect 75596 127744 75638 127784
rect 75678 127744 75720 127784
rect 75760 127744 75769 127784
rect 90503 127744 90512 127784
rect 90552 127744 90594 127784
rect 90634 127744 90676 127784
rect 90716 127744 90758 127784
rect 90798 127744 90840 127784
rect 90880 127744 90889 127784
rect 105623 127744 105632 127784
rect 105672 127744 105714 127784
rect 105754 127744 105796 127784
rect 105836 127744 105878 127784
rect 105918 127744 105960 127784
rect 106000 127744 106009 127784
rect 120743 127744 120752 127784
rect 120792 127744 120834 127784
rect 120874 127744 120916 127784
rect 120956 127744 120998 127784
rect 121038 127744 121080 127784
rect 121120 127744 121129 127784
rect 135863 127744 135872 127784
rect 135912 127744 135954 127784
rect 135994 127744 136036 127784
rect 136076 127744 136118 127784
rect 136158 127744 136200 127784
rect 136240 127744 136249 127784
rect 150983 127744 150992 127784
rect 151032 127744 151074 127784
rect 151114 127744 151156 127784
rect 151196 127744 151238 127784
rect 151278 127744 151320 127784
rect 151360 127744 151369 127784
rect 74143 126988 74152 127028
rect 74192 126988 74234 127028
rect 74274 126988 74316 127028
rect 74356 126988 74398 127028
rect 74438 126988 74480 127028
rect 74520 126988 74529 127028
rect 89263 126988 89272 127028
rect 89312 126988 89354 127028
rect 89394 126988 89436 127028
rect 89476 126988 89518 127028
rect 89558 126988 89600 127028
rect 89640 126988 89649 127028
rect 104383 126988 104392 127028
rect 104432 126988 104474 127028
rect 104514 126988 104556 127028
rect 104596 126988 104638 127028
rect 104678 126988 104720 127028
rect 104760 126988 104769 127028
rect 119503 126988 119512 127028
rect 119552 126988 119594 127028
rect 119634 126988 119676 127028
rect 119716 126988 119758 127028
rect 119798 126988 119840 127028
rect 119880 126988 119889 127028
rect 134623 126988 134632 127028
rect 134672 126988 134714 127028
rect 134754 126988 134796 127028
rect 134836 126988 134878 127028
rect 134918 126988 134960 127028
rect 135000 126988 135009 127028
rect 149743 126988 149752 127028
rect 149792 126988 149834 127028
rect 149874 126988 149916 127028
rect 149956 126988 149998 127028
rect 150038 126988 150080 127028
rect 150120 126988 150129 127028
rect 75383 126232 75392 126272
rect 75432 126232 75474 126272
rect 75514 126232 75556 126272
rect 75596 126232 75638 126272
rect 75678 126232 75720 126272
rect 75760 126232 75769 126272
rect 90503 126232 90512 126272
rect 90552 126232 90594 126272
rect 90634 126232 90676 126272
rect 90716 126232 90758 126272
rect 90798 126232 90840 126272
rect 90880 126232 90889 126272
rect 105623 126232 105632 126272
rect 105672 126232 105714 126272
rect 105754 126232 105796 126272
rect 105836 126232 105878 126272
rect 105918 126232 105960 126272
rect 106000 126232 106009 126272
rect 120743 126232 120752 126272
rect 120792 126232 120834 126272
rect 120874 126232 120916 126272
rect 120956 126232 120998 126272
rect 121038 126232 121080 126272
rect 121120 126232 121129 126272
rect 135863 126232 135872 126272
rect 135912 126232 135954 126272
rect 135994 126232 136036 126272
rect 136076 126232 136118 126272
rect 136158 126232 136200 126272
rect 136240 126232 136249 126272
rect 150983 126232 150992 126272
rect 151032 126232 151074 126272
rect 151114 126232 151156 126272
rect 151196 126232 151238 126272
rect 151278 126232 151320 126272
rect 151360 126232 151369 126272
rect 74143 125476 74152 125516
rect 74192 125476 74234 125516
rect 74274 125476 74316 125516
rect 74356 125476 74398 125516
rect 74438 125476 74480 125516
rect 74520 125476 74529 125516
rect 89263 125476 89272 125516
rect 89312 125476 89354 125516
rect 89394 125476 89436 125516
rect 89476 125476 89518 125516
rect 89558 125476 89600 125516
rect 89640 125476 89649 125516
rect 104383 125476 104392 125516
rect 104432 125476 104474 125516
rect 104514 125476 104556 125516
rect 104596 125476 104638 125516
rect 104678 125476 104720 125516
rect 104760 125476 104769 125516
rect 119503 125476 119512 125516
rect 119552 125476 119594 125516
rect 119634 125476 119676 125516
rect 119716 125476 119758 125516
rect 119798 125476 119840 125516
rect 119880 125476 119889 125516
rect 134623 125476 134632 125516
rect 134672 125476 134714 125516
rect 134754 125476 134796 125516
rect 134836 125476 134878 125516
rect 134918 125476 134960 125516
rect 135000 125476 135009 125516
rect 149743 125476 149752 125516
rect 149792 125476 149834 125516
rect 149874 125476 149916 125516
rect 149956 125476 149998 125516
rect 150038 125476 150080 125516
rect 150120 125476 150129 125516
rect 75383 124720 75392 124760
rect 75432 124720 75474 124760
rect 75514 124720 75556 124760
rect 75596 124720 75638 124760
rect 75678 124720 75720 124760
rect 75760 124720 75769 124760
rect 90503 124720 90512 124760
rect 90552 124720 90594 124760
rect 90634 124720 90676 124760
rect 90716 124720 90758 124760
rect 90798 124720 90840 124760
rect 90880 124720 90889 124760
rect 105623 124720 105632 124760
rect 105672 124720 105714 124760
rect 105754 124720 105796 124760
rect 105836 124720 105878 124760
rect 105918 124720 105960 124760
rect 106000 124720 106009 124760
rect 120743 124720 120752 124760
rect 120792 124720 120834 124760
rect 120874 124720 120916 124760
rect 120956 124720 120998 124760
rect 121038 124720 121080 124760
rect 121120 124720 121129 124760
rect 135863 124720 135872 124760
rect 135912 124720 135954 124760
rect 135994 124720 136036 124760
rect 136076 124720 136118 124760
rect 136158 124720 136200 124760
rect 136240 124720 136249 124760
rect 150983 124720 150992 124760
rect 151032 124720 151074 124760
rect 151114 124720 151156 124760
rect 151196 124720 151238 124760
rect 151278 124720 151320 124760
rect 151360 124720 151369 124760
rect 74143 123964 74152 124004
rect 74192 123964 74234 124004
rect 74274 123964 74316 124004
rect 74356 123964 74398 124004
rect 74438 123964 74480 124004
rect 74520 123964 74529 124004
rect 89263 123964 89272 124004
rect 89312 123964 89354 124004
rect 89394 123964 89436 124004
rect 89476 123964 89518 124004
rect 89558 123964 89600 124004
rect 89640 123964 89649 124004
rect 104383 123964 104392 124004
rect 104432 123964 104474 124004
rect 104514 123964 104556 124004
rect 104596 123964 104638 124004
rect 104678 123964 104720 124004
rect 104760 123964 104769 124004
rect 119503 123964 119512 124004
rect 119552 123964 119594 124004
rect 119634 123964 119676 124004
rect 119716 123964 119758 124004
rect 119798 123964 119840 124004
rect 119880 123964 119889 124004
rect 134623 123964 134632 124004
rect 134672 123964 134714 124004
rect 134754 123964 134796 124004
rect 134836 123964 134878 124004
rect 134918 123964 134960 124004
rect 135000 123964 135009 124004
rect 149743 123964 149752 124004
rect 149792 123964 149834 124004
rect 149874 123964 149916 124004
rect 149956 123964 149998 124004
rect 150038 123964 150080 124004
rect 150120 123964 150129 124004
rect 75383 123208 75392 123248
rect 75432 123208 75474 123248
rect 75514 123208 75556 123248
rect 75596 123208 75638 123248
rect 75678 123208 75720 123248
rect 75760 123208 75769 123248
rect 90503 123208 90512 123248
rect 90552 123208 90594 123248
rect 90634 123208 90676 123248
rect 90716 123208 90758 123248
rect 90798 123208 90840 123248
rect 90880 123208 90889 123248
rect 105623 123208 105632 123248
rect 105672 123208 105714 123248
rect 105754 123208 105796 123248
rect 105836 123208 105878 123248
rect 105918 123208 105960 123248
rect 106000 123208 106009 123248
rect 120743 123208 120752 123248
rect 120792 123208 120834 123248
rect 120874 123208 120916 123248
rect 120956 123208 120998 123248
rect 121038 123208 121080 123248
rect 121120 123208 121129 123248
rect 135863 123208 135872 123248
rect 135912 123208 135954 123248
rect 135994 123208 136036 123248
rect 136076 123208 136118 123248
rect 136158 123208 136200 123248
rect 136240 123208 136249 123248
rect 150983 123208 150992 123248
rect 151032 123208 151074 123248
rect 151114 123208 151156 123248
rect 151196 123208 151238 123248
rect 151278 123208 151320 123248
rect 151360 123208 151369 123248
rect 74143 122452 74152 122492
rect 74192 122452 74234 122492
rect 74274 122452 74316 122492
rect 74356 122452 74398 122492
rect 74438 122452 74480 122492
rect 74520 122452 74529 122492
rect 89263 122452 89272 122492
rect 89312 122452 89354 122492
rect 89394 122452 89436 122492
rect 89476 122452 89518 122492
rect 89558 122452 89600 122492
rect 89640 122452 89649 122492
rect 104383 122452 104392 122492
rect 104432 122452 104474 122492
rect 104514 122452 104556 122492
rect 104596 122452 104638 122492
rect 104678 122452 104720 122492
rect 104760 122452 104769 122492
rect 119503 122452 119512 122492
rect 119552 122452 119594 122492
rect 119634 122452 119676 122492
rect 119716 122452 119758 122492
rect 119798 122452 119840 122492
rect 119880 122452 119889 122492
rect 134623 122452 134632 122492
rect 134672 122452 134714 122492
rect 134754 122452 134796 122492
rect 134836 122452 134878 122492
rect 134918 122452 134960 122492
rect 135000 122452 135009 122492
rect 149743 122452 149752 122492
rect 149792 122452 149834 122492
rect 149874 122452 149916 122492
rect 149956 122452 149998 122492
rect 150038 122452 150080 122492
rect 150120 122452 150129 122492
rect 75383 121696 75392 121736
rect 75432 121696 75474 121736
rect 75514 121696 75556 121736
rect 75596 121696 75638 121736
rect 75678 121696 75720 121736
rect 75760 121696 75769 121736
rect 90503 121696 90512 121736
rect 90552 121696 90594 121736
rect 90634 121696 90676 121736
rect 90716 121696 90758 121736
rect 90798 121696 90840 121736
rect 90880 121696 90889 121736
rect 105623 121696 105632 121736
rect 105672 121696 105714 121736
rect 105754 121696 105796 121736
rect 105836 121696 105878 121736
rect 105918 121696 105960 121736
rect 106000 121696 106009 121736
rect 120743 121696 120752 121736
rect 120792 121696 120834 121736
rect 120874 121696 120916 121736
rect 120956 121696 120998 121736
rect 121038 121696 121080 121736
rect 121120 121696 121129 121736
rect 135863 121696 135872 121736
rect 135912 121696 135954 121736
rect 135994 121696 136036 121736
rect 136076 121696 136118 121736
rect 136158 121696 136200 121736
rect 136240 121696 136249 121736
rect 150983 121696 150992 121736
rect 151032 121696 151074 121736
rect 151114 121696 151156 121736
rect 151196 121696 151238 121736
rect 151278 121696 151320 121736
rect 151360 121696 151369 121736
rect 74143 120940 74152 120980
rect 74192 120940 74234 120980
rect 74274 120940 74316 120980
rect 74356 120940 74398 120980
rect 74438 120940 74480 120980
rect 74520 120940 74529 120980
rect 89263 120940 89272 120980
rect 89312 120940 89354 120980
rect 89394 120940 89436 120980
rect 89476 120940 89518 120980
rect 89558 120940 89600 120980
rect 89640 120940 89649 120980
rect 104383 120940 104392 120980
rect 104432 120940 104474 120980
rect 104514 120940 104556 120980
rect 104596 120940 104638 120980
rect 104678 120940 104720 120980
rect 104760 120940 104769 120980
rect 119503 120940 119512 120980
rect 119552 120940 119594 120980
rect 119634 120940 119676 120980
rect 119716 120940 119758 120980
rect 119798 120940 119840 120980
rect 119880 120940 119889 120980
rect 134623 120940 134632 120980
rect 134672 120940 134714 120980
rect 134754 120940 134796 120980
rect 134836 120940 134878 120980
rect 134918 120940 134960 120980
rect 135000 120940 135009 120980
rect 149743 120940 149752 120980
rect 149792 120940 149834 120980
rect 149874 120940 149916 120980
rect 149956 120940 149998 120980
rect 150038 120940 150080 120980
rect 150120 120940 150129 120980
rect 75383 120184 75392 120224
rect 75432 120184 75474 120224
rect 75514 120184 75556 120224
rect 75596 120184 75638 120224
rect 75678 120184 75720 120224
rect 75760 120184 75769 120224
rect 90503 120184 90512 120224
rect 90552 120184 90594 120224
rect 90634 120184 90676 120224
rect 90716 120184 90758 120224
rect 90798 120184 90840 120224
rect 90880 120184 90889 120224
rect 105623 120184 105632 120224
rect 105672 120184 105714 120224
rect 105754 120184 105796 120224
rect 105836 120184 105878 120224
rect 105918 120184 105960 120224
rect 106000 120184 106009 120224
rect 120743 120184 120752 120224
rect 120792 120184 120834 120224
rect 120874 120184 120916 120224
rect 120956 120184 120998 120224
rect 121038 120184 121080 120224
rect 121120 120184 121129 120224
rect 135863 120184 135872 120224
rect 135912 120184 135954 120224
rect 135994 120184 136036 120224
rect 136076 120184 136118 120224
rect 136158 120184 136200 120224
rect 136240 120184 136249 120224
rect 150983 120184 150992 120224
rect 151032 120184 151074 120224
rect 151114 120184 151156 120224
rect 151196 120184 151238 120224
rect 151278 120184 151320 120224
rect 151360 120184 151369 120224
rect 64099 120016 64108 120056
rect 64148 120016 160032 120056
rect 74143 119428 74152 119468
rect 74192 119428 74234 119468
rect 74274 119428 74316 119468
rect 74356 119428 74398 119468
rect 74438 119428 74480 119468
rect 74520 119428 74529 119468
rect 89263 119428 89272 119468
rect 89312 119428 89354 119468
rect 89394 119428 89436 119468
rect 89476 119428 89518 119468
rect 89558 119428 89600 119468
rect 89640 119428 89649 119468
rect 104383 119428 104392 119468
rect 104432 119428 104474 119468
rect 104514 119428 104556 119468
rect 104596 119428 104638 119468
rect 104678 119428 104720 119468
rect 104760 119428 104769 119468
rect 119503 119428 119512 119468
rect 119552 119428 119594 119468
rect 119634 119428 119676 119468
rect 119716 119428 119758 119468
rect 119798 119428 119840 119468
rect 119880 119428 119889 119468
rect 134623 119428 134632 119468
rect 134672 119428 134714 119468
rect 134754 119428 134796 119468
rect 134836 119428 134878 119468
rect 134918 119428 134960 119468
rect 135000 119428 135009 119468
rect 149743 119428 149752 119468
rect 149792 119428 149834 119468
rect 149874 119428 149916 119468
rect 149956 119428 149998 119468
rect 150038 119428 150080 119468
rect 150120 119428 150129 119468
rect 75383 118672 75392 118712
rect 75432 118672 75474 118712
rect 75514 118672 75556 118712
rect 75596 118672 75638 118712
rect 75678 118672 75720 118712
rect 75760 118672 75769 118712
rect 90503 118672 90512 118712
rect 90552 118672 90594 118712
rect 90634 118672 90676 118712
rect 90716 118672 90758 118712
rect 90798 118672 90840 118712
rect 90880 118672 90889 118712
rect 105623 118672 105632 118712
rect 105672 118672 105714 118712
rect 105754 118672 105796 118712
rect 105836 118672 105878 118712
rect 105918 118672 105960 118712
rect 106000 118672 106009 118712
rect 120743 118672 120752 118712
rect 120792 118672 120834 118712
rect 120874 118672 120916 118712
rect 120956 118672 120998 118712
rect 121038 118672 121080 118712
rect 121120 118672 121129 118712
rect 135863 118672 135872 118712
rect 135912 118672 135954 118712
rect 135994 118672 136036 118712
rect 136076 118672 136118 118712
rect 136158 118672 136200 118712
rect 136240 118672 136249 118712
rect 150983 118672 150992 118712
rect 151032 118672 151074 118712
rect 151114 118672 151156 118712
rect 151196 118672 151238 118712
rect 151278 118672 151320 118712
rect 151360 118672 151369 118712
rect 74143 117916 74152 117956
rect 74192 117916 74234 117956
rect 74274 117916 74316 117956
rect 74356 117916 74398 117956
rect 74438 117916 74480 117956
rect 74520 117916 74529 117956
rect 89263 117916 89272 117956
rect 89312 117916 89354 117956
rect 89394 117916 89436 117956
rect 89476 117916 89518 117956
rect 89558 117916 89600 117956
rect 89640 117916 89649 117956
rect 104383 117916 104392 117956
rect 104432 117916 104474 117956
rect 104514 117916 104556 117956
rect 104596 117916 104638 117956
rect 104678 117916 104720 117956
rect 104760 117916 104769 117956
rect 119503 117916 119512 117956
rect 119552 117916 119594 117956
rect 119634 117916 119676 117956
rect 119716 117916 119758 117956
rect 119798 117916 119840 117956
rect 119880 117916 119889 117956
rect 134623 117916 134632 117956
rect 134672 117916 134714 117956
rect 134754 117916 134796 117956
rect 134836 117916 134878 117956
rect 134918 117916 134960 117956
rect 135000 117916 135009 117956
rect 149743 117916 149752 117956
rect 149792 117916 149834 117956
rect 149874 117916 149916 117956
rect 149956 117916 149998 117956
rect 150038 117916 150080 117956
rect 150120 117916 150129 117956
rect 75383 117160 75392 117200
rect 75432 117160 75474 117200
rect 75514 117160 75556 117200
rect 75596 117160 75638 117200
rect 75678 117160 75720 117200
rect 75760 117160 75769 117200
rect 90503 117160 90512 117200
rect 90552 117160 90594 117200
rect 90634 117160 90676 117200
rect 90716 117160 90758 117200
rect 90798 117160 90840 117200
rect 90880 117160 90889 117200
rect 105623 117160 105632 117200
rect 105672 117160 105714 117200
rect 105754 117160 105796 117200
rect 105836 117160 105878 117200
rect 105918 117160 105960 117200
rect 106000 117160 106009 117200
rect 120743 117160 120752 117200
rect 120792 117160 120834 117200
rect 120874 117160 120916 117200
rect 120956 117160 120998 117200
rect 121038 117160 121080 117200
rect 121120 117160 121129 117200
rect 135863 117160 135872 117200
rect 135912 117160 135954 117200
rect 135994 117160 136036 117200
rect 136076 117160 136118 117200
rect 136158 117160 136200 117200
rect 136240 117160 136249 117200
rect 150983 117160 150992 117200
rect 151032 117160 151074 117200
rect 151114 117160 151156 117200
rect 151196 117160 151238 117200
rect 151278 117160 151320 117200
rect 151360 117160 151369 117200
rect 74143 116404 74152 116444
rect 74192 116404 74234 116444
rect 74274 116404 74316 116444
rect 74356 116404 74398 116444
rect 74438 116404 74480 116444
rect 74520 116404 74529 116444
rect 89263 116404 89272 116444
rect 89312 116404 89354 116444
rect 89394 116404 89436 116444
rect 89476 116404 89518 116444
rect 89558 116404 89600 116444
rect 89640 116404 89649 116444
rect 104383 116404 104392 116444
rect 104432 116404 104474 116444
rect 104514 116404 104556 116444
rect 104596 116404 104638 116444
rect 104678 116404 104720 116444
rect 104760 116404 104769 116444
rect 119503 116404 119512 116444
rect 119552 116404 119594 116444
rect 119634 116404 119676 116444
rect 119716 116404 119758 116444
rect 119798 116404 119840 116444
rect 119880 116404 119889 116444
rect 134623 116404 134632 116444
rect 134672 116404 134714 116444
rect 134754 116404 134796 116444
rect 134836 116404 134878 116444
rect 134918 116404 134960 116444
rect 135000 116404 135009 116444
rect 149743 116404 149752 116444
rect 149792 116404 149834 116444
rect 149874 116404 149916 116444
rect 149956 116404 149998 116444
rect 150038 116404 150080 116444
rect 150120 116404 150129 116444
rect 75383 115648 75392 115688
rect 75432 115648 75474 115688
rect 75514 115648 75556 115688
rect 75596 115648 75638 115688
rect 75678 115648 75720 115688
rect 75760 115648 75769 115688
rect 90503 115648 90512 115688
rect 90552 115648 90594 115688
rect 90634 115648 90676 115688
rect 90716 115648 90758 115688
rect 90798 115648 90840 115688
rect 90880 115648 90889 115688
rect 105623 115648 105632 115688
rect 105672 115648 105714 115688
rect 105754 115648 105796 115688
rect 105836 115648 105878 115688
rect 105918 115648 105960 115688
rect 106000 115648 106009 115688
rect 120743 115648 120752 115688
rect 120792 115648 120834 115688
rect 120874 115648 120916 115688
rect 120956 115648 120998 115688
rect 121038 115648 121080 115688
rect 121120 115648 121129 115688
rect 135863 115648 135872 115688
rect 135912 115648 135954 115688
rect 135994 115648 136036 115688
rect 136076 115648 136118 115688
rect 136158 115648 136200 115688
rect 136240 115648 136249 115688
rect 150983 115648 150992 115688
rect 151032 115648 151074 115688
rect 151114 115648 151156 115688
rect 151196 115648 151238 115688
rect 151278 115648 151320 115688
rect 151360 115648 151369 115688
rect 74143 114892 74152 114932
rect 74192 114892 74234 114932
rect 74274 114892 74316 114932
rect 74356 114892 74398 114932
rect 74438 114892 74480 114932
rect 74520 114892 74529 114932
rect 89263 114892 89272 114932
rect 89312 114892 89354 114932
rect 89394 114892 89436 114932
rect 89476 114892 89518 114932
rect 89558 114892 89600 114932
rect 89640 114892 89649 114932
rect 104383 114892 104392 114932
rect 104432 114892 104474 114932
rect 104514 114892 104556 114932
rect 104596 114892 104638 114932
rect 104678 114892 104720 114932
rect 104760 114892 104769 114932
rect 119503 114892 119512 114932
rect 119552 114892 119594 114932
rect 119634 114892 119676 114932
rect 119716 114892 119758 114932
rect 119798 114892 119840 114932
rect 119880 114892 119889 114932
rect 134623 114892 134632 114932
rect 134672 114892 134714 114932
rect 134754 114892 134796 114932
rect 134836 114892 134878 114932
rect 134918 114892 134960 114932
rect 135000 114892 135009 114932
rect 149743 114892 149752 114932
rect 149792 114892 149834 114932
rect 149874 114892 149916 114932
rect 149956 114892 149998 114932
rect 150038 114892 150080 114932
rect 150120 114892 150129 114932
rect 75383 114136 75392 114176
rect 75432 114136 75474 114176
rect 75514 114136 75556 114176
rect 75596 114136 75638 114176
rect 75678 114136 75720 114176
rect 75760 114136 75769 114176
rect 90503 114136 90512 114176
rect 90552 114136 90594 114176
rect 90634 114136 90676 114176
rect 90716 114136 90758 114176
rect 90798 114136 90840 114176
rect 90880 114136 90889 114176
rect 105623 114136 105632 114176
rect 105672 114136 105714 114176
rect 105754 114136 105796 114176
rect 105836 114136 105878 114176
rect 105918 114136 105960 114176
rect 106000 114136 106009 114176
rect 120743 114136 120752 114176
rect 120792 114136 120834 114176
rect 120874 114136 120916 114176
rect 120956 114136 120998 114176
rect 121038 114136 121080 114176
rect 121120 114136 121129 114176
rect 135863 114136 135872 114176
rect 135912 114136 135954 114176
rect 135994 114136 136036 114176
rect 136076 114136 136118 114176
rect 136158 114136 136200 114176
rect 136240 114136 136249 114176
rect 150983 114136 150992 114176
rect 151032 114136 151074 114176
rect 151114 114136 151156 114176
rect 151196 114136 151238 114176
rect 151278 114136 151320 114176
rect 151360 114136 151369 114176
rect 74143 113380 74152 113420
rect 74192 113380 74234 113420
rect 74274 113380 74316 113420
rect 74356 113380 74398 113420
rect 74438 113380 74480 113420
rect 74520 113380 74529 113420
rect 89263 113380 89272 113420
rect 89312 113380 89354 113420
rect 89394 113380 89436 113420
rect 89476 113380 89518 113420
rect 89558 113380 89600 113420
rect 89640 113380 89649 113420
rect 104383 113380 104392 113420
rect 104432 113380 104474 113420
rect 104514 113380 104556 113420
rect 104596 113380 104638 113420
rect 104678 113380 104720 113420
rect 104760 113380 104769 113420
rect 119503 113380 119512 113420
rect 119552 113380 119594 113420
rect 119634 113380 119676 113420
rect 119716 113380 119758 113420
rect 119798 113380 119840 113420
rect 119880 113380 119889 113420
rect 134623 113380 134632 113420
rect 134672 113380 134714 113420
rect 134754 113380 134796 113420
rect 134836 113380 134878 113420
rect 134918 113380 134960 113420
rect 135000 113380 135009 113420
rect 149743 113380 149752 113420
rect 149792 113380 149834 113420
rect 149874 113380 149916 113420
rect 149956 113380 149998 113420
rect 150038 113380 150080 113420
rect 150120 113380 150129 113420
rect 75383 112624 75392 112664
rect 75432 112624 75474 112664
rect 75514 112624 75556 112664
rect 75596 112624 75638 112664
rect 75678 112624 75720 112664
rect 75760 112624 75769 112664
rect 90503 112624 90512 112664
rect 90552 112624 90594 112664
rect 90634 112624 90676 112664
rect 90716 112624 90758 112664
rect 90798 112624 90840 112664
rect 90880 112624 90889 112664
rect 105623 112624 105632 112664
rect 105672 112624 105714 112664
rect 105754 112624 105796 112664
rect 105836 112624 105878 112664
rect 105918 112624 105960 112664
rect 106000 112624 106009 112664
rect 120743 112624 120752 112664
rect 120792 112624 120834 112664
rect 120874 112624 120916 112664
rect 120956 112624 120998 112664
rect 121038 112624 121080 112664
rect 121120 112624 121129 112664
rect 135863 112624 135872 112664
rect 135912 112624 135954 112664
rect 135994 112624 136036 112664
rect 136076 112624 136118 112664
rect 136158 112624 136200 112664
rect 136240 112624 136249 112664
rect 150983 112624 150992 112664
rect 151032 112624 151074 112664
rect 151114 112624 151156 112664
rect 151196 112624 151238 112664
rect 151278 112624 151320 112664
rect 151360 112624 151369 112664
rect 74143 111868 74152 111908
rect 74192 111868 74234 111908
rect 74274 111868 74316 111908
rect 74356 111868 74398 111908
rect 74438 111868 74480 111908
rect 74520 111868 74529 111908
rect 89263 111868 89272 111908
rect 89312 111868 89354 111908
rect 89394 111868 89436 111908
rect 89476 111868 89518 111908
rect 89558 111868 89600 111908
rect 89640 111868 89649 111908
rect 104383 111868 104392 111908
rect 104432 111868 104474 111908
rect 104514 111868 104556 111908
rect 104596 111868 104638 111908
rect 104678 111868 104720 111908
rect 104760 111868 104769 111908
rect 119503 111868 119512 111908
rect 119552 111868 119594 111908
rect 119634 111868 119676 111908
rect 119716 111868 119758 111908
rect 119798 111868 119840 111908
rect 119880 111868 119889 111908
rect 134623 111868 134632 111908
rect 134672 111868 134714 111908
rect 134754 111868 134796 111908
rect 134836 111868 134878 111908
rect 134918 111868 134960 111908
rect 135000 111868 135009 111908
rect 149743 111868 149752 111908
rect 149792 111868 149834 111908
rect 149874 111868 149916 111908
rect 149956 111868 149998 111908
rect 150038 111868 150080 111908
rect 150120 111868 150129 111908
rect 75383 111112 75392 111152
rect 75432 111112 75474 111152
rect 75514 111112 75556 111152
rect 75596 111112 75638 111152
rect 75678 111112 75720 111152
rect 75760 111112 75769 111152
rect 90503 111112 90512 111152
rect 90552 111112 90594 111152
rect 90634 111112 90676 111152
rect 90716 111112 90758 111152
rect 90798 111112 90840 111152
rect 90880 111112 90889 111152
rect 105623 111112 105632 111152
rect 105672 111112 105714 111152
rect 105754 111112 105796 111152
rect 105836 111112 105878 111152
rect 105918 111112 105960 111152
rect 106000 111112 106009 111152
rect 120743 111112 120752 111152
rect 120792 111112 120834 111152
rect 120874 111112 120916 111152
rect 120956 111112 120998 111152
rect 121038 111112 121080 111152
rect 121120 111112 121129 111152
rect 135863 111112 135872 111152
rect 135912 111112 135954 111152
rect 135994 111112 136036 111152
rect 136076 111112 136118 111152
rect 136158 111112 136200 111152
rect 136240 111112 136249 111152
rect 150983 111112 150992 111152
rect 151032 111112 151074 111152
rect 151114 111112 151156 111152
rect 151196 111112 151238 111152
rect 151278 111112 151320 111152
rect 151360 111112 151369 111152
rect 74143 110356 74152 110396
rect 74192 110356 74234 110396
rect 74274 110356 74316 110396
rect 74356 110356 74398 110396
rect 74438 110356 74480 110396
rect 74520 110356 74529 110396
rect 89263 110356 89272 110396
rect 89312 110356 89354 110396
rect 89394 110356 89436 110396
rect 89476 110356 89518 110396
rect 89558 110356 89600 110396
rect 89640 110356 89649 110396
rect 104383 110356 104392 110396
rect 104432 110356 104474 110396
rect 104514 110356 104556 110396
rect 104596 110356 104638 110396
rect 104678 110356 104720 110396
rect 104760 110356 104769 110396
rect 119503 110356 119512 110396
rect 119552 110356 119594 110396
rect 119634 110356 119676 110396
rect 119716 110356 119758 110396
rect 119798 110356 119840 110396
rect 119880 110356 119889 110396
rect 134623 110356 134632 110396
rect 134672 110356 134714 110396
rect 134754 110356 134796 110396
rect 134836 110356 134878 110396
rect 134918 110356 134960 110396
rect 135000 110356 135009 110396
rect 149743 110356 149752 110396
rect 149792 110356 149834 110396
rect 149874 110356 149916 110396
rect 149956 110356 149998 110396
rect 150038 110356 150080 110396
rect 150120 110356 150129 110396
rect 75383 109600 75392 109640
rect 75432 109600 75474 109640
rect 75514 109600 75556 109640
rect 75596 109600 75638 109640
rect 75678 109600 75720 109640
rect 75760 109600 75769 109640
rect 90503 109600 90512 109640
rect 90552 109600 90594 109640
rect 90634 109600 90676 109640
rect 90716 109600 90758 109640
rect 90798 109600 90840 109640
rect 90880 109600 90889 109640
rect 105623 109600 105632 109640
rect 105672 109600 105714 109640
rect 105754 109600 105796 109640
rect 105836 109600 105878 109640
rect 105918 109600 105960 109640
rect 106000 109600 106009 109640
rect 120743 109600 120752 109640
rect 120792 109600 120834 109640
rect 120874 109600 120916 109640
rect 120956 109600 120998 109640
rect 121038 109600 121080 109640
rect 121120 109600 121129 109640
rect 135863 109600 135872 109640
rect 135912 109600 135954 109640
rect 135994 109600 136036 109640
rect 136076 109600 136118 109640
rect 136158 109600 136200 109640
rect 136240 109600 136249 109640
rect 150983 109600 150992 109640
rect 151032 109600 151074 109640
rect 151114 109600 151156 109640
rect 151196 109600 151238 109640
rect 151278 109600 151320 109640
rect 151360 109600 151369 109640
rect 74143 108844 74152 108884
rect 74192 108844 74234 108884
rect 74274 108844 74316 108884
rect 74356 108844 74398 108884
rect 74438 108844 74480 108884
rect 74520 108844 74529 108884
rect 89263 108844 89272 108884
rect 89312 108844 89354 108884
rect 89394 108844 89436 108884
rect 89476 108844 89518 108884
rect 89558 108844 89600 108884
rect 89640 108844 89649 108884
rect 104383 108844 104392 108884
rect 104432 108844 104474 108884
rect 104514 108844 104556 108884
rect 104596 108844 104638 108884
rect 104678 108844 104720 108884
rect 104760 108844 104769 108884
rect 119503 108844 119512 108884
rect 119552 108844 119594 108884
rect 119634 108844 119676 108884
rect 119716 108844 119758 108884
rect 119798 108844 119840 108884
rect 119880 108844 119889 108884
rect 134623 108844 134632 108884
rect 134672 108844 134714 108884
rect 134754 108844 134796 108884
rect 134836 108844 134878 108884
rect 134918 108844 134960 108884
rect 135000 108844 135009 108884
rect 149743 108844 149752 108884
rect 149792 108844 149834 108884
rect 149874 108844 149916 108884
rect 149956 108844 149998 108884
rect 150038 108844 150080 108884
rect 150120 108844 150129 108884
rect 75383 108088 75392 108128
rect 75432 108088 75474 108128
rect 75514 108088 75556 108128
rect 75596 108088 75638 108128
rect 75678 108088 75720 108128
rect 75760 108088 75769 108128
rect 90503 108088 90512 108128
rect 90552 108088 90594 108128
rect 90634 108088 90676 108128
rect 90716 108088 90758 108128
rect 90798 108088 90840 108128
rect 90880 108088 90889 108128
rect 105623 108088 105632 108128
rect 105672 108088 105714 108128
rect 105754 108088 105796 108128
rect 105836 108088 105878 108128
rect 105918 108088 105960 108128
rect 106000 108088 106009 108128
rect 120743 108088 120752 108128
rect 120792 108088 120834 108128
rect 120874 108088 120916 108128
rect 120956 108088 120998 108128
rect 121038 108088 121080 108128
rect 121120 108088 121129 108128
rect 135863 108088 135872 108128
rect 135912 108088 135954 108128
rect 135994 108088 136036 108128
rect 136076 108088 136118 108128
rect 136158 108088 136200 108128
rect 136240 108088 136249 108128
rect 150983 108088 150992 108128
rect 151032 108088 151074 108128
rect 151114 108088 151156 108128
rect 151196 108088 151238 108128
rect 151278 108088 151320 108128
rect 151360 108088 151369 108128
rect 74143 107332 74152 107372
rect 74192 107332 74234 107372
rect 74274 107332 74316 107372
rect 74356 107332 74398 107372
rect 74438 107332 74480 107372
rect 74520 107332 74529 107372
rect 89263 107332 89272 107372
rect 89312 107332 89354 107372
rect 89394 107332 89436 107372
rect 89476 107332 89518 107372
rect 89558 107332 89600 107372
rect 89640 107332 89649 107372
rect 104383 107332 104392 107372
rect 104432 107332 104474 107372
rect 104514 107332 104556 107372
rect 104596 107332 104638 107372
rect 104678 107332 104720 107372
rect 104760 107332 104769 107372
rect 119503 107332 119512 107372
rect 119552 107332 119594 107372
rect 119634 107332 119676 107372
rect 119716 107332 119758 107372
rect 119798 107332 119840 107372
rect 119880 107332 119889 107372
rect 134623 107332 134632 107372
rect 134672 107332 134714 107372
rect 134754 107332 134796 107372
rect 134836 107332 134878 107372
rect 134918 107332 134960 107372
rect 135000 107332 135009 107372
rect 149743 107332 149752 107372
rect 149792 107332 149834 107372
rect 149874 107332 149916 107372
rect 149956 107332 149998 107372
rect 150038 107332 150080 107372
rect 150120 107332 150129 107372
rect 75383 106576 75392 106616
rect 75432 106576 75474 106616
rect 75514 106576 75556 106616
rect 75596 106576 75638 106616
rect 75678 106576 75720 106616
rect 75760 106576 75769 106616
rect 90503 106576 90512 106616
rect 90552 106576 90594 106616
rect 90634 106576 90676 106616
rect 90716 106576 90758 106616
rect 90798 106576 90840 106616
rect 90880 106576 90889 106616
rect 105623 106576 105632 106616
rect 105672 106576 105714 106616
rect 105754 106576 105796 106616
rect 105836 106576 105878 106616
rect 105918 106576 105960 106616
rect 106000 106576 106009 106616
rect 120743 106576 120752 106616
rect 120792 106576 120834 106616
rect 120874 106576 120916 106616
rect 120956 106576 120998 106616
rect 121038 106576 121080 106616
rect 121120 106576 121129 106616
rect 135863 106576 135872 106616
rect 135912 106576 135954 106616
rect 135994 106576 136036 106616
rect 136076 106576 136118 106616
rect 136158 106576 136200 106616
rect 136240 106576 136249 106616
rect 150983 106576 150992 106616
rect 151032 106576 151074 106616
rect 151114 106576 151156 106616
rect 151196 106576 151238 106616
rect 151278 106576 151320 106616
rect 151360 106576 151369 106616
rect 74143 105820 74152 105860
rect 74192 105820 74234 105860
rect 74274 105820 74316 105860
rect 74356 105820 74398 105860
rect 74438 105820 74480 105860
rect 74520 105820 74529 105860
rect 89263 105820 89272 105860
rect 89312 105820 89354 105860
rect 89394 105820 89436 105860
rect 89476 105820 89518 105860
rect 89558 105820 89600 105860
rect 89640 105820 89649 105860
rect 104383 105820 104392 105860
rect 104432 105820 104474 105860
rect 104514 105820 104556 105860
rect 104596 105820 104638 105860
rect 104678 105820 104720 105860
rect 104760 105820 104769 105860
rect 119503 105820 119512 105860
rect 119552 105820 119594 105860
rect 119634 105820 119676 105860
rect 119716 105820 119758 105860
rect 119798 105820 119840 105860
rect 119880 105820 119889 105860
rect 134623 105820 134632 105860
rect 134672 105820 134714 105860
rect 134754 105820 134796 105860
rect 134836 105820 134878 105860
rect 134918 105820 134960 105860
rect 135000 105820 135009 105860
rect 149743 105820 149752 105860
rect 149792 105820 149834 105860
rect 149874 105820 149916 105860
rect 149956 105820 149998 105860
rect 150038 105820 150080 105860
rect 150120 105820 150129 105860
rect 75383 105064 75392 105104
rect 75432 105064 75474 105104
rect 75514 105064 75556 105104
rect 75596 105064 75638 105104
rect 75678 105064 75720 105104
rect 75760 105064 75769 105104
rect 90503 105064 90512 105104
rect 90552 105064 90594 105104
rect 90634 105064 90676 105104
rect 90716 105064 90758 105104
rect 90798 105064 90840 105104
rect 90880 105064 90889 105104
rect 105623 105064 105632 105104
rect 105672 105064 105714 105104
rect 105754 105064 105796 105104
rect 105836 105064 105878 105104
rect 105918 105064 105960 105104
rect 106000 105064 106009 105104
rect 120743 105064 120752 105104
rect 120792 105064 120834 105104
rect 120874 105064 120916 105104
rect 120956 105064 120998 105104
rect 121038 105064 121080 105104
rect 121120 105064 121129 105104
rect 135863 105064 135872 105104
rect 135912 105064 135954 105104
rect 135994 105064 136036 105104
rect 136076 105064 136118 105104
rect 136158 105064 136200 105104
rect 136240 105064 136249 105104
rect 150983 105064 150992 105104
rect 151032 105064 151074 105104
rect 151114 105064 151156 105104
rect 151196 105064 151238 105104
rect 151278 105064 151320 105104
rect 151360 105064 151369 105104
rect 74143 104308 74152 104348
rect 74192 104308 74234 104348
rect 74274 104308 74316 104348
rect 74356 104308 74398 104348
rect 74438 104308 74480 104348
rect 74520 104308 74529 104348
rect 89263 104308 89272 104348
rect 89312 104308 89354 104348
rect 89394 104308 89436 104348
rect 89476 104308 89518 104348
rect 89558 104308 89600 104348
rect 89640 104308 89649 104348
rect 104383 104308 104392 104348
rect 104432 104308 104474 104348
rect 104514 104308 104556 104348
rect 104596 104308 104638 104348
rect 104678 104308 104720 104348
rect 104760 104308 104769 104348
rect 119503 104308 119512 104348
rect 119552 104308 119594 104348
rect 119634 104308 119676 104348
rect 119716 104308 119758 104348
rect 119798 104308 119840 104348
rect 119880 104308 119889 104348
rect 134623 104308 134632 104348
rect 134672 104308 134714 104348
rect 134754 104308 134796 104348
rect 134836 104308 134878 104348
rect 134918 104308 134960 104348
rect 135000 104308 135009 104348
rect 149743 104308 149752 104348
rect 149792 104308 149834 104348
rect 149874 104308 149916 104348
rect 149956 104308 149998 104348
rect 150038 104308 150080 104348
rect 150120 104308 150129 104348
rect 64099 103972 64108 104012
rect 64148 103972 160032 104012
rect 75383 103552 75392 103592
rect 75432 103552 75474 103592
rect 75514 103552 75556 103592
rect 75596 103552 75638 103592
rect 75678 103552 75720 103592
rect 75760 103552 75769 103592
rect 90503 103552 90512 103592
rect 90552 103552 90594 103592
rect 90634 103552 90676 103592
rect 90716 103552 90758 103592
rect 90798 103552 90840 103592
rect 90880 103552 90889 103592
rect 105623 103552 105632 103592
rect 105672 103552 105714 103592
rect 105754 103552 105796 103592
rect 105836 103552 105878 103592
rect 105918 103552 105960 103592
rect 106000 103552 106009 103592
rect 120743 103552 120752 103592
rect 120792 103552 120834 103592
rect 120874 103552 120916 103592
rect 120956 103552 120998 103592
rect 121038 103552 121080 103592
rect 121120 103552 121129 103592
rect 135863 103552 135872 103592
rect 135912 103552 135954 103592
rect 135994 103552 136036 103592
rect 136076 103552 136118 103592
rect 136158 103552 136200 103592
rect 136240 103552 136249 103592
rect 150983 103552 150992 103592
rect 151032 103552 151074 103592
rect 151114 103552 151156 103592
rect 151196 103552 151238 103592
rect 151278 103552 151320 103592
rect 151360 103552 151369 103592
rect 74143 102796 74152 102836
rect 74192 102796 74234 102836
rect 74274 102796 74316 102836
rect 74356 102796 74398 102836
rect 74438 102796 74480 102836
rect 74520 102796 74529 102836
rect 89263 102796 89272 102836
rect 89312 102796 89354 102836
rect 89394 102796 89436 102836
rect 89476 102796 89518 102836
rect 89558 102796 89600 102836
rect 89640 102796 89649 102836
rect 104383 102796 104392 102836
rect 104432 102796 104474 102836
rect 104514 102796 104556 102836
rect 104596 102796 104638 102836
rect 104678 102796 104720 102836
rect 104760 102796 104769 102836
rect 119503 102796 119512 102836
rect 119552 102796 119594 102836
rect 119634 102796 119676 102836
rect 119716 102796 119758 102836
rect 119798 102796 119840 102836
rect 119880 102796 119889 102836
rect 134623 102796 134632 102836
rect 134672 102796 134714 102836
rect 134754 102796 134796 102836
rect 134836 102796 134878 102836
rect 134918 102796 134960 102836
rect 135000 102796 135009 102836
rect 149743 102796 149752 102836
rect 149792 102796 149834 102836
rect 149874 102796 149916 102836
rect 149956 102796 149998 102836
rect 150038 102796 150080 102836
rect 150120 102796 150129 102836
rect 75383 102040 75392 102080
rect 75432 102040 75474 102080
rect 75514 102040 75556 102080
rect 75596 102040 75638 102080
rect 75678 102040 75720 102080
rect 75760 102040 75769 102080
rect 90503 102040 90512 102080
rect 90552 102040 90594 102080
rect 90634 102040 90676 102080
rect 90716 102040 90758 102080
rect 90798 102040 90840 102080
rect 90880 102040 90889 102080
rect 105623 102040 105632 102080
rect 105672 102040 105714 102080
rect 105754 102040 105796 102080
rect 105836 102040 105878 102080
rect 105918 102040 105960 102080
rect 106000 102040 106009 102080
rect 120743 102040 120752 102080
rect 120792 102040 120834 102080
rect 120874 102040 120916 102080
rect 120956 102040 120998 102080
rect 121038 102040 121080 102080
rect 121120 102040 121129 102080
rect 135863 102040 135872 102080
rect 135912 102040 135954 102080
rect 135994 102040 136036 102080
rect 136076 102040 136118 102080
rect 136158 102040 136200 102080
rect 136240 102040 136249 102080
rect 150983 102040 150992 102080
rect 151032 102040 151074 102080
rect 151114 102040 151156 102080
rect 151196 102040 151238 102080
rect 151278 102040 151320 102080
rect 151360 102040 151369 102080
rect 74143 101284 74152 101324
rect 74192 101284 74234 101324
rect 74274 101284 74316 101324
rect 74356 101284 74398 101324
rect 74438 101284 74480 101324
rect 74520 101284 74529 101324
rect 89263 101284 89272 101324
rect 89312 101284 89354 101324
rect 89394 101284 89436 101324
rect 89476 101284 89518 101324
rect 89558 101284 89600 101324
rect 89640 101284 89649 101324
rect 104383 101284 104392 101324
rect 104432 101284 104474 101324
rect 104514 101284 104556 101324
rect 104596 101284 104638 101324
rect 104678 101284 104720 101324
rect 104760 101284 104769 101324
rect 119503 101284 119512 101324
rect 119552 101284 119594 101324
rect 119634 101284 119676 101324
rect 119716 101284 119758 101324
rect 119798 101284 119840 101324
rect 119880 101284 119889 101324
rect 134623 101284 134632 101324
rect 134672 101284 134714 101324
rect 134754 101284 134796 101324
rect 134836 101284 134878 101324
rect 134918 101284 134960 101324
rect 135000 101284 135009 101324
rect 149743 101284 149752 101324
rect 149792 101284 149834 101324
rect 149874 101284 149916 101324
rect 149956 101284 149998 101324
rect 150038 101284 150080 101324
rect 150120 101284 150129 101324
rect 75383 100528 75392 100568
rect 75432 100528 75474 100568
rect 75514 100528 75556 100568
rect 75596 100528 75638 100568
rect 75678 100528 75720 100568
rect 75760 100528 75769 100568
rect 90503 100528 90512 100568
rect 90552 100528 90594 100568
rect 90634 100528 90676 100568
rect 90716 100528 90758 100568
rect 90798 100528 90840 100568
rect 90880 100528 90889 100568
rect 105623 100528 105632 100568
rect 105672 100528 105714 100568
rect 105754 100528 105796 100568
rect 105836 100528 105878 100568
rect 105918 100528 105960 100568
rect 106000 100528 106009 100568
rect 120743 100528 120752 100568
rect 120792 100528 120834 100568
rect 120874 100528 120916 100568
rect 120956 100528 120998 100568
rect 121038 100528 121080 100568
rect 121120 100528 121129 100568
rect 135863 100528 135872 100568
rect 135912 100528 135954 100568
rect 135994 100528 136036 100568
rect 136076 100528 136118 100568
rect 136158 100528 136200 100568
rect 136240 100528 136249 100568
rect 150983 100528 150992 100568
rect 151032 100528 151074 100568
rect 151114 100528 151156 100568
rect 151196 100528 151238 100568
rect 151278 100528 151320 100568
rect 151360 100528 151369 100568
rect 74143 99772 74152 99812
rect 74192 99772 74234 99812
rect 74274 99772 74316 99812
rect 74356 99772 74398 99812
rect 74438 99772 74480 99812
rect 74520 99772 74529 99812
rect 89263 99772 89272 99812
rect 89312 99772 89354 99812
rect 89394 99772 89436 99812
rect 89476 99772 89518 99812
rect 89558 99772 89600 99812
rect 89640 99772 89649 99812
rect 104383 99772 104392 99812
rect 104432 99772 104474 99812
rect 104514 99772 104556 99812
rect 104596 99772 104638 99812
rect 104678 99772 104720 99812
rect 104760 99772 104769 99812
rect 119503 99772 119512 99812
rect 119552 99772 119594 99812
rect 119634 99772 119676 99812
rect 119716 99772 119758 99812
rect 119798 99772 119840 99812
rect 119880 99772 119889 99812
rect 134623 99772 134632 99812
rect 134672 99772 134714 99812
rect 134754 99772 134796 99812
rect 134836 99772 134878 99812
rect 134918 99772 134960 99812
rect 135000 99772 135009 99812
rect 149743 99772 149752 99812
rect 149792 99772 149834 99812
rect 149874 99772 149916 99812
rect 149956 99772 149998 99812
rect 150038 99772 150080 99812
rect 150120 99772 150129 99812
rect 75383 99016 75392 99056
rect 75432 99016 75474 99056
rect 75514 99016 75556 99056
rect 75596 99016 75638 99056
rect 75678 99016 75720 99056
rect 75760 99016 75769 99056
rect 90503 99016 90512 99056
rect 90552 99016 90594 99056
rect 90634 99016 90676 99056
rect 90716 99016 90758 99056
rect 90798 99016 90840 99056
rect 90880 99016 90889 99056
rect 105623 99016 105632 99056
rect 105672 99016 105714 99056
rect 105754 99016 105796 99056
rect 105836 99016 105878 99056
rect 105918 99016 105960 99056
rect 106000 99016 106009 99056
rect 120743 99016 120752 99056
rect 120792 99016 120834 99056
rect 120874 99016 120916 99056
rect 120956 99016 120998 99056
rect 121038 99016 121080 99056
rect 121120 99016 121129 99056
rect 135863 99016 135872 99056
rect 135912 99016 135954 99056
rect 135994 99016 136036 99056
rect 136076 99016 136118 99056
rect 136158 99016 136200 99056
rect 136240 99016 136249 99056
rect 150983 99016 150992 99056
rect 151032 99016 151074 99056
rect 151114 99016 151156 99056
rect 151196 99016 151238 99056
rect 151278 99016 151320 99056
rect 151360 99016 151369 99056
rect 74143 98260 74152 98300
rect 74192 98260 74234 98300
rect 74274 98260 74316 98300
rect 74356 98260 74398 98300
rect 74438 98260 74480 98300
rect 74520 98260 74529 98300
rect 89263 98260 89272 98300
rect 89312 98260 89354 98300
rect 89394 98260 89436 98300
rect 89476 98260 89518 98300
rect 89558 98260 89600 98300
rect 89640 98260 89649 98300
rect 104383 98260 104392 98300
rect 104432 98260 104474 98300
rect 104514 98260 104556 98300
rect 104596 98260 104638 98300
rect 104678 98260 104720 98300
rect 104760 98260 104769 98300
rect 119503 98260 119512 98300
rect 119552 98260 119594 98300
rect 119634 98260 119676 98300
rect 119716 98260 119758 98300
rect 119798 98260 119840 98300
rect 119880 98260 119889 98300
rect 134623 98260 134632 98300
rect 134672 98260 134714 98300
rect 134754 98260 134796 98300
rect 134836 98260 134878 98300
rect 134918 98260 134960 98300
rect 135000 98260 135009 98300
rect 149743 98260 149752 98300
rect 149792 98260 149834 98300
rect 149874 98260 149916 98300
rect 149956 98260 149998 98300
rect 150038 98260 150080 98300
rect 150120 98260 150129 98300
rect 75383 97504 75392 97544
rect 75432 97504 75474 97544
rect 75514 97504 75556 97544
rect 75596 97504 75638 97544
rect 75678 97504 75720 97544
rect 75760 97504 75769 97544
rect 90503 97504 90512 97544
rect 90552 97504 90594 97544
rect 90634 97504 90676 97544
rect 90716 97504 90758 97544
rect 90798 97504 90840 97544
rect 90880 97504 90889 97544
rect 105623 97504 105632 97544
rect 105672 97504 105714 97544
rect 105754 97504 105796 97544
rect 105836 97504 105878 97544
rect 105918 97504 105960 97544
rect 106000 97504 106009 97544
rect 120743 97504 120752 97544
rect 120792 97504 120834 97544
rect 120874 97504 120916 97544
rect 120956 97504 120998 97544
rect 121038 97504 121080 97544
rect 121120 97504 121129 97544
rect 135863 97504 135872 97544
rect 135912 97504 135954 97544
rect 135994 97504 136036 97544
rect 136076 97504 136118 97544
rect 136158 97504 136200 97544
rect 136240 97504 136249 97544
rect 150983 97504 150992 97544
rect 151032 97504 151074 97544
rect 151114 97504 151156 97544
rect 151196 97504 151238 97544
rect 151278 97504 151320 97544
rect 151360 97504 151369 97544
rect 74143 96748 74152 96788
rect 74192 96748 74234 96788
rect 74274 96748 74316 96788
rect 74356 96748 74398 96788
rect 74438 96748 74480 96788
rect 74520 96748 74529 96788
rect 89263 96748 89272 96788
rect 89312 96748 89354 96788
rect 89394 96748 89436 96788
rect 89476 96748 89518 96788
rect 89558 96748 89600 96788
rect 89640 96748 89649 96788
rect 104383 96748 104392 96788
rect 104432 96748 104474 96788
rect 104514 96748 104556 96788
rect 104596 96748 104638 96788
rect 104678 96748 104720 96788
rect 104760 96748 104769 96788
rect 119503 96748 119512 96788
rect 119552 96748 119594 96788
rect 119634 96748 119676 96788
rect 119716 96748 119758 96788
rect 119798 96748 119840 96788
rect 119880 96748 119889 96788
rect 134623 96748 134632 96788
rect 134672 96748 134714 96788
rect 134754 96748 134796 96788
rect 134836 96748 134878 96788
rect 134918 96748 134960 96788
rect 135000 96748 135009 96788
rect 149743 96748 149752 96788
rect 149792 96748 149834 96788
rect 149874 96748 149916 96788
rect 149956 96748 149998 96788
rect 150038 96748 150080 96788
rect 150120 96748 150129 96788
rect 75383 95992 75392 96032
rect 75432 95992 75474 96032
rect 75514 95992 75556 96032
rect 75596 95992 75638 96032
rect 75678 95992 75720 96032
rect 75760 95992 75769 96032
rect 90503 95992 90512 96032
rect 90552 95992 90594 96032
rect 90634 95992 90676 96032
rect 90716 95992 90758 96032
rect 90798 95992 90840 96032
rect 90880 95992 90889 96032
rect 105623 95992 105632 96032
rect 105672 95992 105714 96032
rect 105754 95992 105796 96032
rect 105836 95992 105878 96032
rect 105918 95992 105960 96032
rect 106000 95992 106009 96032
rect 120743 95992 120752 96032
rect 120792 95992 120834 96032
rect 120874 95992 120916 96032
rect 120956 95992 120998 96032
rect 121038 95992 121080 96032
rect 121120 95992 121129 96032
rect 135863 95992 135872 96032
rect 135912 95992 135954 96032
rect 135994 95992 136036 96032
rect 136076 95992 136118 96032
rect 136158 95992 136200 96032
rect 136240 95992 136249 96032
rect 150983 95992 150992 96032
rect 151032 95992 151074 96032
rect 151114 95992 151156 96032
rect 151196 95992 151238 96032
rect 151278 95992 151320 96032
rect 151360 95992 151369 96032
rect 74143 95236 74152 95276
rect 74192 95236 74234 95276
rect 74274 95236 74316 95276
rect 74356 95236 74398 95276
rect 74438 95236 74480 95276
rect 74520 95236 74529 95276
rect 89263 95236 89272 95276
rect 89312 95236 89354 95276
rect 89394 95236 89436 95276
rect 89476 95236 89518 95276
rect 89558 95236 89600 95276
rect 89640 95236 89649 95276
rect 104383 95236 104392 95276
rect 104432 95236 104474 95276
rect 104514 95236 104556 95276
rect 104596 95236 104638 95276
rect 104678 95236 104720 95276
rect 104760 95236 104769 95276
rect 119503 95236 119512 95276
rect 119552 95236 119594 95276
rect 119634 95236 119676 95276
rect 119716 95236 119758 95276
rect 119798 95236 119840 95276
rect 119880 95236 119889 95276
rect 134623 95236 134632 95276
rect 134672 95236 134714 95276
rect 134754 95236 134796 95276
rect 134836 95236 134878 95276
rect 134918 95236 134960 95276
rect 135000 95236 135009 95276
rect 149743 95236 149752 95276
rect 149792 95236 149834 95276
rect 149874 95236 149916 95276
rect 149956 95236 149998 95276
rect 150038 95236 150080 95276
rect 150120 95236 150129 95276
rect 75383 94480 75392 94520
rect 75432 94480 75474 94520
rect 75514 94480 75556 94520
rect 75596 94480 75638 94520
rect 75678 94480 75720 94520
rect 75760 94480 75769 94520
rect 90503 94480 90512 94520
rect 90552 94480 90594 94520
rect 90634 94480 90676 94520
rect 90716 94480 90758 94520
rect 90798 94480 90840 94520
rect 90880 94480 90889 94520
rect 105623 94480 105632 94520
rect 105672 94480 105714 94520
rect 105754 94480 105796 94520
rect 105836 94480 105878 94520
rect 105918 94480 105960 94520
rect 106000 94480 106009 94520
rect 120743 94480 120752 94520
rect 120792 94480 120834 94520
rect 120874 94480 120916 94520
rect 120956 94480 120998 94520
rect 121038 94480 121080 94520
rect 121120 94480 121129 94520
rect 135863 94480 135872 94520
rect 135912 94480 135954 94520
rect 135994 94480 136036 94520
rect 136076 94480 136118 94520
rect 136158 94480 136200 94520
rect 136240 94480 136249 94520
rect 150983 94480 150992 94520
rect 151032 94480 151074 94520
rect 151114 94480 151156 94520
rect 151196 94480 151238 94520
rect 151278 94480 151320 94520
rect 151360 94480 151369 94520
rect 74143 93724 74152 93764
rect 74192 93724 74234 93764
rect 74274 93724 74316 93764
rect 74356 93724 74398 93764
rect 74438 93724 74480 93764
rect 74520 93724 74529 93764
rect 89263 93724 89272 93764
rect 89312 93724 89354 93764
rect 89394 93724 89436 93764
rect 89476 93724 89518 93764
rect 89558 93724 89600 93764
rect 89640 93724 89649 93764
rect 104383 93724 104392 93764
rect 104432 93724 104474 93764
rect 104514 93724 104556 93764
rect 104596 93724 104638 93764
rect 104678 93724 104720 93764
rect 104760 93724 104769 93764
rect 119503 93724 119512 93764
rect 119552 93724 119594 93764
rect 119634 93724 119676 93764
rect 119716 93724 119758 93764
rect 119798 93724 119840 93764
rect 119880 93724 119889 93764
rect 134623 93724 134632 93764
rect 134672 93724 134714 93764
rect 134754 93724 134796 93764
rect 134836 93724 134878 93764
rect 134918 93724 134960 93764
rect 135000 93724 135009 93764
rect 149743 93724 149752 93764
rect 149792 93724 149834 93764
rect 149874 93724 149916 93764
rect 149956 93724 149998 93764
rect 150038 93724 150080 93764
rect 150120 93724 150129 93764
rect 75383 92968 75392 93008
rect 75432 92968 75474 93008
rect 75514 92968 75556 93008
rect 75596 92968 75638 93008
rect 75678 92968 75720 93008
rect 75760 92968 75769 93008
rect 90503 92968 90512 93008
rect 90552 92968 90594 93008
rect 90634 92968 90676 93008
rect 90716 92968 90758 93008
rect 90798 92968 90840 93008
rect 90880 92968 90889 93008
rect 105623 92968 105632 93008
rect 105672 92968 105714 93008
rect 105754 92968 105796 93008
rect 105836 92968 105878 93008
rect 105918 92968 105960 93008
rect 106000 92968 106009 93008
rect 120743 92968 120752 93008
rect 120792 92968 120834 93008
rect 120874 92968 120916 93008
rect 120956 92968 120998 93008
rect 121038 92968 121080 93008
rect 121120 92968 121129 93008
rect 135863 92968 135872 93008
rect 135912 92968 135954 93008
rect 135994 92968 136036 93008
rect 136076 92968 136118 93008
rect 136158 92968 136200 93008
rect 136240 92968 136249 93008
rect 150983 92968 150992 93008
rect 151032 92968 151074 93008
rect 151114 92968 151156 93008
rect 151196 92968 151238 93008
rect 151278 92968 151320 93008
rect 151360 92968 151369 93008
rect 74143 92212 74152 92252
rect 74192 92212 74234 92252
rect 74274 92212 74316 92252
rect 74356 92212 74398 92252
rect 74438 92212 74480 92252
rect 74520 92212 74529 92252
rect 89263 92212 89272 92252
rect 89312 92212 89354 92252
rect 89394 92212 89436 92252
rect 89476 92212 89518 92252
rect 89558 92212 89600 92252
rect 89640 92212 89649 92252
rect 104383 92212 104392 92252
rect 104432 92212 104474 92252
rect 104514 92212 104556 92252
rect 104596 92212 104638 92252
rect 104678 92212 104720 92252
rect 104760 92212 104769 92252
rect 119503 92212 119512 92252
rect 119552 92212 119594 92252
rect 119634 92212 119676 92252
rect 119716 92212 119758 92252
rect 119798 92212 119840 92252
rect 119880 92212 119889 92252
rect 134623 92212 134632 92252
rect 134672 92212 134714 92252
rect 134754 92212 134796 92252
rect 134836 92212 134878 92252
rect 134918 92212 134960 92252
rect 135000 92212 135009 92252
rect 149743 92212 149752 92252
rect 149792 92212 149834 92252
rect 149874 92212 149916 92252
rect 149956 92212 149998 92252
rect 150038 92212 150080 92252
rect 150120 92212 150129 92252
rect 75383 91456 75392 91496
rect 75432 91456 75474 91496
rect 75514 91456 75556 91496
rect 75596 91456 75638 91496
rect 75678 91456 75720 91496
rect 75760 91456 75769 91496
rect 90503 91456 90512 91496
rect 90552 91456 90594 91496
rect 90634 91456 90676 91496
rect 90716 91456 90758 91496
rect 90798 91456 90840 91496
rect 90880 91456 90889 91496
rect 105623 91456 105632 91496
rect 105672 91456 105714 91496
rect 105754 91456 105796 91496
rect 105836 91456 105878 91496
rect 105918 91456 105960 91496
rect 106000 91456 106009 91496
rect 120743 91456 120752 91496
rect 120792 91456 120834 91496
rect 120874 91456 120916 91496
rect 120956 91456 120998 91496
rect 121038 91456 121080 91496
rect 121120 91456 121129 91496
rect 135863 91456 135872 91496
rect 135912 91456 135954 91496
rect 135994 91456 136036 91496
rect 136076 91456 136118 91496
rect 136158 91456 136200 91496
rect 136240 91456 136249 91496
rect 150983 91456 150992 91496
rect 151032 91456 151074 91496
rect 151114 91456 151156 91496
rect 151196 91456 151238 91496
rect 151278 91456 151320 91496
rect 151360 91456 151369 91496
rect 74143 90700 74152 90740
rect 74192 90700 74234 90740
rect 74274 90700 74316 90740
rect 74356 90700 74398 90740
rect 74438 90700 74480 90740
rect 74520 90700 74529 90740
rect 89263 90700 89272 90740
rect 89312 90700 89354 90740
rect 89394 90700 89436 90740
rect 89476 90700 89518 90740
rect 89558 90700 89600 90740
rect 89640 90700 89649 90740
rect 104383 90700 104392 90740
rect 104432 90700 104474 90740
rect 104514 90700 104556 90740
rect 104596 90700 104638 90740
rect 104678 90700 104720 90740
rect 104760 90700 104769 90740
rect 119503 90700 119512 90740
rect 119552 90700 119594 90740
rect 119634 90700 119676 90740
rect 119716 90700 119758 90740
rect 119798 90700 119840 90740
rect 119880 90700 119889 90740
rect 134623 90700 134632 90740
rect 134672 90700 134714 90740
rect 134754 90700 134796 90740
rect 134836 90700 134878 90740
rect 134918 90700 134960 90740
rect 135000 90700 135009 90740
rect 149743 90700 149752 90740
rect 149792 90700 149834 90740
rect 149874 90700 149916 90740
rect 149956 90700 149998 90740
rect 150038 90700 150080 90740
rect 150120 90700 150129 90740
rect 75383 89944 75392 89984
rect 75432 89944 75474 89984
rect 75514 89944 75556 89984
rect 75596 89944 75638 89984
rect 75678 89944 75720 89984
rect 75760 89944 75769 89984
rect 90503 89944 90512 89984
rect 90552 89944 90594 89984
rect 90634 89944 90676 89984
rect 90716 89944 90758 89984
rect 90798 89944 90840 89984
rect 90880 89944 90889 89984
rect 105623 89944 105632 89984
rect 105672 89944 105714 89984
rect 105754 89944 105796 89984
rect 105836 89944 105878 89984
rect 105918 89944 105960 89984
rect 106000 89944 106009 89984
rect 120743 89944 120752 89984
rect 120792 89944 120834 89984
rect 120874 89944 120916 89984
rect 120956 89944 120998 89984
rect 121038 89944 121080 89984
rect 121120 89944 121129 89984
rect 135863 89944 135872 89984
rect 135912 89944 135954 89984
rect 135994 89944 136036 89984
rect 136076 89944 136118 89984
rect 136158 89944 136200 89984
rect 136240 89944 136249 89984
rect 150983 89944 150992 89984
rect 151032 89944 151074 89984
rect 151114 89944 151156 89984
rect 151196 89944 151238 89984
rect 151278 89944 151320 89984
rect 151360 89944 151369 89984
rect 74143 89188 74152 89228
rect 74192 89188 74234 89228
rect 74274 89188 74316 89228
rect 74356 89188 74398 89228
rect 74438 89188 74480 89228
rect 74520 89188 74529 89228
rect 89263 89188 89272 89228
rect 89312 89188 89354 89228
rect 89394 89188 89436 89228
rect 89476 89188 89518 89228
rect 89558 89188 89600 89228
rect 89640 89188 89649 89228
rect 104383 89188 104392 89228
rect 104432 89188 104474 89228
rect 104514 89188 104556 89228
rect 104596 89188 104638 89228
rect 104678 89188 104720 89228
rect 104760 89188 104769 89228
rect 119503 89188 119512 89228
rect 119552 89188 119594 89228
rect 119634 89188 119676 89228
rect 119716 89188 119758 89228
rect 119798 89188 119840 89228
rect 119880 89188 119889 89228
rect 134623 89188 134632 89228
rect 134672 89188 134714 89228
rect 134754 89188 134796 89228
rect 134836 89188 134878 89228
rect 134918 89188 134960 89228
rect 135000 89188 135009 89228
rect 149743 89188 149752 89228
rect 149792 89188 149834 89228
rect 149874 89188 149916 89228
rect 149956 89188 149998 89228
rect 150038 89188 150080 89228
rect 150120 89188 150129 89228
rect 75383 88432 75392 88472
rect 75432 88432 75474 88472
rect 75514 88432 75556 88472
rect 75596 88432 75638 88472
rect 75678 88432 75720 88472
rect 75760 88432 75769 88472
rect 90503 88432 90512 88472
rect 90552 88432 90594 88472
rect 90634 88432 90676 88472
rect 90716 88432 90758 88472
rect 90798 88432 90840 88472
rect 90880 88432 90889 88472
rect 105623 88432 105632 88472
rect 105672 88432 105714 88472
rect 105754 88432 105796 88472
rect 105836 88432 105878 88472
rect 105918 88432 105960 88472
rect 106000 88432 106009 88472
rect 120743 88432 120752 88472
rect 120792 88432 120834 88472
rect 120874 88432 120916 88472
rect 120956 88432 120998 88472
rect 121038 88432 121080 88472
rect 121120 88432 121129 88472
rect 135863 88432 135872 88472
rect 135912 88432 135954 88472
rect 135994 88432 136036 88472
rect 136076 88432 136118 88472
rect 136158 88432 136200 88472
rect 136240 88432 136249 88472
rect 150983 88432 150992 88472
rect 151032 88432 151074 88472
rect 151114 88432 151156 88472
rect 151196 88432 151238 88472
rect 151278 88432 151320 88472
rect 151360 88432 151369 88472
rect 64099 88012 64108 88052
rect 64148 88012 160032 88052
rect 74143 87676 74152 87716
rect 74192 87676 74234 87716
rect 74274 87676 74316 87716
rect 74356 87676 74398 87716
rect 74438 87676 74480 87716
rect 74520 87676 74529 87716
rect 89263 87676 89272 87716
rect 89312 87676 89354 87716
rect 89394 87676 89436 87716
rect 89476 87676 89518 87716
rect 89558 87676 89600 87716
rect 89640 87676 89649 87716
rect 104383 87676 104392 87716
rect 104432 87676 104474 87716
rect 104514 87676 104556 87716
rect 104596 87676 104638 87716
rect 104678 87676 104720 87716
rect 104760 87676 104769 87716
rect 119503 87676 119512 87716
rect 119552 87676 119594 87716
rect 119634 87676 119676 87716
rect 119716 87676 119758 87716
rect 119798 87676 119840 87716
rect 119880 87676 119889 87716
rect 134623 87676 134632 87716
rect 134672 87676 134714 87716
rect 134754 87676 134796 87716
rect 134836 87676 134878 87716
rect 134918 87676 134960 87716
rect 135000 87676 135009 87716
rect 149743 87676 149752 87716
rect 149792 87676 149834 87716
rect 149874 87676 149916 87716
rect 149956 87676 149998 87716
rect 150038 87676 150080 87716
rect 150120 87676 150129 87716
rect 75383 86920 75392 86960
rect 75432 86920 75474 86960
rect 75514 86920 75556 86960
rect 75596 86920 75638 86960
rect 75678 86920 75720 86960
rect 75760 86920 75769 86960
rect 90503 86920 90512 86960
rect 90552 86920 90594 86960
rect 90634 86920 90676 86960
rect 90716 86920 90758 86960
rect 90798 86920 90840 86960
rect 90880 86920 90889 86960
rect 105623 86920 105632 86960
rect 105672 86920 105714 86960
rect 105754 86920 105796 86960
rect 105836 86920 105878 86960
rect 105918 86920 105960 86960
rect 106000 86920 106009 86960
rect 120743 86920 120752 86960
rect 120792 86920 120834 86960
rect 120874 86920 120916 86960
rect 120956 86920 120998 86960
rect 121038 86920 121080 86960
rect 121120 86920 121129 86960
rect 135863 86920 135872 86960
rect 135912 86920 135954 86960
rect 135994 86920 136036 86960
rect 136076 86920 136118 86960
rect 136158 86920 136200 86960
rect 136240 86920 136249 86960
rect 150983 86920 150992 86960
rect 151032 86920 151074 86960
rect 151114 86920 151156 86960
rect 151196 86920 151238 86960
rect 151278 86920 151320 86960
rect 151360 86920 151369 86960
rect 74143 86164 74152 86204
rect 74192 86164 74234 86204
rect 74274 86164 74316 86204
rect 74356 86164 74398 86204
rect 74438 86164 74480 86204
rect 74520 86164 74529 86204
rect 89263 86164 89272 86204
rect 89312 86164 89354 86204
rect 89394 86164 89436 86204
rect 89476 86164 89518 86204
rect 89558 86164 89600 86204
rect 89640 86164 89649 86204
rect 104383 86164 104392 86204
rect 104432 86164 104474 86204
rect 104514 86164 104556 86204
rect 104596 86164 104638 86204
rect 104678 86164 104720 86204
rect 104760 86164 104769 86204
rect 119503 86164 119512 86204
rect 119552 86164 119594 86204
rect 119634 86164 119676 86204
rect 119716 86164 119758 86204
rect 119798 86164 119840 86204
rect 119880 86164 119889 86204
rect 134623 86164 134632 86204
rect 134672 86164 134714 86204
rect 134754 86164 134796 86204
rect 134836 86164 134878 86204
rect 134918 86164 134960 86204
rect 135000 86164 135009 86204
rect 149743 86164 149752 86204
rect 149792 86164 149834 86204
rect 149874 86164 149916 86204
rect 149956 86164 149998 86204
rect 150038 86164 150080 86204
rect 150120 86164 150129 86204
rect 75383 85408 75392 85448
rect 75432 85408 75474 85448
rect 75514 85408 75556 85448
rect 75596 85408 75638 85448
rect 75678 85408 75720 85448
rect 75760 85408 75769 85448
rect 90503 85408 90512 85448
rect 90552 85408 90594 85448
rect 90634 85408 90676 85448
rect 90716 85408 90758 85448
rect 90798 85408 90840 85448
rect 90880 85408 90889 85448
rect 105623 85408 105632 85448
rect 105672 85408 105714 85448
rect 105754 85408 105796 85448
rect 105836 85408 105878 85448
rect 105918 85408 105960 85448
rect 106000 85408 106009 85448
rect 120743 85408 120752 85448
rect 120792 85408 120834 85448
rect 120874 85408 120916 85448
rect 120956 85408 120998 85448
rect 121038 85408 121080 85448
rect 121120 85408 121129 85448
rect 135863 85408 135872 85448
rect 135912 85408 135954 85448
rect 135994 85408 136036 85448
rect 136076 85408 136118 85448
rect 136158 85408 136200 85448
rect 136240 85408 136249 85448
rect 150983 85408 150992 85448
rect 151032 85408 151074 85448
rect 151114 85408 151156 85448
rect 151196 85408 151238 85448
rect 151278 85408 151320 85448
rect 151360 85408 151369 85448
rect 74143 84652 74152 84692
rect 74192 84652 74234 84692
rect 74274 84652 74316 84692
rect 74356 84652 74398 84692
rect 74438 84652 74480 84692
rect 74520 84652 74529 84692
rect 89263 84652 89272 84692
rect 89312 84652 89354 84692
rect 89394 84652 89436 84692
rect 89476 84652 89518 84692
rect 89558 84652 89600 84692
rect 89640 84652 89649 84692
rect 104383 84652 104392 84692
rect 104432 84652 104474 84692
rect 104514 84652 104556 84692
rect 104596 84652 104638 84692
rect 104678 84652 104720 84692
rect 104760 84652 104769 84692
rect 119503 84652 119512 84692
rect 119552 84652 119594 84692
rect 119634 84652 119676 84692
rect 119716 84652 119758 84692
rect 119798 84652 119840 84692
rect 119880 84652 119889 84692
rect 134623 84652 134632 84692
rect 134672 84652 134714 84692
rect 134754 84652 134796 84692
rect 134836 84652 134878 84692
rect 134918 84652 134960 84692
rect 135000 84652 135009 84692
rect 149743 84652 149752 84692
rect 149792 84652 149834 84692
rect 149874 84652 149916 84692
rect 149956 84652 149998 84692
rect 150038 84652 150080 84692
rect 150120 84652 150129 84692
rect 75383 83896 75392 83936
rect 75432 83896 75474 83936
rect 75514 83896 75556 83936
rect 75596 83896 75638 83936
rect 75678 83896 75720 83936
rect 75760 83896 75769 83936
rect 90503 83896 90512 83936
rect 90552 83896 90594 83936
rect 90634 83896 90676 83936
rect 90716 83896 90758 83936
rect 90798 83896 90840 83936
rect 90880 83896 90889 83936
rect 105623 83896 105632 83936
rect 105672 83896 105714 83936
rect 105754 83896 105796 83936
rect 105836 83896 105878 83936
rect 105918 83896 105960 83936
rect 106000 83896 106009 83936
rect 120743 83896 120752 83936
rect 120792 83896 120834 83936
rect 120874 83896 120916 83936
rect 120956 83896 120998 83936
rect 121038 83896 121080 83936
rect 121120 83896 121129 83936
rect 135863 83896 135872 83936
rect 135912 83896 135954 83936
rect 135994 83896 136036 83936
rect 136076 83896 136118 83936
rect 136158 83896 136200 83936
rect 136240 83896 136249 83936
rect 150983 83896 150992 83936
rect 151032 83896 151074 83936
rect 151114 83896 151156 83936
rect 151196 83896 151238 83936
rect 151278 83896 151320 83936
rect 151360 83896 151369 83936
rect 74143 83140 74152 83180
rect 74192 83140 74234 83180
rect 74274 83140 74316 83180
rect 74356 83140 74398 83180
rect 74438 83140 74480 83180
rect 74520 83140 74529 83180
rect 89263 83140 89272 83180
rect 89312 83140 89354 83180
rect 89394 83140 89436 83180
rect 89476 83140 89518 83180
rect 89558 83140 89600 83180
rect 89640 83140 89649 83180
rect 104383 83140 104392 83180
rect 104432 83140 104474 83180
rect 104514 83140 104556 83180
rect 104596 83140 104638 83180
rect 104678 83140 104720 83180
rect 104760 83140 104769 83180
rect 119503 83140 119512 83180
rect 119552 83140 119594 83180
rect 119634 83140 119676 83180
rect 119716 83140 119758 83180
rect 119798 83140 119840 83180
rect 119880 83140 119889 83180
rect 134623 83140 134632 83180
rect 134672 83140 134714 83180
rect 134754 83140 134796 83180
rect 134836 83140 134878 83180
rect 134918 83140 134960 83180
rect 135000 83140 135009 83180
rect 149743 83140 149752 83180
rect 149792 83140 149834 83180
rect 149874 83140 149916 83180
rect 149956 83140 149998 83180
rect 150038 83140 150080 83180
rect 150120 83140 150129 83180
rect 75383 82384 75392 82424
rect 75432 82384 75474 82424
rect 75514 82384 75556 82424
rect 75596 82384 75638 82424
rect 75678 82384 75720 82424
rect 75760 82384 75769 82424
rect 90503 82384 90512 82424
rect 90552 82384 90594 82424
rect 90634 82384 90676 82424
rect 90716 82384 90758 82424
rect 90798 82384 90840 82424
rect 90880 82384 90889 82424
rect 105623 82384 105632 82424
rect 105672 82384 105714 82424
rect 105754 82384 105796 82424
rect 105836 82384 105878 82424
rect 105918 82384 105960 82424
rect 106000 82384 106009 82424
rect 120743 82384 120752 82424
rect 120792 82384 120834 82424
rect 120874 82384 120916 82424
rect 120956 82384 120998 82424
rect 121038 82384 121080 82424
rect 121120 82384 121129 82424
rect 135863 82384 135872 82424
rect 135912 82384 135954 82424
rect 135994 82384 136036 82424
rect 136076 82384 136118 82424
rect 136158 82384 136200 82424
rect 136240 82384 136249 82424
rect 150983 82384 150992 82424
rect 151032 82384 151074 82424
rect 151114 82384 151156 82424
rect 151196 82384 151238 82424
rect 151278 82384 151320 82424
rect 151360 82384 151369 82424
rect 74143 81628 74152 81668
rect 74192 81628 74234 81668
rect 74274 81628 74316 81668
rect 74356 81628 74398 81668
rect 74438 81628 74480 81668
rect 74520 81628 74529 81668
rect 89263 81628 89272 81668
rect 89312 81628 89354 81668
rect 89394 81628 89436 81668
rect 89476 81628 89518 81668
rect 89558 81628 89600 81668
rect 89640 81628 89649 81668
rect 104383 81628 104392 81668
rect 104432 81628 104474 81668
rect 104514 81628 104556 81668
rect 104596 81628 104638 81668
rect 104678 81628 104720 81668
rect 104760 81628 104769 81668
rect 119503 81628 119512 81668
rect 119552 81628 119594 81668
rect 119634 81628 119676 81668
rect 119716 81628 119758 81668
rect 119798 81628 119840 81668
rect 119880 81628 119889 81668
rect 134623 81628 134632 81668
rect 134672 81628 134714 81668
rect 134754 81628 134796 81668
rect 134836 81628 134878 81668
rect 134918 81628 134960 81668
rect 135000 81628 135009 81668
rect 149743 81628 149752 81668
rect 149792 81628 149834 81668
rect 149874 81628 149916 81668
rect 149956 81628 149998 81668
rect 150038 81628 150080 81668
rect 150120 81628 150129 81668
rect 75383 80872 75392 80912
rect 75432 80872 75474 80912
rect 75514 80872 75556 80912
rect 75596 80872 75638 80912
rect 75678 80872 75720 80912
rect 75760 80872 75769 80912
rect 90503 80872 90512 80912
rect 90552 80872 90594 80912
rect 90634 80872 90676 80912
rect 90716 80872 90758 80912
rect 90798 80872 90840 80912
rect 90880 80872 90889 80912
rect 105623 80872 105632 80912
rect 105672 80872 105714 80912
rect 105754 80872 105796 80912
rect 105836 80872 105878 80912
rect 105918 80872 105960 80912
rect 106000 80872 106009 80912
rect 120743 80872 120752 80912
rect 120792 80872 120834 80912
rect 120874 80872 120916 80912
rect 120956 80872 120998 80912
rect 121038 80872 121080 80912
rect 121120 80872 121129 80912
rect 135863 80872 135872 80912
rect 135912 80872 135954 80912
rect 135994 80872 136036 80912
rect 136076 80872 136118 80912
rect 136158 80872 136200 80912
rect 136240 80872 136249 80912
rect 150983 80872 150992 80912
rect 151032 80872 151074 80912
rect 151114 80872 151156 80912
rect 151196 80872 151238 80912
rect 151278 80872 151320 80912
rect 151360 80872 151369 80912
rect 74143 80116 74152 80156
rect 74192 80116 74234 80156
rect 74274 80116 74316 80156
rect 74356 80116 74398 80156
rect 74438 80116 74480 80156
rect 74520 80116 74529 80156
rect 89263 80116 89272 80156
rect 89312 80116 89354 80156
rect 89394 80116 89436 80156
rect 89476 80116 89518 80156
rect 89558 80116 89600 80156
rect 89640 80116 89649 80156
rect 104383 80116 104392 80156
rect 104432 80116 104474 80156
rect 104514 80116 104556 80156
rect 104596 80116 104638 80156
rect 104678 80116 104720 80156
rect 104760 80116 104769 80156
rect 119503 80116 119512 80156
rect 119552 80116 119594 80156
rect 119634 80116 119676 80156
rect 119716 80116 119758 80156
rect 119798 80116 119840 80156
rect 119880 80116 119889 80156
rect 134623 80116 134632 80156
rect 134672 80116 134714 80156
rect 134754 80116 134796 80156
rect 134836 80116 134878 80156
rect 134918 80116 134960 80156
rect 135000 80116 135009 80156
rect 149743 80116 149752 80156
rect 149792 80116 149834 80156
rect 149874 80116 149916 80156
rect 149956 80116 149998 80156
rect 150038 80116 150080 80156
rect 150120 80116 150129 80156
rect 75383 79360 75392 79400
rect 75432 79360 75474 79400
rect 75514 79360 75556 79400
rect 75596 79360 75638 79400
rect 75678 79360 75720 79400
rect 75760 79360 75769 79400
rect 90503 79360 90512 79400
rect 90552 79360 90594 79400
rect 90634 79360 90676 79400
rect 90716 79360 90758 79400
rect 90798 79360 90840 79400
rect 90880 79360 90889 79400
rect 105623 79360 105632 79400
rect 105672 79360 105714 79400
rect 105754 79360 105796 79400
rect 105836 79360 105878 79400
rect 105918 79360 105960 79400
rect 106000 79360 106009 79400
rect 120743 79360 120752 79400
rect 120792 79360 120834 79400
rect 120874 79360 120916 79400
rect 120956 79360 120998 79400
rect 121038 79360 121080 79400
rect 121120 79360 121129 79400
rect 135863 79360 135872 79400
rect 135912 79360 135954 79400
rect 135994 79360 136036 79400
rect 136076 79360 136118 79400
rect 136158 79360 136200 79400
rect 136240 79360 136249 79400
rect 150983 79360 150992 79400
rect 151032 79360 151074 79400
rect 151114 79360 151156 79400
rect 151196 79360 151238 79400
rect 151278 79360 151320 79400
rect 151360 79360 151369 79400
rect 74143 78604 74152 78644
rect 74192 78604 74234 78644
rect 74274 78604 74316 78644
rect 74356 78604 74398 78644
rect 74438 78604 74480 78644
rect 74520 78604 74529 78644
rect 89263 78604 89272 78644
rect 89312 78604 89354 78644
rect 89394 78604 89436 78644
rect 89476 78604 89518 78644
rect 89558 78604 89600 78644
rect 89640 78604 89649 78644
rect 104383 78604 104392 78644
rect 104432 78604 104474 78644
rect 104514 78604 104556 78644
rect 104596 78604 104638 78644
rect 104678 78604 104720 78644
rect 104760 78604 104769 78644
rect 119503 78604 119512 78644
rect 119552 78604 119594 78644
rect 119634 78604 119676 78644
rect 119716 78604 119758 78644
rect 119798 78604 119840 78644
rect 119880 78604 119889 78644
rect 134623 78604 134632 78644
rect 134672 78604 134714 78644
rect 134754 78604 134796 78644
rect 134836 78604 134878 78644
rect 134918 78604 134960 78644
rect 135000 78604 135009 78644
rect 149743 78604 149752 78644
rect 149792 78604 149834 78644
rect 149874 78604 149916 78644
rect 149956 78604 149998 78644
rect 150038 78604 150080 78644
rect 150120 78604 150129 78644
rect 75383 77848 75392 77888
rect 75432 77848 75474 77888
rect 75514 77848 75556 77888
rect 75596 77848 75638 77888
rect 75678 77848 75720 77888
rect 75760 77848 75769 77888
rect 90503 77848 90512 77888
rect 90552 77848 90594 77888
rect 90634 77848 90676 77888
rect 90716 77848 90758 77888
rect 90798 77848 90840 77888
rect 90880 77848 90889 77888
rect 105623 77848 105632 77888
rect 105672 77848 105714 77888
rect 105754 77848 105796 77888
rect 105836 77848 105878 77888
rect 105918 77848 105960 77888
rect 106000 77848 106009 77888
rect 120743 77848 120752 77888
rect 120792 77848 120834 77888
rect 120874 77848 120916 77888
rect 120956 77848 120998 77888
rect 121038 77848 121080 77888
rect 121120 77848 121129 77888
rect 135863 77848 135872 77888
rect 135912 77848 135954 77888
rect 135994 77848 136036 77888
rect 136076 77848 136118 77888
rect 136158 77848 136200 77888
rect 136240 77848 136249 77888
rect 150983 77848 150992 77888
rect 151032 77848 151074 77888
rect 151114 77848 151156 77888
rect 151196 77848 151238 77888
rect 151278 77848 151320 77888
rect 151360 77848 151369 77888
rect 74143 77092 74152 77132
rect 74192 77092 74234 77132
rect 74274 77092 74316 77132
rect 74356 77092 74398 77132
rect 74438 77092 74480 77132
rect 74520 77092 74529 77132
rect 89263 77092 89272 77132
rect 89312 77092 89354 77132
rect 89394 77092 89436 77132
rect 89476 77092 89518 77132
rect 89558 77092 89600 77132
rect 89640 77092 89649 77132
rect 104383 77092 104392 77132
rect 104432 77092 104474 77132
rect 104514 77092 104556 77132
rect 104596 77092 104638 77132
rect 104678 77092 104720 77132
rect 104760 77092 104769 77132
rect 119503 77092 119512 77132
rect 119552 77092 119594 77132
rect 119634 77092 119676 77132
rect 119716 77092 119758 77132
rect 119798 77092 119840 77132
rect 119880 77092 119889 77132
rect 134623 77092 134632 77132
rect 134672 77092 134714 77132
rect 134754 77092 134796 77132
rect 134836 77092 134878 77132
rect 134918 77092 134960 77132
rect 135000 77092 135009 77132
rect 149743 77092 149752 77132
rect 149792 77092 149834 77132
rect 149874 77092 149916 77132
rect 149956 77092 149998 77132
rect 150038 77092 150080 77132
rect 150120 77092 150129 77132
rect 75383 76336 75392 76376
rect 75432 76336 75474 76376
rect 75514 76336 75556 76376
rect 75596 76336 75638 76376
rect 75678 76336 75720 76376
rect 75760 76336 75769 76376
rect 90503 76336 90512 76376
rect 90552 76336 90594 76376
rect 90634 76336 90676 76376
rect 90716 76336 90758 76376
rect 90798 76336 90840 76376
rect 90880 76336 90889 76376
rect 105623 76336 105632 76376
rect 105672 76336 105714 76376
rect 105754 76336 105796 76376
rect 105836 76336 105878 76376
rect 105918 76336 105960 76376
rect 106000 76336 106009 76376
rect 120743 76336 120752 76376
rect 120792 76336 120834 76376
rect 120874 76336 120916 76376
rect 120956 76336 120998 76376
rect 121038 76336 121080 76376
rect 121120 76336 121129 76376
rect 135863 76336 135872 76376
rect 135912 76336 135954 76376
rect 135994 76336 136036 76376
rect 136076 76336 136118 76376
rect 136158 76336 136200 76376
rect 136240 76336 136249 76376
rect 150983 76336 150992 76376
rect 151032 76336 151074 76376
rect 151114 76336 151156 76376
rect 151196 76336 151238 76376
rect 151278 76336 151320 76376
rect 151360 76336 151369 76376
rect 74143 75580 74152 75620
rect 74192 75580 74234 75620
rect 74274 75580 74316 75620
rect 74356 75580 74398 75620
rect 74438 75580 74480 75620
rect 74520 75580 74529 75620
rect 89263 75580 89272 75620
rect 89312 75580 89354 75620
rect 89394 75580 89436 75620
rect 89476 75580 89518 75620
rect 89558 75580 89600 75620
rect 89640 75580 89649 75620
rect 104383 75580 104392 75620
rect 104432 75580 104474 75620
rect 104514 75580 104556 75620
rect 104596 75580 104638 75620
rect 104678 75580 104720 75620
rect 104760 75580 104769 75620
rect 119503 75580 119512 75620
rect 119552 75580 119594 75620
rect 119634 75580 119676 75620
rect 119716 75580 119758 75620
rect 119798 75580 119840 75620
rect 119880 75580 119889 75620
rect 134623 75580 134632 75620
rect 134672 75580 134714 75620
rect 134754 75580 134796 75620
rect 134836 75580 134878 75620
rect 134918 75580 134960 75620
rect 135000 75580 135009 75620
rect 149743 75580 149752 75620
rect 149792 75580 149834 75620
rect 149874 75580 149916 75620
rect 149956 75580 149998 75620
rect 150038 75580 150080 75620
rect 150120 75580 150129 75620
rect 75383 74824 75392 74864
rect 75432 74824 75474 74864
rect 75514 74824 75556 74864
rect 75596 74824 75638 74864
rect 75678 74824 75720 74864
rect 75760 74824 75769 74864
rect 90503 74824 90512 74864
rect 90552 74824 90594 74864
rect 90634 74824 90676 74864
rect 90716 74824 90758 74864
rect 90798 74824 90840 74864
rect 90880 74824 90889 74864
rect 105623 74824 105632 74864
rect 105672 74824 105714 74864
rect 105754 74824 105796 74864
rect 105836 74824 105878 74864
rect 105918 74824 105960 74864
rect 106000 74824 106009 74864
rect 120743 74824 120752 74864
rect 120792 74824 120834 74864
rect 120874 74824 120916 74864
rect 120956 74824 120998 74864
rect 121038 74824 121080 74864
rect 121120 74824 121129 74864
rect 135863 74824 135872 74864
rect 135912 74824 135954 74864
rect 135994 74824 136036 74864
rect 136076 74824 136118 74864
rect 136158 74824 136200 74864
rect 136240 74824 136249 74864
rect 150983 74824 150992 74864
rect 151032 74824 151074 74864
rect 151114 74824 151156 74864
rect 151196 74824 151238 74864
rect 151278 74824 151320 74864
rect 151360 74824 151369 74864
rect 74143 74068 74152 74108
rect 74192 74068 74234 74108
rect 74274 74068 74316 74108
rect 74356 74068 74398 74108
rect 74438 74068 74480 74108
rect 74520 74068 74529 74108
rect 89263 74068 89272 74108
rect 89312 74068 89354 74108
rect 89394 74068 89436 74108
rect 89476 74068 89518 74108
rect 89558 74068 89600 74108
rect 89640 74068 89649 74108
rect 104383 74068 104392 74108
rect 104432 74068 104474 74108
rect 104514 74068 104556 74108
rect 104596 74068 104638 74108
rect 104678 74068 104720 74108
rect 104760 74068 104769 74108
rect 119503 74068 119512 74108
rect 119552 74068 119594 74108
rect 119634 74068 119676 74108
rect 119716 74068 119758 74108
rect 119798 74068 119840 74108
rect 119880 74068 119889 74108
rect 134623 74068 134632 74108
rect 134672 74068 134714 74108
rect 134754 74068 134796 74108
rect 134836 74068 134878 74108
rect 134918 74068 134960 74108
rect 135000 74068 135009 74108
rect 149743 74068 149752 74108
rect 149792 74068 149834 74108
rect 149874 74068 149916 74108
rect 149956 74068 149998 74108
rect 150038 74068 150080 74108
rect 150120 74068 150129 74108
rect 75383 73312 75392 73352
rect 75432 73312 75474 73352
rect 75514 73312 75556 73352
rect 75596 73312 75638 73352
rect 75678 73312 75720 73352
rect 75760 73312 75769 73352
rect 90503 73312 90512 73352
rect 90552 73312 90594 73352
rect 90634 73312 90676 73352
rect 90716 73312 90758 73352
rect 90798 73312 90840 73352
rect 90880 73312 90889 73352
rect 105623 73312 105632 73352
rect 105672 73312 105714 73352
rect 105754 73312 105796 73352
rect 105836 73312 105878 73352
rect 105918 73312 105960 73352
rect 106000 73312 106009 73352
rect 120743 73312 120752 73352
rect 120792 73312 120834 73352
rect 120874 73312 120916 73352
rect 120956 73312 120998 73352
rect 121038 73312 121080 73352
rect 121120 73312 121129 73352
rect 135863 73312 135872 73352
rect 135912 73312 135954 73352
rect 135994 73312 136036 73352
rect 136076 73312 136118 73352
rect 136158 73312 136200 73352
rect 136240 73312 136249 73352
rect 150983 73312 150992 73352
rect 151032 73312 151074 73352
rect 151114 73312 151156 73352
rect 151196 73312 151238 73352
rect 151278 73312 151320 73352
rect 151360 73312 151369 73352
rect 74143 72556 74152 72596
rect 74192 72556 74234 72596
rect 74274 72556 74316 72596
rect 74356 72556 74398 72596
rect 74438 72556 74480 72596
rect 74520 72556 74529 72596
rect 89263 72556 89272 72596
rect 89312 72556 89354 72596
rect 89394 72556 89436 72596
rect 89476 72556 89518 72596
rect 89558 72556 89600 72596
rect 89640 72556 89649 72596
rect 104383 72556 104392 72596
rect 104432 72556 104474 72596
rect 104514 72556 104556 72596
rect 104596 72556 104638 72596
rect 104678 72556 104720 72596
rect 104760 72556 104769 72596
rect 119503 72556 119512 72596
rect 119552 72556 119594 72596
rect 119634 72556 119676 72596
rect 119716 72556 119758 72596
rect 119798 72556 119840 72596
rect 119880 72556 119889 72596
rect 134623 72556 134632 72596
rect 134672 72556 134714 72596
rect 134754 72556 134796 72596
rect 134836 72556 134878 72596
rect 134918 72556 134960 72596
rect 135000 72556 135009 72596
rect 149743 72556 149752 72596
rect 149792 72556 149834 72596
rect 149874 72556 149916 72596
rect 149956 72556 149998 72596
rect 150038 72556 150080 72596
rect 150120 72556 150129 72596
rect 64099 71968 64108 72008
rect 64148 71968 160032 72008
rect 75383 71800 75392 71840
rect 75432 71800 75474 71840
rect 75514 71800 75556 71840
rect 75596 71800 75638 71840
rect 75678 71800 75720 71840
rect 75760 71800 75769 71840
rect 90503 71800 90512 71840
rect 90552 71800 90594 71840
rect 90634 71800 90676 71840
rect 90716 71800 90758 71840
rect 90798 71800 90840 71840
rect 90880 71800 90889 71840
rect 105623 71800 105632 71840
rect 105672 71800 105714 71840
rect 105754 71800 105796 71840
rect 105836 71800 105878 71840
rect 105918 71800 105960 71840
rect 106000 71800 106009 71840
rect 120743 71800 120752 71840
rect 120792 71800 120834 71840
rect 120874 71800 120916 71840
rect 120956 71800 120998 71840
rect 121038 71800 121080 71840
rect 121120 71800 121129 71840
rect 135863 71800 135872 71840
rect 135912 71800 135954 71840
rect 135994 71800 136036 71840
rect 136076 71800 136118 71840
rect 136158 71800 136200 71840
rect 136240 71800 136249 71840
rect 150983 71800 150992 71840
rect 151032 71800 151074 71840
rect 151114 71800 151156 71840
rect 151196 71800 151238 71840
rect 151278 71800 151320 71840
rect 151360 71800 151369 71840
rect 119980 64156 151564 64196
rect 151604 64156 151613 64196
rect 119980 63971 120020 64156
<< via3 >>
rect 75392 151936 75432 151976
rect 75474 151936 75514 151976
rect 75556 151936 75596 151976
rect 75638 151936 75678 151976
rect 75720 151936 75760 151976
rect 90512 151936 90552 151976
rect 90594 151936 90634 151976
rect 90676 151936 90716 151976
rect 90758 151936 90798 151976
rect 90840 151936 90880 151976
rect 105632 151936 105672 151976
rect 105714 151936 105754 151976
rect 105796 151936 105836 151976
rect 105878 151936 105918 151976
rect 105960 151936 106000 151976
rect 120752 151936 120792 151976
rect 120834 151936 120874 151976
rect 120916 151936 120956 151976
rect 120998 151936 121038 151976
rect 121080 151936 121120 151976
rect 135872 151936 135912 151976
rect 135954 151936 135994 151976
rect 136036 151936 136076 151976
rect 136118 151936 136158 151976
rect 136200 151936 136240 151976
rect 150992 151936 151032 151976
rect 151074 151936 151114 151976
rect 151156 151936 151196 151976
rect 151238 151936 151278 151976
rect 151320 151936 151360 151976
rect 74152 151180 74192 151220
rect 74234 151180 74274 151220
rect 74316 151180 74356 151220
rect 74398 151180 74438 151220
rect 74480 151180 74520 151220
rect 89272 151180 89312 151220
rect 89354 151180 89394 151220
rect 89436 151180 89476 151220
rect 89518 151180 89558 151220
rect 89600 151180 89640 151220
rect 104392 151180 104432 151220
rect 104474 151180 104514 151220
rect 104556 151180 104596 151220
rect 104638 151180 104678 151220
rect 104720 151180 104760 151220
rect 119512 151180 119552 151220
rect 119594 151180 119634 151220
rect 119676 151180 119716 151220
rect 119758 151180 119798 151220
rect 119840 151180 119880 151220
rect 134632 151180 134672 151220
rect 134714 151180 134754 151220
rect 134796 151180 134836 151220
rect 134878 151180 134918 151220
rect 134960 151180 135000 151220
rect 149752 151180 149792 151220
rect 149834 151180 149874 151220
rect 149916 151180 149956 151220
rect 149998 151180 150038 151220
rect 150080 151180 150120 151220
rect 75392 150424 75432 150464
rect 75474 150424 75514 150464
rect 75556 150424 75596 150464
rect 75638 150424 75678 150464
rect 75720 150424 75760 150464
rect 90512 150424 90552 150464
rect 90594 150424 90634 150464
rect 90676 150424 90716 150464
rect 90758 150424 90798 150464
rect 90840 150424 90880 150464
rect 105632 150424 105672 150464
rect 105714 150424 105754 150464
rect 105796 150424 105836 150464
rect 105878 150424 105918 150464
rect 105960 150424 106000 150464
rect 120752 150424 120792 150464
rect 120834 150424 120874 150464
rect 120916 150424 120956 150464
rect 120998 150424 121038 150464
rect 121080 150424 121120 150464
rect 135872 150424 135912 150464
rect 135954 150424 135994 150464
rect 136036 150424 136076 150464
rect 136118 150424 136158 150464
rect 136200 150424 136240 150464
rect 150992 150424 151032 150464
rect 151074 150424 151114 150464
rect 151156 150424 151196 150464
rect 151238 150424 151278 150464
rect 151320 150424 151360 150464
rect 74152 149668 74192 149708
rect 74234 149668 74274 149708
rect 74316 149668 74356 149708
rect 74398 149668 74438 149708
rect 74480 149668 74520 149708
rect 89272 149668 89312 149708
rect 89354 149668 89394 149708
rect 89436 149668 89476 149708
rect 89518 149668 89558 149708
rect 89600 149668 89640 149708
rect 104392 149668 104432 149708
rect 104474 149668 104514 149708
rect 104556 149668 104596 149708
rect 104638 149668 104678 149708
rect 104720 149668 104760 149708
rect 119512 149668 119552 149708
rect 119594 149668 119634 149708
rect 119676 149668 119716 149708
rect 119758 149668 119798 149708
rect 119840 149668 119880 149708
rect 134632 149668 134672 149708
rect 134714 149668 134754 149708
rect 134796 149668 134836 149708
rect 134878 149668 134918 149708
rect 134960 149668 135000 149708
rect 149752 149668 149792 149708
rect 149834 149668 149874 149708
rect 149916 149668 149956 149708
rect 149998 149668 150038 149708
rect 150080 149668 150120 149708
rect 75392 148912 75432 148952
rect 75474 148912 75514 148952
rect 75556 148912 75596 148952
rect 75638 148912 75678 148952
rect 75720 148912 75760 148952
rect 90512 148912 90552 148952
rect 90594 148912 90634 148952
rect 90676 148912 90716 148952
rect 90758 148912 90798 148952
rect 90840 148912 90880 148952
rect 105632 148912 105672 148952
rect 105714 148912 105754 148952
rect 105796 148912 105836 148952
rect 105878 148912 105918 148952
rect 105960 148912 106000 148952
rect 120752 148912 120792 148952
rect 120834 148912 120874 148952
rect 120916 148912 120956 148952
rect 120998 148912 121038 148952
rect 121080 148912 121120 148952
rect 135872 148912 135912 148952
rect 135954 148912 135994 148952
rect 136036 148912 136076 148952
rect 136118 148912 136158 148952
rect 136200 148912 136240 148952
rect 150992 148912 151032 148952
rect 151074 148912 151114 148952
rect 151156 148912 151196 148952
rect 151238 148912 151278 148952
rect 151320 148912 151360 148952
rect 74152 148156 74192 148196
rect 74234 148156 74274 148196
rect 74316 148156 74356 148196
rect 74398 148156 74438 148196
rect 74480 148156 74520 148196
rect 89272 148156 89312 148196
rect 89354 148156 89394 148196
rect 89436 148156 89476 148196
rect 89518 148156 89558 148196
rect 89600 148156 89640 148196
rect 104392 148156 104432 148196
rect 104474 148156 104514 148196
rect 104556 148156 104596 148196
rect 104638 148156 104678 148196
rect 104720 148156 104760 148196
rect 119512 148156 119552 148196
rect 119594 148156 119634 148196
rect 119676 148156 119716 148196
rect 119758 148156 119798 148196
rect 119840 148156 119880 148196
rect 134632 148156 134672 148196
rect 134714 148156 134754 148196
rect 134796 148156 134836 148196
rect 134878 148156 134918 148196
rect 134960 148156 135000 148196
rect 149752 148156 149792 148196
rect 149834 148156 149874 148196
rect 149916 148156 149956 148196
rect 149998 148156 150038 148196
rect 150080 148156 150120 148196
rect 75392 147400 75432 147440
rect 75474 147400 75514 147440
rect 75556 147400 75596 147440
rect 75638 147400 75678 147440
rect 75720 147400 75760 147440
rect 90512 147400 90552 147440
rect 90594 147400 90634 147440
rect 90676 147400 90716 147440
rect 90758 147400 90798 147440
rect 90840 147400 90880 147440
rect 105632 147400 105672 147440
rect 105714 147400 105754 147440
rect 105796 147400 105836 147440
rect 105878 147400 105918 147440
rect 105960 147400 106000 147440
rect 120752 147400 120792 147440
rect 120834 147400 120874 147440
rect 120916 147400 120956 147440
rect 120998 147400 121038 147440
rect 121080 147400 121120 147440
rect 135872 147400 135912 147440
rect 135954 147400 135994 147440
rect 136036 147400 136076 147440
rect 136118 147400 136158 147440
rect 136200 147400 136240 147440
rect 150992 147400 151032 147440
rect 151074 147400 151114 147440
rect 151156 147400 151196 147440
rect 151238 147400 151278 147440
rect 151320 147400 151360 147440
rect 74152 146644 74192 146684
rect 74234 146644 74274 146684
rect 74316 146644 74356 146684
rect 74398 146644 74438 146684
rect 74480 146644 74520 146684
rect 89272 146644 89312 146684
rect 89354 146644 89394 146684
rect 89436 146644 89476 146684
rect 89518 146644 89558 146684
rect 89600 146644 89640 146684
rect 104392 146644 104432 146684
rect 104474 146644 104514 146684
rect 104556 146644 104596 146684
rect 104638 146644 104678 146684
rect 104720 146644 104760 146684
rect 119512 146644 119552 146684
rect 119594 146644 119634 146684
rect 119676 146644 119716 146684
rect 119758 146644 119798 146684
rect 119840 146644 119880 146684
rect 134632 146644 134672 146684
rect 134714 146644 134754 146684
rect 134796 146644 134836 146684
rect 134878 146644 134918 146684
rect 134960 146644 135000 146684
rect 149752 146644 149792 146684
rect 149834 146644 149874 146684
rect 149916 146644 149956 146684
rect 149998 146644 150038 146684
rect 150080 146644 150120 146684
rect 75392 145888 75432 145928
rect 75474 145888 75514 145928
rect 75556 145888 75596 145928
rect 75638 145888 75678 145928
rect 75720 145888 75760 145928
rect 90512 145888 90552 145928
rect 90594 145888 90634 145928
rect 90676 145888 90716 145928
rect 90758 145888 90798 145928
rect 90840 145888 90880 145928
rect 105632 145888 105672 145928
rect 105714 145888 105754 145928
rect 105796 145888 105836 145928
rect 105878 145888 105918 145928
rect 105960 145888 106000 145928
rect 120752 145888 120792 145928
rect 120834 145888 120874 145928
rect 120916 145888 120956 145928
rect 120998 145888 121038 145928
rect 121080 145888 121120 145928
rect 135872 145888 135912 145928
rect 135954 145888 135994 145928
rect 136036 145888 136076 145928
rect 136118 145888 136158 145928
rect 136200 145888 136240 145928
rect 150992 145888 151032 145928
rect 151074 145888 151114 145928
rect 151156 145888 151196 145928
rect 151238 145888 151278 145928
rect 151320 145888 151360 145928
rect 74152 145132 74192 145172
rect 74234 145132 74274 145172
rect 74316 145132 74356 145172
rect 74398 145132 74438 145172
rect 74480 145132 74520 145172
rect 89272 145132 89312 145172
rect 89354 145132 89394 145172
rect 89436 145132 89476 145172
rect 89518 145132 89558 145172
rect 89600 145132 89640 145172
rect 104392 145132 104432 145172
rect 104474 145132 104514 145172
rect 104556 145132 104596 145172
rect 104638 145132 104678 145172
rect 104720 145132 104760 145172
rect 119512 145132 119552 145172
rect 119594 145132 119634 145172
rect 119676 145132 119716 145172
rect 119758 145132 119798 145172
rect 119840 145132 119880 145172
rect 134632 145132 134672 145172
rect 134714 145132 134754 145172
rect 134796 145132 134836 145172
rect 134878 145132 134918 145172
rect 134960 145132 135000 145172
rect 149752 145132 149792 145172
rect 149834 145132 149874 145172
rect 149916 145132 149956 145172
rect 149998 145132 150038 145172
rect 150080 145132 150120 145172
rect 75392 144376 75432 144416
rect 75474 144376 75514 144416
rect 75556 144376 75596 144416
rect 75638 144376 75678 144416
rect 75720 144376 75760 144416
rect 90512 144376 90552 144416
rect 90594 144376 90634 144416
rect 90676 144376 90716 144416
rect 90758 144376 90798 144416
rect 90840 144376 90880 144416
rect 105632 144376 105672 144416
rect 105714 144376 105754 144416
rect 105796 144376 105836 144416
rect 105878 144376 105918 144416
rect 105960 144376 106000 144416
rect 120752 144376 120792 144416
rect 120834 144376 120874 144416
rect 120916 144376 120956 144416
rect 120998 144376 121038 144416
rect 121080 144376 121120 144416
rect 135872 144376 135912 144416
rect 135954 144376 135994 144416
rect 136036 144376 136076 144416
rect 136118 144376 136158 144416
rect 136200 144376 136240 144416
rect 150992 144376 151032 144416
rect 151074 144376 151114 144416
rect 151156 144376 151196 144416
rect 151238 144376 151278 144416
rect 151320 144376 151360 144416
rect 74152 143620 74192 143660
rect 74234 143620 74274 143660
rect 74316 143620 74356 143660
rect 74398 143620 74438 143660
rect 74480 143620 74520 143660
rect 89272 143620 89312 143660
rect 89354 143620 89394 143660
rect 89436 143620 89476 143660
rect 89518 143620 89558 143660
rect 89600 143620 89640 143660
rect 104392 143620 104432 143660
rect 104474 143620 104514 143660
rect 104556 143620 104596 143660
rect 104638 143620 104678 143660
rect 104720 143620 104760 143660
rect 119512 143620 119552 143660
rect 119594 143620 119634 143660
rect 119676 143620 119716 143660
rect 119758 143620 119798 143660
rect 119840 143620 119880 143660
rect 134632 143620 134672 143660
rect 134714 143620 134754 143660
rect 134796 143620 134836 143660
rect 134878 143620 134918 143660
rect 134960 143620 135000 143660
rect 149752 143620 149792 143660
rect 149834 143620 149874 143660
rect 149916 143620 149956 143660
rect 149998 143620 150038 143660
rect 150080 143620 150120 143660
rect 75392 142864 75432 142904
rect 75474 142864 75514 142904
rect 75556 142864 75596 142904
rect 75638 142864 75678 142904
rect 75720 142864 75760 142904
rect 90512 142864 90552 142904
rect 90594 142864 90634 142904
rect 90676 142864 90716 142904
rect 90758 142864 90798 142904
rect 90840 142864 90880 142904
rect 105632 142864 105672 142904
rect 105714 142864 105754 142904
rect 105796 142864 105836 142904
rect 105878 142864 105918 142904
rect 105960 142864 106000 142904
rect 120752 142864 120792 142904
rect 120834 142864 120874 142904
rect 120916 142864 120956 142904
rect 120998 142864 121038 142904
rect 121080 142864 121120 142904
rect 135872 142864 135912 142904
rect 135954 142864 135994 142904
rect 136036 142864 136076 142904
rect 136118 142864 136158 142904
rect 136200 142864 136240 142904
rect 150992 142864 151032 142904
rect 151074 142864 151114 142904
rect 151156 142864 151196 142904
rect 151238 142864 151278 142904
rect 151320 142864 151360 142904
rect 74152 142108 74192 142148
rect 74234 142108 74274 142148
rect 74316 142108 74356 142148
rect 74398 142108 74438 142148
rect 74480 142108 74520 142148
rect 89272 142108 89312 142148
rect 89354 142108 89394 142148
rect 89436 142108 89476 142148
rect 89518 142108 89558 142148
rect 89600 142108 89640 142148
rect 104392 142108 104432 142148
rect 104474 142108 104514 142148
rect 104556 142108 104596 142148
rect 104638 142108 104678 142148
rect 104720 142108 104760 142148
rect 119512 142108 119552 142148
rect 119594 142108 119634 142148
rect 119676 142108 119716 142148
rect 119758 142108 119798 142148
rect 119840 142108 119880 142148
rect 134632 142108 134672 142148
rect 134714 142108 134754 142148
rect 134796 142108 134836 142148
rect 134878 142108 134918 142148
rect 134960 142108 135000 142148
rect 149752 142108 149792 142148
rect 149834 142108 149874 142148
rect 149916 142108 149956 142148
rect 149998 142108 150038 142148
rect 150080 142108 150120 142148
rect 75392 141352 75432 141392
rect 75474 141352 75514 141392
rect 75556 141352 75596 141392
rect 75638 141352 75678 141392
rect 75720 141352 75760 141392
rect 90512 141352 90552 141392
rect 90594 141352 90634 141392
rect 90676 141352 90716 141392
rect 90758 141352 90798 141392
rect 90840 141352 90880 141392
rect 105632 141352 105672 141392
rect 105714 141352 105754 141392
rect 105796 141352 105836 141392
rect 105878 141352 105918 141392
rect 105960 141352 106000 141392
rect 120752 141352 120792 141392
rect 120834 141352 120874 141392
rect 120916 141352 120956 141392
rect 120998 141352 121038 141392
rect 121080 141352 121120 141392
rect 135872 141352 135912 141392
rect 135954 141352 135994 141392
rect 136036 141352 136076 141392
rect 136118 141352 136158 141392
rect 136200 141352 136240 141392
rect 150992 141352 151032 141392
rect 151074 141352 151114 141392
rect 151156 141352 151196 141392
rect 151238 141352 151278 141392
rect 151320 141352 151360 141392
rect 74152 140596 74192 140636
rect 74234 140596 74274 140636
rect 74316 140596 74356 140636
rect 74398 140596 74438 140636
rect 74480 140596 74520 140636
rect 89272 140596 89312 140636
rect 89354 140596 89394 140636
rect 89436 140596 89476 140636
rect 89518 140596 89558 140636
rect 89600 140596 89640 140636
rect 104392 140596 104432 140636
rect 104474 140596 104514 140636
rect 104556 140596 104596 140636
rect 104638 140596 104678 140636
rect 104720 140596 104760 140636
rect 119512 140596 119552 140636
rect 119594 140596 119634 140636
rect 119676 140596 119716 140636
rect 119758 140596 119798 140636
rect 119840 140596 119880 140636
rect 134632 140596 134672 140636
rect 134714 140596 134754 140636
rect 134796 140596 134836 140636
rect 134878 140596 134918 140636
rect 134960 140596 135000 140636
rect 149752 140596 149792 140636
rect 149834 140596 149874 140636
rect 149916 140596 149956 140636
rect 149998 140596 150038 140636
rect 150080 140596 150120 140636
rect 75392 139840 75432 139880
rect 75474 139840 75514 139880
rect 75556 139840 75596 139880
rect 75638 139840 75678 139880
rect 75720 139840 75760 139880
rect 90512 139840 90552 139880
rect 90594 139840 90634 139880
rect 90676 139840 90716 139880
rect 90758 139840 90798 139880
rect 90840 139840 90880 139880
rect 105632 139840 105672 139880
rect 105714 139840 105754 139880
rect 105796 139840 105836 139880
rect 105878 139840 105918 139880
rect 105960 139840 106000 139880
rect 120752 139840 120792 139880
rect 120834 139840 120874 139880
rect 120916 139840 120956 139880
rect 120998 139840 121038 139880
rect 121080 139840 121120 139880
rect 135872 139840 135912 139880
rect 135954 139840 135994 139880
rect 136036 139840 136076 139880
rect 136118 139840 136158 139880
rect 136200 139840 136240 139880
rect 150992 139840 151032 139880
rect 151074 139840 151114 139880
rect 151156 139840 151196 139880
rect 151238 139840 151278 139880
rect 151320 139840 151360 139880
rect 74152 139084 74192 139124
rect 74234 139084 74274 139124
rect 74316 139084 74356 139124
rect 74398 139084 74438 139124
rect 74480 139084 74520 139124
rect 89272 139084 89312 139124
rect 89354 139084 89394 139124
rect 89436 139084 89476 139124
rect 89518 139084 89558 139124
rect 89600 139084 89640 139124
rect 104392 139084 104432 139124
rect 104474 139084 104514 139124
rect 104556 139084 104596 139124
rect 104638 139084 104678 139124
rect 104720 139084 104760 139124
rect 119512 139084 119552 139124
rect 119594 139084 119634 139124
rect 119676 139084 119716 139124
rect 119758 139084 119798 139124
rect 119840 139084 119880 139124
rect 134632 139084 134672 139124
rect 134714 139084 134754 139124
rect 134796 139084 134836 139124
rect 134878 139084 134918 139124
rect 134960 139084 135000 139124
rect 149752 139084 149792 139124
rect 149834 139084 149874 139124
rect 149916 139084 149956 139124
rect 149998 139084 150038 139124
rect 150080 139084 150120 139124
rect 75392 138328 75432 138368
rect 75474 138328 75514 138368
rect 75556 138328 75596 138368
rect 75638 138328 75678 138368
rect 75720 138328 75760 138368
rect 90512 138328 90552 138368
rect 90594 138328 90634 138368
rect 90676 138328 90716 138368
rect 90758 138328 90798 138368
rect 90840 138328 90880 138368
rect 105632 138328 105672 138368
rect 105714 138328 105754 138368
rect 105796 138328 105836 138368
rect 105878 138328 105918 138368
rect 105960 138328 106000 138368
rect 120752 138328 120792 138368
rect 120834 138328 120874 138368
rect 120916 138328 120956 138368
rect 120998 138328 121038 138368
rect 121080 138328 121120 138368
rect 135872 138328 135912 138368
rect 135954 138328 135994 138368
rect 136036 138328 136076 138368
rect 136118 138328 136158 138368
rect 136200 138328 136240 138368
rect 150992 138328 151032 138368
rect 151074 138328 151114 138368
rect 151156 138328 151196 138368
rect 151238 138328 151278 138368
rect 151320 138328 151360 138368
rect 74152 137572 74192 137612
rect 74234 137572 74274 137612
rect 74316 137572 74356 137612
rect 74398 137572 74438 137612
rect 74480 137572 74520 137612
rect 89272 137572 89312 137612
rect 89354 137572 89394 137612
rect 89436 137572 89476 137612
rect 89518 137572 89558 137612
rect 89600 137572 89640 137612
rect 104392 137572 104432 137612
rect 104474 137572 104514 137612
rect 104556 137572 104596 137612
rect 104638 137572 104678 137612
rect 104720 137572 104760 137612
rect 119512 137572 119552 137612
rect 119594 137572 119634 137612
rect 119676 137572 119716 137612
rect 119758 137572 119798 137612
rect 119840 137572 119880 137612
rect 134632 137572 134672 137612
rect 134714 137572 134754 137612
rect 134796 137572 134836 137612
rect 134878 137572 134918 137612
rect 134960 137572 135000 137612
rect 149752 137572 149792 137612
rect 149834 137572 149874 137612
rect 149916 137572 149956 137612
rect 149998 137572 150038 137612
rect 150080 137572 150120 137612
rect 75392 136816 75432 136856
rect 75474 136816 75514 136856
rect 75556 136816 75596 136856
rect 75638 136816 75678 136856
rect 75720 136816 75760 136856
rect 90512 136816 90552 136856
rect 90594 136816 90634 136856
rect 90676 136816 90716 136856
rect 90758 136816 90798 136856
rect 90840 136816 90880 136856
rect 105632 136816 105672 136856
rect 105714 136816 105754 136856
rect 105796 136816 105836 136856
rect 105878 136816 105918 136856
rect 105960 136816 106000 136856
rect 120752 136816 120792 136856
rect 120834 136816 120874 136856
rect 120916 136816 120956 136856
rect 120998 136816 121038 136856
rect 121080 136816 121120 136856
rect 135872 136816 135912 136856
rect 135954 136816 135994 136856
rect 136036 136816 136076 136856
rect 136118 136816 136158 136856
rect 136200 136816 136240 136856
rect 150992 136816 151032 136856
rect 151074 136816 151114 136856
rect 151156 136816 151196 136856
rect 151238 136816 151278 136856
rect 151320 136816 151360 136856
rect 74152 136060 74192 136100
rect 74234 136060 74274 136100
rect 74316 136060 74356 136100
rect 74398 136060 74438 136100
rect 74480 136060 74520 136100
rect 89272 136060 89312 136100
rect 89354 136060 89394 136100
rect 89436 136060 89476 136100
rect 89518 136060 89558 136100
rect 89600 136060 89640 136100
rect 104392 136060 104432 136100
rect 104474 136060 104514 136100
rect 104556 136060 104596 136100
rect 104638 136060 104678 136100
rect 104720 136060 104760 136100
rect 119512 136060 119552 136100
rect 119594 136060 119634 136100
rect 119676 136060 119716 136100
rect 119758 136060 119798 136100
rect 119840 136060 119880 136100
rect 134632 136060 134672 136100
rect 134714 136060 134754 136100
rect 134796 136060 134836 136100
rect 134878 136060 134918 136100
rect 134960 136060 135000 136100
rect 149752 136060 149792 136100
rect 149834 136060 149874 136100
rect 149916 136060 149956 136100
rect 149998 136060 150038 136100
rect 150080 136060 150120 136100
rect 75392 135304 75432 135344
rect 75474 135304 75514 135344
rect 75556 135304 75596 135344
rect 75638 135304 75678 135344
rect 75720 135304 75760 135344
rect 90512 135304 90552 135344
rect 90594 135304 90634 135344
rect 90676 135304 90716 135344
rect 90758 135304 90798 135344
rect 90840 135304 90880 135344
rect 105632 135304 105672 135344
rect 105714 135304 105754 135344
rect 105796 135304 105836 135344
rect 105878 135304 105918 135344
rect 105960 135304 106000 135344
rect 120752 135304 120792 135344
rect 120834 135304 120874 135344
rect 120916 135304 120956 135344
rect 120998 135304 121038 135344
rect 121080 135304 121120 135344
rect 135872 135304 135912 135344
rect 135954 135304 135994 135344
rect 136036 135304 136076 135344
rect 136118 135304 136158 135344
rect 136200 135304 136240 135344
rect 150992 135304 151032 135344
rect 151074 135304 151114 135344
rect 151156 135304 151196 135344
rect 151238 135304 151278 135344
rect 151320 135304 151360 135344
rect 74152 134548 74192 134588
rect 74234 134548 74274 134588
rect 74316 134548 74356 134588
rect 74398 134548 74438 134588
rect 74480 134548 74520 134588
rect 89272 134548 89312 134588
rect 89354 134548 89394 134588
rect 89436 134548 89476 134588
rect 89518 134548 89558 134588
rect 89600 134548 89640 134588
rect 104392 134548 104432 134588
rect 104474 134548 104514 134588
rect 104556 134548 104596 134588
rect 104638 134548 104678 134588
rect 104720 134548 104760 134588
rect 119512 134548 119552 134588
rect 119594 134548 119634 134588
rect 119676 134548 119716 134588
rect 119758 134548 119798 134588
rect 119840 134548 119880 134588
rect 134632 134548 134672 134588
rect 134714 134548 134754 134588
rect 134796 134548 134836 134588
rect 134878 134548 134918 134588
rect 134960 134548 135000 134588
rect 149752 134548 149792 134588
rect 149834 134548 149874 134588
rect 149916 134548 149956 134588
rect 149998 134548 150038 134588
rect 150080 134548 150120 134588
rect 75392 133792 75432 133832
rect 75474 133792 75514 133832
rect 75556 133792 75596 133832
rect 75638 133792 75678 133832
rect 75720 133792 75760 133832
rect 90512 133792 90552 133832
rect 90594 133792 90634 133832
rect 90676 133792 90716 133832
rect 90758 133792 90798 133832
rect 90840 133792 90880 133832
rect 105632 133792 105672 133832
rect 105714 133792 105754 133832
rect 105796 133792 105836 133832
rect 105878 133792 105918 133832
rect 105960 133792 106000 133832
rect 120752 133792 120792 133832
rect 120834 133792 120874 133832
rect 120916 133792 120956 133832
rect 120998 133792 121038 133832
rect 121080 133792 121120 133832
rect 135872 133792 135912 133832
rect 135954 133792 135994 133832
rect 136036 133792 136076 133832
rect 136118 133792 136158 133832
rect 136200 133792 136240 133832
rect 150992 133792 151032 133832
rect 151074 133792 151114 133832
rect 151156 133792 151196 133832
rect 151238 133792 151278 133832
rect 151320 133792 151360 133832
rect 74152 133036 74192 133076
rect 74234 133036 74274 133076
rect 74316 133036 74356 133076
rect 74398 133036 74438 133076
rect 74480 133036 74520 133076
rect 89272 133036 89312 133076
rect 89354 133036 89394 133076
rect 89436 133036 89476 133076
rect 89518 133036 89558 133076
rect 89600 133036 89640 133076
rect 104392 133036 104432 133076
rect 104474 133036 104514 133076
rect 104556 133036 104596 133076
rect 104638 133036 104678 133076
rect 104720 133036 104760 133076
rect 119512 133036 119552 133076
rect 119594 133036 119634 133076
rect 119676 133036 119716 133076
rect 119758 133036 119798 133076
rect 119840 133036 119880 133076
rect 134632 133036 134672 133076
rect 134714 133036 134754 133076
rect 134796 133036 134836 133076
rect 134878 133036 134918 133076
rect 134960 133036 135000 133076
rect 149752 133036 149792 133076
rect 149834 133036 149874 133076
rect 149916 133036 149956 133076
rect 149998 133036 150038 133076
rect 150080 133036 150120 133076
rect 75392 132280 75432 132320
rect 75474 132280 75514 132320
rect 75556 132280 75596 132320
rect 75638 132280 75678 132320
rect 75720 132280 75760 132320
rect 90512 132280 90552 132320
rect 90594 132280 90634 132320
rect 90676 132280 90716 132320
rect 90758 132280 90798 132320
rect 90840 132280 90880 132320
rect 105632 132280 105672 132320
rect 105714 132280 105754 132320
rect 105796 132280 105836 132320
rect 105878 132280 105918 132320
rect 105960 132280 106000 132320
rect 120752 132280 120792 132320
rect 120834 132280 120874 132320
rect 120916 132280 120956 132320
rect 120998 132280 121038 132320
rect 121080 132280 121120 132320
rect 135872 132280 135912 132320
rect 135954 132280 135994 132320
rect 136036 132280 136076 132320
rect 136118 132280 136158 132320
rect 136200 132280 136240 132320
rect 150992 132280 151032 132320
rect 151074 132280 151114 132320
rect 151156 132280 151196 132320
rect 151238 132280 151278 132320
rect 151320 132280 151360 132320
rect 74152 131524 74192 131564
rect 74234 131524 74274 131564
rect 74316 131524 74356 131564
rect 74398 131524 74438 131564
rect 74480 131524 74520 131564
rect 89272 131524 89312 131564
rect 89354 131524 89394 131564
rect 89436 131524 89476 131564
rect 89518 131524 89558 131564
rect 89600 131524 89640 131564
rect 104392 131524 104432 131564
rect 104474 131524 104514 131564
rect 104556 131524 104596 131564
rect 104638 131524 104678 131564
rect 104720 131524 104760 131564
rect 119512 131524 119552 131564
rect 119594 131524 119634 131564
rect 119676 131524 119716 131564
rect 119758 131524 119798 131564
rect 119840 131524 119880 131564
rect 134632 131524 134672 131564
rect 134714 131524 134754 131564
rect 134796 131524 134836 131564
rect 134878 131524 134918 131564
rect 134960 131524 135000 131564
rect 149752 131524 149792 131564
rect 149834 131524 149874 131564
rect 149916 131524 149956 131564
rect 149998 131524 150038 131564
rect 150080 131524 150120 131564
rect 75392 130768 75432 130808
rect 75474 130768 75514 130808
rect 75556 130768 75596 130808
rect 75638 130768 75678 130808
rect 75720 130768 75760 130808
rect 90512 130768 90552 130808
rect 90594 130768 90634 130808
rect 90676 130768 90716 130808
rect 90758 130768 90798 130808
rect 90840 130768 90880 130808
rect 105632 130768 105672 130808
rect 105714 130768 105754 130808
rect 105796 130768 105836 130808
rect 105878 130768 105918 130808
rect 105960 130768 106000 130808
rect 120752 130768 120792 130808
rect 120834 130768 120874 130808
rect 120916 130768 120956 130808
rect 120998 130768 121038 130808
rect 121080 130768 121120 130808
rect 135872 130768 135912 130808
rect 135954 130768 135994 130808
rect 136036 130768 136076 130808
rect 136118 130768 136158 130808
rect 136200 130768 136240 130808
rect 150992 130768 151032 130808
rect 151074 130768 151114 130808
rect 151156 130768 151196 130808
rect 151238 130768 151278 130808
rect 151320 130768 151360 130808
rect 74152 130012 74192 130052
rect 74234 130012 74274 130052
rect 74316 130012 74356 130052
rect 74398 130012 74438 130052
rect 74480 130012 74520 130052
rect 89272 130012 89312 130052
rect 89354 130012 89394 130052
rect 89436 130012 89476 130052
rect 89518 130012 89558 130052
rect 89600 130012 89640 130052
rect 104392 130012 104432 130052
rect 104474 130012 104514 130052
rect 104556 130012 104596 130052
rect 104638 130012 104678 130052
rect 104720 130012 104760 130052
rect 119512 130012 119552 130052
rect 119594 130012 119634 130052
rect 119676 130012 119716 130052
rect 119758 130012 119798 130052
rect 119840 130012 119880 130052
rect 134632 130012 134672 130052
rect 134714 130012 134754 130052
rect 134796 130012 134836 130052
rect 134878 130012 134918 130052
rect 134960 130012 135000 130052
rect 149752 130012 149792 130052
rect 149834 130012 149874 130052
rect 149916 130012 149956 130052
rect 149998 130012 150038 130052
rect 150080 130012 150120 130052
rect 75392 129256 75432 129296
rect 75474 129256 75514 129296
rect 75556 129256 75596 129296
rect 75638 129256 75678 129296
rect 75720 129256 75760 129296
rect 90512 129256 90552 129296
rect 90594 129256 90634 129296
rect 90676 129256 90716 129296
rect 90758 129256 90798 129296
rect 90840 129256 90880 129296
rect 105632 129256 105672 129296
rect 105714 129256 105754 129296
rect 105796 129256 105836 129296
rect 105878 129256 105918 129296
rect 105960 129256 106000 129296
rect 120752 129256 120792 129296
rect 120834 129256 120874 129296
rect 120916 129256 120956 129296
rect 120998 129256 121038 129296
rect 121080 129256 121120 129296
rect 135872 129256 135912 129296
rect 135954 129256 135994 129296
rect 136036 129256 136076 129296
rect 136118 129256 136158 129296
rect 136200 129256 136240 129296
rect 150992 129256 151032 129296
rect 151074 129256 151114 129296
rect 151156 129256 151196 129296
rect 151238 129256 151278 129296
rect 151320 129256 151360 129296
rect 74152 128500 74192 128540
rect 74234 128500 74274 128540
rect 74316 128500 74356 128540
rect 74398 128500 74438 128540
rect 74480 128500 74520 128540
rect 89272 128500 89312 128540
rect 89354 128500 89394 128540
rect 89436 128500 89476 128540
rect 89518 128500 89558 128540
rect 89600 128500 89640 128540
rect 104392 128500 104432 128540
rect 104474 128500 104514 128540
rect 104556 128500 104596 128540
rect 104638 128500 104678 128540
rect 104720 128500 104760 128540
rect 119512 128500 119552 128540
rect 119594 128500 119634 128540
rect 119676 128500 119716 128540
rect 119758 128500 119798 128540
rect 119840 128500 119880 128540
rect 134632 128500 134672 128540
rect 134714 128500 134754 128540
rect 134796 128500 134836 128540
rect 134878 128500 134918 128540
rect 134960 128500 135000 128540
rect 149752 128500 149792 128540
rect 149834 128500 149874 128540
rect 149916 128500 149956 128540
rect 149998 128500 150038 128540
rect 150080 128500 150120 128540
rect 75392 127744 75432 127784
rect 75474 127744 75514 127784
rect 75556 127744 75596 127784
rect 75638 127744 75678 127784
rect 75720 127744 75760 127784
rect 90512 127744 90552 127784
rect 90594 127744 90634 127784
rect 90676 127744 90716 127784
rect 90758 127744 90798 127784
rect 90840 127744 90880 127784
rect 105632 127744 105672 127784
rect 105714 127744 105754 127784
rect 105796 127744 105836 127784
rect 105878 127744 105918 127784
rect 105960 127744 106000 127784
rect 120752 127744 120792 127784
rect 120834 127744 120874 127784
rect 120916 127744 120956 127784
rect 120998 127744 121038 127784
rect 121080 127744 121120 127784
rect 135872 127744 135912 127784
rect 135954 127744 135994 127784
rect 136036 127744 136076 127784
rect 136118 127744 136158 127784
rect 136200 127744 136240 127784
rect 150992 127744 151032 127784
rect 151074 127744 151114 127784
rect 151156 127744 151196 127784
rect 151238 127744 151278 127784
rect 151320 127744 151360 127784
rect 74152 126988 74192 127028
rect 74234 126988 74274 127028
rect 74316 126988 74356 127028
rect 74398 126988 74438 127028
rect 74480 126988 74520 127028
rect 89272 126988 89312 127028
rect 89354 126988 89394 127028
rect 89436 126988 89476 127028
rect 89518 126988 89558 127028
rect 89600 126988 89640 127028
rect 104392 126988 104432 127028
rect 104474 126988 104514 127028
rect 104556 126988 104596 127028
rect 104638 126988 104678 127028
rect 104720 126988 104760 127028
rect 119512 126988 119552 127028
rect 119594 126988 119634 127028
rect 119676 126988 119716 127028
rect 119758 126988 119798 127028
rect 119840 126988 119880 127028
rect 134632 126988 134672 127028
rect 134714 126988 134754 127028
rect 134796 126988 134836 127028
rect 134878 126988 134918 127028
rect 134960 126988 135000 127028
rect 149752 126988 149792 127028
rect 149834 126988 149874 127028
rect 149916 126988 149956 127028
rect 149998 126988 150038 127028
rect 150080 126988 150120 127028
rect 75392 126232 75432 126272
rect 75474 126232 75514 126272
rect 75556 126232 75596 126272
rect 75638 126232 75678 126272
rect 75720 126232 75760 126272
rect 90512 126232 90552 126272
rect 90594 126232 90634 126272
rect 90676 126232 90716 126272
rect 90758 126232 90798 126272
rect 90840 126232 90880 126272
rect 105632 126232 105672 126272
rect 105714 126232 105754 126272
rect 105796 126232 105836 126272
rect 105878 126232 105918 126272
rect 105960 126232 106000 126272
rect 120752 126232 120792 126272
rect 120834 126232 120874 126272
rect 120916 126232 120956 126272
rect 120998 126232 121038 126272
rect 121080 126232 121120 126272
rect 135872 126232 135912 126272
rect 135954 126232 135994 126272
rect 136036 126232 136076 126272
rect 136118 126232 136158 126272
rect 136200 126232 136240 126272
rect 150992 126232 151032 126272
rect 151074 126232 151114 126272
rect 151156 126232 151196 126272
rect 151238 126232 151278 126272
rect 151320 126232 151360 126272
rect 74152 125476 74192 125516
rect 74234 125476 74274 125516
rect 74316 125476 74356 125516
rect 74398 125476 74438 125516
rect 74480 125476 74520 125516
rect 89272 125476 89312 125516
rect 89354 125476 89394 125516
rect 89436 125476 89476 125516
rect 89518 125476 89558 125516
rect 89600 125476 89640 125516
rect 104392 125476 104432 125516
rect 104474 125476 104514 125516
rect 104556 125476 104596 125516
rect 104638 125476 104678 125516
rect 104720 125476 104760 125516
rect 119512 125476 119552 125516
rect 119594 125476 119634 125516
rect 119676 125476 119716 125516
rect 119758 125476 119798 125516
rect 119840 125476 119880 125516
rect 134632 125476 134672 125516
rect 134714 125476 134754 125516
rect 134796 125476 134836 125516
rect 134878 125476 134918 125516
rect 134960 125476 135000 125516
rect 149752 125476 149792 125516
rect 149834 125476 149874 125516
rect 149916 125476 149956 125516
rect 149998 125476 150038 125516
rect 150080 125476 150120 125516
rect 75392 124720 75432 124760
rect 75474 124720 75514 124760
rect 75556 124720 75596 124760
rect 75638 124720 75678 124760
rect 75720 124720 75760 124760
rect 90512 124720 90552 124760
rect 90594 124720 90634 124760
rect 90676 124720 90716 124760
rect 90758 124720 90798 124760
rect 90840 124720 90880 124760
rect 105632 124720 105672 124760
rect 105714 124720 105754 124760
rect 105796 124720 105836 124760
rect 105878 124720 105918 124760
rect 105960 124720 106000 124760
rect 120752 124720 120792 124760
rect 120834 124720 120874 124760
rect 120916 124720 120956 124760
rect 120998 124720 121038 124760
rect 121080 124720 121120 124760
rect 135872 124720 135912 124760
rect 135954 124720 135994 124760
rect 136036 124720 136076 124760
rect 136118 124720 136158 124760
rect 136200 124720 136240 124760
rect 150992 124720 151032 124760
rect 151074 124720 151114 124760
rect 151156 124720 151196 124760
rect 151238 124720 151278 124760
rect 151320 124720 151360 124760
rect 74152 123964 74192 124004
rect 74234 123964 74274 124004
rect 74316 123964 74356 124004
rect 74398 123964 74438 124004
rect 74480 123964 74520 124004
rect 89272 123964 89312 124004
rect 89354 123964 89394 124004
rect 89436 123964 89476 124004
rect 89518 123964 89558 124004
rect 89600 123964 89640 124004
rect 104392 123964 104432 124004
rect 104474 123964 104514 124004
rect 104556 123964 104596 124004
rect 104638 123964 104678 124004
rect 104720 123964 104760 124004
rect 119512 123964 119552 124004
rect 119594 123964 119634 124004
rect 119676 123964 119716 124004
rect 119758 123964 119798 124004
rect 119840 123964 119880 124004
rect 134632 123964 134672 124004
rect 134714 123964 134754 124004
rect 134796 123964 134836 124004
rect 134878 123964 134918 124004
rect 134960 123964 135000 124004
rect 149752 123964 149792 124004
rect 149834 123964 149874 124004
rect 149916 123964 149956 124004
rect 149998 123964 150038 124004
rect 150080 123964 150120 124004
rect 75392 123208 75432 123248
rect 75474 123208 75514 123248
rect 75556 123208 75596 123248
rect 75638 123208 75678 123248
rect 75720 123208 75760 123248
rect 90512 123208 90552 123248
rect 90594 123208 90634 123248
rect 90676 123208 90716 123248
rect 90758 123208 90798 123248
rect 90840 123208 90880 123248
rect 105632 123208 105672 123248
rect 105714 123208 105754 123248
rect 105796 123208 105836 123248
rect 105878 123208 105918 123248
rect 105960 123208 106000 123248
rect 120752 123208 120792 123248
rect 120834 123208 120874 123248
rect 120916 123208 120956 123248
rect 120998 123208 121038 123248
rect 121080 123208 121120 123248
rect 135872 123208 135912 123248
rect 135954 123208 135994 123248
rect 136036 123208 136076 123248
rect 136118 123208 136158 123248
rect 136200 123208 136240 123248
rect 150992 123208 151032 123248
rect 151074 123208 151114 123248
rect 151156 123208 151196 123248
rect 151238 123208 151278 123248
rect 151320 123208 151360 123248
rect 74152 122452 74192 122492
rect 74234 122452 74274 122492
rect 74316 122452 74356 122492
rect 74398 122452 74438 122492
rect 74480 122452 74520 122492
rect 89272 122452 89312 122492
rect 89354 122452 89394 122492
rect 89436 122452 89476 122492
rect 89518 122452 89558 122492
rect 89600 122452 89640 122492
rect 104392 122452 104432 122492
rect 104474 122452 104514 122492
rect 104556 122452 104596 122492
rect 104638 122452 104678 122492
rect 104720 122452 104760 122492
rect 119512 122452 119552 122492
rect 119594 122452 119634 122492
rect 119676 122452 119716 122492
rect 119758 122452 119798 122492
rect 119840 122452 119880 122492
rect 134632 122452 134672 122492
rect 134714 122452 134754 122492
rect 134796 122452 134836 122492
rect 134878 122452 134918 122492
rect 134960 122452 135000 122492
rect 149752 122452 149792 122492
rect 149834 122452 149874 122492
rect 149916 122452 149956 122492
rect 149998 122452 150038 122492
rect 150080 122452 150120 122492
rect 75392 121696 75432 121736
rect 75474 121696 75514 121736
rect 75556 121696 75596 121736
rect 75638 121696 75678 121736
rect 75720 121696 75760 121736
rect 90512 121696 90552 121736
rect 90594 121696 90634 121736
rect 90676 121696 90716 121736
rect 90758 121696 90798 121736
rect 90840 121696 90880 121736
rect 105632 121696 105672 121736
rect 105714 121696 105754 121736
rect 105796 121696 105836 121736
rect 105878 121696 105918 121736
rect 105960 121696 106000 121736
rect 120752 121696 120792 121736
rect 120834 121696 120874 121736
rect 120916 121696 120956 121736
rect 120998 121696 121038 121736
rect 121080 121696 121120 121736
rect 135872 121696 135912 121736
rect 135954 121696 135994 121736
rect 136036 121696 136076 121736
rect 136118 121696 136158 121736
rect 136200 121696 136240 121736
rect 150992 121696 151032 121736
rect 151074 121696 151114 121736
rect 151156 121696 151196 121736
rect 151238 121696 151278 121736
rect 151320 121696 151360 121736
rect 74152 120940 74192 120980
rect 74234 120940 74274 120980
rect 74316 120940 74356 120980
rect 74398 120940 74438 120980
rect 74480 120940 74520 120980
rect 89272 120940 89312 120980
rect 89354 120940 89394 120980
rect 89436 120940 89476 120980
rect 89518 120940 89558 120980
rect 89600 120940 89640 120980
rect 104392 120940 104432 120980
rect 104474 120940 104514 120980
rect 104556 120940 104596 120980
rect 104638 120940 104678 120980
rect 104720 120940 104760 120980
rect 119512 120940 119552 120980
rect 119594 120940 119634 120980
rect 119676 120940 119716 120980
rect 119758 120940 119798 120980
rect 119840 120940 119880 120980
rect 134632 120940 134672 120980
rect 134714 120940 134754 120980
rect 134796 120940 134836 120980
rect 134878 120940 134918 120980
rect 134960 120940 135000 120980
rect 149752 120940 149792 120980
rect 149834 120940 149874 120980
rect 149916 120940 149956 120980
rect 149998 120940 150038 120980
rect 150080 120940 150120 120980
rect 75392 120184 75432 120224
rect 75474 120184 75514 120224
rect 75556 120184 75596 120224
rect 75638 120184 75678 120224
rect 75720 120184 75760 120224
rect 90512 120184 90552 120224
rect 90594 120184 90634 120224
rect 90676 120184 90716 120224
rect 90758 120184 90798 120224
rect 90840 120184 90880 120224
rect 105632 120184 105672 120224
rect 105714 120184 105754 120224
rect 105796 120184 105836 120224
rect 105878 120184 105918 120224
rect 105960 120184 106000 120224
rect 120752 120184 120792 120224
rect 120834 120184 120874 120224
rect 120916 120184 120956 120224
rect 120998 120184 121038 120224
rect 121080 120184 121120 120224
rect 135872 120184 135912 120224
rect 135954 120184 135994 120224
rect 136036 120184 136076 120224
rect 136118 120184 136158 120224
rect 136200 120184 136240 120224
rect 150992 120184 151032 120224
rect 151074 120184 151114 120224
rect 151156 120184 151196 120224
rect 151238 120184 151278 120224
rect 151320 120184 151360 120224
rect 74152 119428 74192 119468
rect 74234 119428 74274 119468
rect 74316 119428 74356 119468
rect 74398 119428 74438 119468
rect 74480 119428 74520 119468
rect 89272 119428 89312 119468
rect 89354 119428 89394 119468
rect 89436 119428 89476 119468
rect 89518 119428 89558 119468
rect 89600 119428 89640 119468
rect 104392 119428 104432 119468
rect 104474 119428 104514 119468
rect 104556 119428 104596 119468
rect 104638 119428 104678 119468
rect 104720 119428 104760 119468
rect 119512 119428 119552 119468
rect 119594 119428 119634 119468
rect 119676 119428 119716 119468
rect 119758 119428 119798 119468
rect 119840 119428 119880 119468
rect 134632 119428 134672 119468
rect 134714 119428 134754 119468
rect 134796 119428 134836 119468
rect 134878 119428 134918 119468
rect 134960 119428 135000 119468
rect 149752 119428 149792 119468
rect 149834 119428 149874 119468
rect 149916 119428 149956 119468
rect 149998 119428 150038 119468
rect 150080 119428 150120 119468
rect 75392 118672 75432 118712
rect 75474 118672 75514 118712
rect 75556 118672 75596 118712
rect 75638 118672 75678 118712
rect 75720 118672 75760 118712
rect 90512 118672 90552 118712
rect 90594 118672 90634 118712
rect 90676 118672 90716 118712
rect 90758 118672 90798 118712
rect 90840 118672 90880 118712
rect 105632 118672 105672 118712
rect 105714 118672 105754 118712
rect 105796 118672 105836 118712
rect 105878 118672 105918 118712
rect 105960 118672 106000 118712
rect 120752 118672 120792 118712
rect 120834 118672 120874 118712
rect 120916 118672 120956 118712
rect 120998 118672 121038 118712
rect 121080 118672 121120 118712
rect 135872 118672 135912 118712
rect 135954 118672 135994 118712
rect 136036 118672 136076 118712
rect 136118 118672 136158 118712
rect 136200 118672 136240 118712
rect 150992 118672 151032 118712
rect 151074 118672 151114 118712
rect 151156 118672 151196 118712
rect 151238 118672 151278 118712
rect 151320 118672 151360 118712
rect 74152 117916 74192 117956
rect 74234 117916 74274 117956
rect 74316 117916 74356 117956
rect 74398 117916 74438 117956
rect 74480 117916 74520 117956
rect 89272 117916 89312 117956
rect 89354 117916 89394 117956
rect 89436 117916 89476 117956
rect 89518 117916 89558 117956
rect 89600 117916 89640 117956
rect 104392 117916 104432 117956
rect 104474 117916 104514 117956
rect 104556 117916 104596 117956
rect 104638 117916 104678 117956
rect 104720 117916 104760 117956
rect 119512 117916 119552 117956
rect 119594 117916 119634 117956
rect 119676 117916 119716 117956
rect 119758 117916 119798 117956
rect 119840 117916 119880 117956
rect 134632 117916 134672 117956
rect 134714 117916 134754 117956
rect 134796 117916 134836 117956
rect 134878 117916 134918 117956
rect 134960 117916 135000 117956
rect 149752 117916 149792 117956
rect 149834 117916 149874 117956
rect 149916 117916 149956 117956
rect 149998 117916 150038 117956
rect 150080 117916 150120 117956
rect 75392 117160 75432 117200
rect 75474 117160 75514 117200
rect 75556 117160 75596 117200
rect 75638 117160 75678 117200
rect 75720 117160 75760 117200
rect 90512 117160 90552 117200
rect 90594 117160 90634 117200
rect 90676 117160 90716 117200
rect 90758 117160 90798 117200
rect 90840 117160 90880 117200
rect 105632 117160 105672 117200
rect 105714 117160 105754 117200
rect 105796 117160 105836 117200
rect 105878 117160 105918 117200
rect 105960 117160 106000 117200
rect 120752 117160 120792 117200
rect 120834 117160 120874 117200
rect 120916 117160 120956 117200
rect 120998 117160 121038 117200
rect 121080 117160 121120 117200
rect 135872 117160 135912 117200
rect 135954 117160 135994 117200
rect 136036 117160 136076 117200
rect 136118 117160 136158 117200
rect 136200 117160 136240 117200
rect 150992 117160 151032 117200
rect 151074 117160 151114 117200
rect 151156 117160 151196 117200
rect 151238 117160 151278 117200
rect 151320 117160 151360 117200
rect 74152 116404 74192 116444
rect 74234 116404 74274 116444
rect 74316 116404 74356 116444
rect 74398 116404 74438 116444
rect 74480 116404 74520 116444
rect 89272 116404 89312 116444
rect 89354 116404 89394 116444
rect 89436 116404 89476 116444
rect 89518 116404 89558 116444
rect 89600 116404 89640 116444
rect 104392 116404 104432 116444
rect 104474 116404 104514 116444
rect 104556 116404 104596 116444
rect 104638 116404 104678 116444
rect 104720 116404 104760 116444
rect 119512 116404 119552 116444
rect 119594 116404 119634 116444
rect 119676 116404 119716 116444
rect 119758 116404 119798 116444
rect 119840 116404 119880 116444
rect 134632 116404 134672 116444
rect 134714 116404 134754 116444
rect 134796 116404 134836 116444
rect 134878 116404 134918 116444
rect 134960 116404 135000 116444
rect 149752 116404 149792 116444
rect 149834 116404 149874 116444
rect 149916 116404 149956 116444
rect 149998 116404 150038 116444
rect 150080 116404 150120 116444
rect 75392 115648 75432 115688
rect 75474 115648 75514 115688
rect 75556 115648 75596 115688
rect 75638 115648 75678 115688
rect 75720 115648 75760 115688
rect 90512 115648 90552 115688
rect 90594 115648 90634 115688
rect 90676 115648 90716 115688
rect 90758 115648 90798 115688
rect 90840 115648 90880 115688
rect 105632 115648 105672 115688
rect 105714 115648 105754 115688
rect 105796 115648 105836 115688
rect 105878 115648 105918 115688
rect 105960 115648 106000 115688
rect 120752 115648 120792 115688
rect 120834 115648 120874 115688
rect 120916 115648 120956 115688
rect 120998 115648 121038 115688
rect 121080 115648 121120 115688
rect 135872 115648 135912 115688
rect 135954 115648 135994 115688
rect 136036 115648 136076 115688
rect 136118 115648 136158 115688
rect 136200 115648 136240 115688
rect 150992 115648 151032 115688
rect 151074 115648 151114 115688
rect 151156 115648 151196 115688
rect 151238 115648 151278 115688
rect 151320 115648 151360 115688
rect 74152 114892 74192 114932
rect 74234 114892 74274 114932
rect 74316 114892 74356 114932
rect 74398 114892 74438 114932
rect 74480 114892 74520 114932
rect 89272 114892 89312 114932
rect 89354 114892 89394 114932
rect 89436 114892 89476 114932
rect 89518 114892 89558 114932
rect 89600 114892 89640 114932
rect 104392 114892 104432 114932
rect 104474 114892 104514 114932
rect 104556 114892 104596 114932
rect 104638 114892 104678 114932
rect 104720 114892 104760 114932
rect 119512 114892 119552 114932
rect 119594 114892 119634 114932
rect 119676 114892 119716 114932
rect 119758 114892 119798 114932
rect 119840 114892 119880 114932
rect 134632 114892 134672 114932
rect 134714 114892 134754 114932
rect 134796 114892 134836 114932
rect 134878 114892 134918 114932
rect 134960 114892 135000 114932
rect 149752 114892 149792 114932
rect 149834 114892 149874 114932
rect 149916 114892 149956 114932
rect 149998 114892 150038 114932
rect 150080 114892 150120 114932
rect 75392 114136 75432 114176
rect 75474 114136 75514 114176
rect 75556 114136 75596 114176
rect 75638 114136 75678 114176
rect 75720 114136 75760 114176
rect 90512 114136 90552 114176
rect 90594 114136 90634 114176
rect 90676 114136 90716 114176
rect 90758 114136 90798 114176
rect 90840 114136 90880 114176
rect 105632 114136 105672 114176
rect 105714 114136 105754 114176
rect 105796 114136 105836 114176
rect 105878 114136 105918 114176
rect 105960 114136 106000 114176
rect 120752 114136 120792 114176
rect 120834 114136 120874 114176
rect 120916 114136 120956 114176
rect 120998 114136 121038 114176
rect 121080 114136 121120 114176
rect 135872 114136 135912 114176
rect 135954 114136 135994 114176
rect 136036 114136 136076 114176
rect 136118 114136 136158 114176
rect 136200 114136 136240 114176
rect 150992 114136 151032 114176
rect 151074 114136 151114 114176
rect 151156 114136 151196 114176
rect 151238 114136 151278 114176
rect 151320 114136 151360 114176
rect 74152 113380 74192 113420
rect 74234 113380 74274 113420
rect 74316 113380 74356 113420
rect 74398 113380 74438 113420
rect 74480 113380 74520 113420
rect 89272 113380 89312 113420
rect 89354 113380 89394 113420
rect 89436 113380 89476 113420
rect 89518 113380 89558 113420
rect 89600 113380 89640 113420
rect 104392 113380 104432 113420
rect 104474 113380 104514 113420
rect 104556 113380 104596 113420
rect 104638 113380 104678 113420
rect 104720 113380 104760 113420
rect 119512 113380 119552 113420
rect 119594 113380 119634 113420
rect 119676 113380 119716 113420
rect 119758 113380 119798 113420
rect 119840 113380 119880 113420
rect 134632 113380 134672 113420
rect 134714 113380 134754 113420
rect 134796 113380 134836 113420
rect 134878 113380 134918 113420
rect 134960 113380 135000 113420
rect 149752 113380 149792 113420
rect 149834 113380 149874 113420
rect 149916 113380 149956 113420
rect 149998 113380 150038 113420
rect 150080 113380 150120 113420
rect 75392 112624 75432 112664
rect 75474 112624 75514 112664
rect 75556 112624 75596 112664
rect 75638 112624 75678 112664
rect 75720 112624 75760 112664
rect 90512 112624 90552 112664
rect 90594 112624 90634 112664
rect 90676 112624 90716 112664
rect 90758 112624 90798 112664
rect 90840 112624 90880 112664
rect 105632 112624 105672 112664
rect 105714 112624 105754 112664
rect 105796 112624 105836 112664
rect 105878 112624 105918 112664
rect 105960 112624 106000 112664
rect 120752 112624 120792 112664
rect 120834 112624 120874 112664
rect 120916 112624 120956 112664
rect 120998 112624 121038 112664
rect 121080 112624 121120 112664
rect 135872 112624 135912 112664
rect 135954 112624 135994 112664
rect 136036 112624 136076 112664
rect 136118 112624 136158 112664
rect 136200 112624 136240 112664
rect 150992 112624 151032 112664
rect 151074 112624 151114 112664
rect 151156 112624 151196 112664
rect 151238 112624 151278 112664
rect 151320 112624 151360 112664
rect 74152 111868 74192 111908
rect 74234 111868 74274 111908
rect 74316 111868 74356 111908
rect 74398 111868 74438 111908
rect 74480 111868 74520 111908
rect 89272 111868 89312 111908
rect 89354 111868 89394 111908
rect 89436 111868 89476 111908
rect 89518 111868 89558 111908
rect 89600 111868 89640 111908
rect 104392 111868 104432 111908
rect 104474 111868 104514 111908
rect 104556 111868 104596 111908
rect 104638 111868 104678 111908
rect 104720 111868 104760 111908
rect 119512 111868 119552 111908
rect 119594 111868 119634 111908
rect 119676 111868 119716 111908
rect 119758 111868 119798 111908
rect 119840 111868 119880 111908
rect 134632 111868 134672 111908
rect 134714 111868 134754 111908
rect 134796 111868 134836 111908
rect 134878 111868 134918 111908
rect 134960 111868 135000 111908
rect 149752 111868 149792 111908
rect 149834 111868 149874 111908
rect 149916 111868 149956 111908
rect 149998 111868 150038 111908
rect 150080 111868 150120 111908
rect 75392 111112 75432 111152
rect 75474 111112 75514 111152
rect 75556 111112 75596 111152
rect 75638 111112 75678 111152
rect 75720 111112 75760 111152
rect 90512 111112 90552 111152
rect 90594 111112 90634 111152
rect 90676 111112 90716 111152
rect 90758 111112 90798 111152
rect 90840 111112 90880 111152
rect 105632 111112 105672 111152
rect 105714 111112 105754 111152
rect 105796 111112 105836 111152
rect 105878 111112 105918 111152
rect 105960 111112 106000 111152
rect 120752 111112 120792 111152
rect 120834 111112 120874 111152
rect 120916 111112 120956 111152
rect 120998 111112 121038 111152
rect 121080 111112 121120 111152
rect 135872 111112 135912 111152
rect 135954 111112 135994 111152
rect 136036 111112 136076 111152
rect 136118 111112 136158 111152
rect 136200 111112 136240 111152
rect 150992 111112 151032 111152
rect 151074 111112 151114 111152
rect 151156 111112 151196 111152
rect 151238 111112 151278 111152
rect 151320 111112 151360 111152
rect 74152 110356 74192 110396
rect 74234 110356 74274 110396
rect 74316 110356 74356 110396
rect 74398 110356 74438 110396
rect 74480 110356 74520 110396
rect 89272 110356 89312 110396
rect 89354 110356 89394 110396
rect 89436 110356 89476 110396
rect 89518 110356 89558 110396
rect 89600 110356 89640 110396
rect 104392 110356 104432 110396
rect 104474 110356 104514 110396
rect 104556 110356 104596 110396
rect 104638 110356 104678 110396
rect 104720 110356 104760 110396
rect 119512 110356 119552 110396
rect 119594 110356 119634 110396
rect 119676 110356 119716 110396
rect 119758 110356 119798 110396
rect 119840 110356 119880 110396
rect 134632 110356 134672 110396
rect 134714 110356 134754 110396
rect 134796 110356 134836 110396
rect 134878 110356 134918 110396
rect 134960 110356 135000 110396
rect 149752 110356 149792 110396
rect 149834 110356 149874 110396
rect 149916 110356 149956 110396
rect 149998 110356 150038 110396
rect 150080 110356 150120 110396
rect 75392 109600 75432 109640
rect 75474 109600 75514 109640
rect 75556 109600 75596 109640
rect 75638 109600 75678 109640
rect 75720 109600 75760 109640
rect 90512 109600 90552 109640
rect 90594 109600 90634 109640
rect 90676 109600 90716 109640
rect 90758 109600 90798 109640
rect 90840 109600 90880 109640
rect 105632 109600 105672 109640
rect 105714 109600 105754 109640
rect 105796 109600 105836 109640
rect 105878 109600 105918 109640
rect 105960 109600 106000 109640
rect 120752 109600 120792 109640
rect 120834 109600 120874 109640
rect 120916 109600 120956 109640
rect 120998 109600 121038 109640
rect 121080 109600 121120 109640
rect 135872 109600 135912 109640
rect 135954 109600 135994 109640
rect 136036 109600 136076 109640
rect 136118 109600 136158 109640
rect 136200 109600 136240 109640
rect 150992 109600 151032 109640
rect 151074 109600 151114 109640
rect 151156 109600 151196 109640
rect 151238 109600 151278 109640
rect 151320 109600 151360 109640
rect 74152 108844 74192 108884
rect 74234 108844 74274 108884
rect 74316 108844 74356 108884
rect 74398 108844 74438 108884
rect 74480 108844 74520 108884
rect 89272 108844 89312 108884
rect 89354 108844 89394 108884
rect 89436 108844 89476 108884
rect 89518 108844 89558 108884
rect 89600 108844 89640 108884
rect 104392 108844 104432 108884
rect 104474 108844 104514 108884
rect 104556 108844 104596 108884
rect 104638 108844 104678 108884
rect 104720 108844 104760 108884
rect 119512 108844 119552 108884
rect 119594 108844 119634 108884
rect 119676 108844 119716 108884
rect 119758 108844 119798 108884
rect 119840 108844 119880 108884
rect 134632 108844 134672 108884
rect 134714 108844 134754 108884
rect 134796 108844 134836 108884
rect 134878 108844 134918 108884
rect 134960 108844 135000 108884
rect 149752 108844 149792 108884
rect 149834 108844 149874 108884
rect 149916 108844 149956 108884
rect 149998 108844 150038 108884
rect 150080 108844 150120 108884
rect 75392 108088 75432 108128
rect 75474 108088 75514 108128
rect 75556 108088 75596 108128
rect 75638 108088 75678 108128
rect 75720 108088 75760 108128
rect 90512 108088 90552 108128
rect 90594 108088 90634 108128
rect 90676 108088 90716 108128
rect 90758 108088 90798 108128
rect 90840 108088 90880 108128
rect 105632 108088 105672 108128
rect 105714 108088 105754 108128
rect 105796 108088 105836 108128
rect 105878 108088 105918 108128
rect 105960 108088 106000 108128
rect 120752 108088 120792 108128
rect 120834 108088 120874 108128
rect 120916 108088 120956 108128
rect 120998 108088 121038 108128
rect 121080 108088 121120 108128
rect 135872 108088 135912 108128
rect 135954 108088 135994 108128
rect 136036 108088 136076 108128
rect 136118 108088 136158 108128
rect 136200 108088 136240 108128
rect 150992 108088 151032 108128
rect 151074 108088 151114 108128
rect 151156 108088 151196 108128
rect 151238 108088 151278 108128
rect 151320 108088 151360 108128
rect 74152 107332 74192 107372
rect 74234 107332 74274 107372
rect 74316 107332 74356 107372
rect 74398 107332 74438 107372
rect 74480 107332 74520 107372
rect 89272 107332 89312 107372
rect 89354 107332 89394 107372
rect 89436 107332 89476 107372
rect 89518 107332 89558 107372
rect 89600 107332 89640 107372
rect 104392 107332 104432 107372
rect 104474 107332 104514 107372
rect 104556 107332 104596 107372
rect 104638 107332 104678 107372
rect 104720 107332 104760 107372
rect 119512 107332 119552 107372
rect 119594 107332 119634 107372
rect 119676 107332 119716 107372
rect 119758 107332 119798 107372
rect 119840 107332 119880 107372
rect 134632 107332 134672 107372
rect 134714 107332 134754 107372
rect 134796 107332 134836 107372
rect 134878 107332 134918 107372
rect 134960 107332 135000 107372
rect 149752 107332 149792 107372
rect 149834 107332 149874 107372
rect 149916 107332 149956 107372
rect 149998 107332 150038 107372
rect 150080 107332 150120 107372
rect 75392 106576 75432 106616
rect 75474 106576 75514 106616
rect 75556 106576 75596 106616
rect 75638 106576 75678 106616
rect 75720 106576 75760 106616
rect 90512 106576 90552 106616
rect 90594 106576 90634 106616
rect 90676 106576 90716 106616
rect 90758 106576 90798 106616
rect 90840 106576 90880 106616
rect 105632 106576 105672 106616
rect 105714 106576 105754 106616
rect 105796 106576 105836 106616
rect 105878 106576 105918 106616
rect 105960 106576 106000 106616
rect 120752 106576 120792 106616
rect 120834 106576 120874 106616
rect 120916 106576 120956 106616
rect 120998 106576 121038 106616
rect 121080 106576 121120 106616
rect 135872 106576 135912 106616
rect 135954 106576 135994 106616
rect 136036 106576 136076 106616
rect 136118 106576 136158 106616
rect 136200 106576 136240 106616
rect 150992 106576 151032 106616
rect 151074 106576 151114 106616
rect 151156 106576 151196 106616
rect 151238 106576 151278 106616
rect 151320 106576 151360 106616
rect 74152 105820 74192 105860
rect 74234 105820 74274 105860
rect 74316 105820 74356 105860
rect 74398 105820 74438 105860
rect 74480 105820 74520 105860
rect 89272 105820 89312 105860
rect 89354 105820 89394 105860
rect 89436 105820 89476 105860
rect 89518 105820 89558 105860
rect 89600 105820 89640 105860
rect 104392 105820 104432 105860
rect 104474 105820 104514 105860
rect 104556 105820 104596 105860
rect 104638 105820 104678 105860
rect 104720 105820 104760 105860
rect 119512 105820 119552 105860
rect 119594 105820 119634 105860
rect 119676 105820 119716 105860
rect 119758 105820 119798 105860
rect 119840 105820 119880 105860
rect 134632 105820 134672 105860
rect 134714 105820 134754 105860
rect 134796 105820 134836 105860
rect 134878 105820 134918 105860
rect 134960 105820 135000 105860
rect 149752 105820 149792 105860
rect 149834 105820 149874 105860
rect 149916 105820 149956 105860
rect 149998 105820 150038 105860
rect 150080 105820 150120 105860
rect 75392 105064 75432 105104
rect 75474 105064 75514 105104
rect 75556 105064 75596 105104
rect 75638 105064 75678 105104
rect 75720 105064 75760 105104
rect 90512 105064 90552 105104
rect 90594 105064 90634 105104
rect 90676 105064 90716 105104
rect 90758 105064 90798 105104
rect 90840 105064 90880 105104
rect 105632 105064 105672 105104
rect 105714 105064 105754 105104
rect 105796 105064 105836 105104
rect 105878 105064 105918 105104
rect 105960 105064 106000 105104
rect 120752 105064 120792 105104
rect 120834 105064 120874 105104
rect 120916 105064 120956 105104
rect 120998 105064 121038 105104
rect 121080 105064 121120 105104
rect 135872 105064 135912 105104
rect 135954 105064 135994 105104
rect 136036 105064 136076 105104
rect 136118 105064 136158 105104
rect 136200 105064 136240 105104
rect 150992 105064 151032 105104
rect 151074 105064 151114 105104
rect 151156 105064 151196 105104
rect 151238 105064 151278 105104
rect 151320 105064 151360 105104
rect 74152 104308 74192 104348
rect 74234 104308 74274 104348
rect 74316 104308 74356 104348
rect 74398 104308 74438 104348
rect 74480 104308 74520 104348
rect 89272 104308 89312 104348
rect 89354 104308 89394 104348
rect 89436 104308 89476 104348
rect 89518 104308 89558 104348
rect 89600 104308 89640 104348
rect 104392 104308 104432 104348
rect 104474 104308 104514 104348
rect 104556 104308 104596 104348
rect 104638 104308 104678 104348
rect 104720 104308 104760 104348
rect 119512 104308 119552 104348
rect 119594 104308 119634 104348
rect 119676 104308 119716 104348
rect 119758 104308 119798 104348
rect 119840 104308 119880 104348
rect 134632 104308 134672 104348
rect 134714 104308 134754 104348
rect 134796 104308 134836 104348
rect 134878 104308 134918 104348
rect 134960 104308 135000 104348
rect 149752 104308 149792 104348
rect 149834 104308 149874 104348
rect 149916 104308 149956 104348
rect 149998 104308 150038 104348
rect 150080 104308 150120 104348
rect 75392 103552 75432 103592
rect 75474 103552 75514 103592
rect 75556 103552 75596 103592
rect 75638 103552 75678 103592
rect 75720 103552 75760 103592
rect 90512 103552 90552 103592
rect 90594 103552 90634 103592
rect 90676 103552 90716 103592
rect 90758 103552 90798 103592
rect 90840 103552 90880 103592
rect 105632 103552 105672 103592
rect 105714 103552 105754 103592
rect 105796 103552 105836 103592
rect 105878 103552 105918 103592
rect 105960 103552 106000 103592
rect 120752 103552 120792 103592
rect 120834 103552 120874 103592
rect 120916 103552 120956 103592
rect 120998 103552 121038 103592
rect 121080 103552 121120 103592
rect 135872 103552 135912 103592
rect 135954 103552 135994 103592
rect 136036 103552 136076 103592
rect 136118 103552 136158 103592
rect 136200 103552 136240 103592
rect 150992 103552 151032 103592
rect 151074 103552 151114 103592
rect 151156 103552 151196 103592
rect 151238 103552 151278 103592
rect 151320 103552 151360 103592
rect 74152 102796 74192 102836
rect 74234 102796 74274 102836
rect 74316 102796 74356 102836
rect 74398 102796 74438 102836
rect 74480 102796 74520 102836
rect 89272 102796 89312 102836
rect 89354 102796 89394 102836
rect 89436 102796 89476 102836
rect 89518 102796 89558 102836
rect 89600 102796 89640 102836
rect 104392 102796 104432 102836
rect 104474 102796 104514 102836
rect 104556 102796 104596 102836
rect 104638 102796 104678 102836
rect 104720 102796 104760 102836
rect 119512 102796 119552 102836
rect 119594 102796 119634 102836
rect 119676 102796 119716 102836
rect 119758 102796 119798 102836
rect 119840 102796 119880 102836
rect 134632 102796 134672 102836
rect 134714 102796 134754 102836
rect 134796 102796 134836 102836
rect 134878 102796 134918 102836
rect 134960 102796 135000 102836
rect 149752 102796 149792 102836
rect 149834 102796 149874 102836
rect 149916 102796 149956 102836
rect 149998 102796 150038 102836
rect 150080 102796 150120 102836
rect 75392 102040 75432 102080
rect 75474 102040 75514 102080
rect 75556 102040 75596 102080
rect 75638 102040 75678 102080
rect 75720 102040 75760 102080
rect 90512 102040 90552 102080
rect 90594 102040 90634 102080
rect 90676 102040 90716 102080
rect 90758 102040 90798 102080
rect 90840 102040 90880 102080
rect 105632 102040 105672 102080
rect 105714 102040 105754 102080
rect 105796 102040 105836 102080
rect 105878 102040 105918 102080
rect 105960 102040 106000 102080
rect 120752 102040 120792 102080
rect 120834 102040 120874 102080
rect 120916 102040 120956 102080
rect 120998 102040 121038 102080
rect 121080 102040 121120 102080
rect 135872 102040 135912 102080
rect 135954 102040 135994 102080
rect 136036 102040 136076 102080
rect 136118 102040 136158 102080
rect 136200 102040 136240 102080
rect 150992 102040 151032 102080
rect 151074 102040 151114 102080
rect 151156 102040 151196 102080
rect 151238 102040 151278 102080
rect 151320 102040 151360 102080
rect 74152 101284 74192 101324
rect 74234 101284 74274 101324
rect 74316 101284 74356 101324
rect 74398 101284 74438 101324
rect 74480 101284 74520 101324
rect 89272 101284 89312 101324
rect 89354 101284 89394 101324
rect 89436 101284 89476 101324
rect 89518 101284 89558 101324
rect 89600 101284 89640 101324
rect 104392 101284 104432 101324
rect 104474 101284 104514 101324
rect 104556 101284 104596 101324
rect 104638 101284 104678 101324
rect 104720 101284 104760 101324
rect 119512 101284 119552 101324
rect 119594 101284 119634 101324
rect 119676 101284 119716 101324
rect 119758 101284 119798 101324
rect 119840 101284 119880 101324
rect 134632 101284 134672 101324
rect 134714 101284 134754 101324
rect 134796 101284 134836 101324
rect 134878 101284 134918 101324
rect 134960 101284 135000 101324
rect 149752 101284 149792 101324
rect 149834 101284 149874 101324
rect 149916 101284 149956 101324
rect 149998 101284 150038 101324
rect 150080 101284 150120 101324
rect 75392 100528 75432 100568
rect 75474 100528 75514 100568
rect 75556 100528 75596 100568
rect 75638 100528 75678 100568
rect 75720 100528 75760 100568
rect 90512 100528 90552 100568
rect 90594 100528 90634 100568
rect 90676 100528 90716 100568
rect 90758 100528 90798 100568
rect 90840 100528 90880 100568
rect 105632 100528 105672 100568
rect 105714 100528 105754 100568
rect 105796 100528 105836 100568
rect 105878 100528 105918 100568
rect 105960 100528 106000 100568
rect 120752 100528 120792 100568
rect 120834 100528 120874 100568
rect 120916 100528 120956 100568
rect 120998 100528 121038 100568
rect 121080 100528 121120 100568
rect 135872 100528 135912 100568
rect 135954 100528 135994 100568
rect 136036 100528 136076 100568
rect 136118 100528 136158 100568
rect 136200 100528 136240 100568
rect 150992 100528 151032 100568
rect 151074 100528 151114 100568
rect 151156 100528 151196 100568
rect 151238 100528 151278 100568
rect 151320 100528 151360 100568
rect 74152 99772 74192 99812
rect 74234 99772 74274 99812
rect 74316 99772 74356 99812
rect 74398 99772 74438 99812
rect 74480 99772 74520 99812
rect 89272 99772 89312 99812
rect 89354 99772 89394 99812
rect 89436 99772 89476 99812
rect 89518 99772 89558 99812
rect 89600 99772 89640 99812
rect 104392 99772 104432 99812
rect 104474 99772 104514 99812
rect 104556 99772 104596 99812
rect 104638 99772 104678 99812
rect 104720 99772 104760 99812
rect 119512 99772 119552 99812
rect 119594 99772 119634 99812
rect 119676 99772 119716 99812
rect 119758 99772 119798 99812
rect 119840 99772 119880 99812
rect 134632 99772 134672 99812
rect 134714 99772 134754 99812
rect 134796 99772 134836 99812
rect 134878 99772 134918 99812
rect 134960 99772 135000 99812
rect 149752 99772 149792 99812
rect 149834 99772 149874 99812
rect 149916 99772 149956 99812
rect 149998 99772 150038 99812
rect 150080 99772 150120 99812
rect 75392 99016 75432 99056
rect 75474 99016 75514 99056
rect 75556 99016 75596 99056
rect 75638 99016 75678 99056
rect 75720 99016 75760 99056
rect 90512 99016 90552 99056
rect 90594 99016 90634 99056
rect 90676 99016 90716 99056
rect 90758 99016 90798 99056
rect 90840 99016 90880 99056
rect 105632 99016 105672 99056
rect 105714 99016 105754 99056
rect 105796 99016 105836 99056
rect 105878 99016 105918 99056
rect 105960 99016 106000 99056
rect 120752 99016 120792 99056
rect 120834 99016 120874 99056
rect 120916 99016 120956 99056
rect 120998 99016 121038 99056
rect 121080 99016 121120 99056
rect 135872 99016 135912 99056
rect 135954 99016 135994 99056
rect 136036 99016 136076 99056
rect 136118 99016 136158 99056
rect 136200 99016 136240 99056
rect 150992 99016 151032 99056
rect 151074 99016 151114 99056
rect 151156 99016 151196 99056
rect 151238 99016 151278 99056
rect 151320 99016 151360 99056
rect 74152 98260 74192 98300
rect 74234 98260 74274 98300
rect 74316 98260 74356 98300
rect 74398 98260 74438 98300
rect 74480 98260 74520 98300
rect 89272 98260 89312 98300
rect 89354 98260 89394 98300
rect 89436 98260 89476 98300
rect 89518 98260 89558 98300
rect 89600 98260 89640 98300
rect 104392 98260 104432 98300
rect 104474 98260 104514 98300
rect 104556 98260 104596 98300
rect 104638 98260 104678 98300
rect 104720 98260 104760 98300
rect 119512 98260 119552 98300
rect 119594 98260 119634 98300
rect 119676 98260 119716 98300
rect 119758 98260 119798 98300
rect 119840 98260 119880 98300
rect 134632 98260 134672 98300
rect 134714 98260 134754 98300
rect 134796 98260 134836 98300
rect 134878 98260 134918 98300
rect 134960 98260 135000 98300
rect 149752 98260 149792 98300
rect 149834 98260 149874 98300
rect 149916 98260 149956 98300
rect 149998 98260 150038 98300
rect 150080 98260 150120 98300
rect 75392 97504 75432 97544
rect 75474 97504 75514 97544
rect 75556 97504 75596 97544
rect 75638 97504 75678 97544
rect 75720 97504 75760 97544
rect 90512 97504 90552 97544
rect 90594 97504 90634 97544
rect 90676 97504 90716 97544
rect 90758 97504 90798 97544
rect 90840 97504 90880 97544
rect 105632 97504 105672 97544
rect 105714 97504 105754 97544
rect 105796 97504 105836 97544
rect 105878 97504 105918 97544
rect 105960 97504 106000 97544
rect 120752 97504 120792 97544
rect 120834 97504 120874 97544
rect 120916 97504 120956 97544
rect 120998 97504 121038 97544
rect 121080 97504 121120 97544
rect 135872 97504 135912 97544
rect 135954 97504 135994 97544
rect 136036 97504 136076 97544
rect 136118 97504 136158 97544
rect 136200 97504 136240 97544
rect 150992 97504 151032 97544
rect 151074 97504 151114 97544
rect 151156 97504 151196 97544
rect 151238 97504 151278 97544
rect 151320 97504 151360 97544
rect 74152 96748 74192 96788
rect 74234 96748 74274 96788
rect 74316 96748 74356 96788
rect 74398 96748 74438 96788
rect 74480 96748 74520 96788
rect 89272 96748 89312 96788
rect 89354 96748 89394 96788
rect 89436 96748 89476 96788
rect 89518 96748 89558 96788
rect 89600 96748 89640 96788
rect 104392 96748 104432 96788
rect 104474 96748 104514 96788
rect 104556 96748 104596 96788
rect 104638 96748 104678 96788
rect 104720 96748 104760 96788
rect 119512 96748 119552 96788
rect 119594 96748 119634 96788
rect 119676 96748 119716 96788
rect 119758 96748 119798 96788
rect 119840 96748 119880 96788
rect 134632 96748 134672 96788
rect 134714 96748 134754 96788
rect 134796 96748 134836 96788
rect 134878 96748 134918 96788
rect 134960 96748 135000 96788
rect 149752 96748 149792 96788
rect 149834 96748 149874 96788
rect 149916 96748 149956 96788
rect 149998 96748 150038 96788
rect 150080 96748 150120 96788
rect 75392 95992 75432 96032
rect 75474 95992 75514 96032
rect 75556 95992 75596 96032
rect 75638 95992 75678 96032
rect 75720 95992 75760 96032
rect 90512 95992 90552 96032
rect 90594 95992 90634 96032
rect 90676 95992 90716 96032
rect 90758 95992 90798 96032
rect 90840 95992 90880 96032
rect 105632 95992 105672 96032
rect 105714 95992 105754 96032
rect 105796 95992 105836 96032
rect 105878 95992 105918 96032
rect 105960 95992 106000 96032
rect 120752 95992 120792 96032
rect 120834 95992 120874 96032
rect 120916 95992 120956 96032
rect 120998 95992 121038 96032
rect 121080 95992 121120 96032
rect 135872 95992 135912 96032
rect 135954 95992 135994 96032
rect 136036 95992 136076 96032
rect 136118 95992 136158 96032
rect 136200 95992 136240 96032
rect 150992 95992 151032 96032
rect 151074 95992 151114 96032
rect 151156 95992 151196 96032
rect 151238 95992 151278 96032
rect 151320 95992 151360 96032
rect 74152 95236 74192 95276
rect 74234 95236 74274 95276
rect 74316 95236 74356 95276
rect 74398 95236 74438 95276
rect 74480 95236 74520 95276
rect 89272 95236 89312 95276
rect 89354 95236 89394 95276
rect 89436 95236 89476 95276
rect 89518 95236 89558 95276
rect 89600 95236 89640 95276
rect 104392 95236 104432 95276
rect 104474 95236 104514 95276
rect 104556 95236 104596 95276
rect 104638 95236 104678 95276
rect 104720 95236 104760 95276
rect 119512 95236 119552 95276
rect 119594 95236 119634 95276
rect 119676 95236 119716 95276
rect 119758 95236 119798 95276
rect 119840 95236 119880 95276
rect 134632 95236 134672 95276
rect 134714 95236 134754 95276
rect 134796 95236 134836 95276
rect 134878 95236 134918 95276
rect 134960 95236 135000 95276
rect 149752 95236 149792 95276
rect 149834 95236 149874 95276
rect 149916 95236 149956 95276
rect 149998 95236 150038 95276
rect 150080 95236 150120 95276
rect 75392 94480 75432 94520
rect 75474 94480 75514 94520
rect 75556 94480 75596 94520
rect 75638 94480 75678 94520
rect 75720 94480 75760 94520
rect 90512 94480 90552 94520
rect 90594 94480 90634 94520
rect 90676 94480 90716 94520
rect 90758 94480 90798 94520
rect 90840 94480 90880 94520
rect 105632 94480 105672 94520
rect 105714 94480 105754 94520
rect 105796 94480 105836 94520
rect 105878 94480 105918 94520
rect 105960 94480 106000 94520
rect 120752 94480 120792 94520
rect 120834 94480 120874 94520
rect 120916 94480 120956 94520
rect 120998 94480 121038 94520
rect 121080 94480 121120 94520
rect 135872 94480 135912 94520
rect 135954 94480 135994 94520
rect 136036 94480 136076 94520
rect 136118 94480 136158 94520
rect 136200 94480 136240 94520
rect 150992 94480 151032 94520
rect 151074 94480 151114 94520
rect 151156 94480 151196 94520
rect 151238 94480 151278 94520
rect 151320 94480 151360 94520
rect 74152 93724 74192 93764
rect 74234 93724 74274 93764
rect 74316 93724 74356 93764
rect 74398 93724 74438 93764
rect 74480 93724 74520 93764
rect 89272 93724 89312 93764
rect 89354 93724 89394 93764
rect 89436 93724 89476 93764
rect 89518 93724 89558 93764
rect 89600 93724 89640 93764
rect 104392 93724 104432 93764
rect 104474 93724 104514 93764
rect 104556 93724 104596 93764
rect 104638 93724 104678 93764
rect 104720 93724 104760 93764
rect 119512 93724 119552 93764
rect 119594 93724 119634 93764
rect 119676 93724 119716 93764
rect 119758 93724 119798 93764
rect 119840 93724 119880 93764
rect 134632 93724 134672 93764
rect 134714 93724 134754 93764
rect 134796 93724 134836 93764
rect 134878 93724 134918 93764
rect 134960 93724 135000 93764
rect 149752 93724 149792 93764
rect 149834 93724 149874 93764
rect 149916 93724 149956 93764
rect 149998 93724 150038 93764
rect 150080 93724 150120 93764
rect 75392 92968 75432 93008
rect 75474 92968 75514 93008
rect 75556 92968 75596 93008
rect 75638 92968 75678 93008
rect 75720 92968 75760 93008
rect 90512 92968 90552 93008
rect 90594 92968 90634 93008
rect 90676 92968 90716 93008
rect 90758 92968 90798 93008
rect 90840 92968 90880 93008
rect 105632 92968 105672 93008
rect 105714 92968 105754 93008
rect 105796 92968 105836 93008
rect 105878 92968 105918 93008
rect 105960 92968 106000 93008
rect 120752 92968 120792 93008
rect 120834 92968 120874 93008
rect 120916 92968 120956 93008
rect 120998 92968 121038 93008
rect 121080 92968 121120 93008
rect 135872 92968 135912 93008
rect 135954 92968 135994 93008
rect 136036 92968 136076 93008
rect 136118 92968 136158 93008
rect 136200 92968 136240 93008
rect 150992 92968 151032 93008
rect 151074 92968 151114 93008
rect 151156 92968 151196 93008
rect 151238 92968 151278 93008
rect 151320 92968 151360 93008
rect 74152 92212 74192 92252
rect 74234 92212 74274 92252
rect 74316 92212 74356 92252
rect 74398 92212 74438 92252
rect 74480 92212 74520 92252
rect 89272 92212 89312 92252
rect 89354 92212 89394 92252
rect 89436 92212 89476 92252
rect 89518 92212 89558 92252
rect 89600 92212 89640 92252
rect 104392 92212 104432 92252
rect 104474 92212 104514 92252
rect 104556 92212 104596 92252
rect 104638 92212 104678 92252
rect 104720 92212 104760 92252
rect 119512 92212 119552 92252
rect 119594 92212 119634 92252
rect 119676 92212 119716 92252
rect 119758 92212 119798 92252
rect 119840 92212 119880 92252
rect 134632 92212 134672 92252
rect 134714 92212 134754 92252
rect 134796 92212 134836 92252
rect 134878 92212 134918 92252
rect 134960 92212 135000 92252
rect 149752 92212 149792 92252
rect 149834 92212 149874 92252
rect 149916 92212 149956 92252
rect 149998 92212 150038 92252
rect 150080 92212 150120 92252
rect 75392 91456 75432 91496
rect 75474 91456 75514 91496
rect 75556 91456 75596 91496
rect 75638 91456 75678 91496
rect 75720 91456 75760 91496
rect 90512 91456 90552 91496
rect 90594 91456 90634 91496
rect 90676 91456 90716 91496
rect 90758 91456 90798 91496
rect 90840 91456 90880 91496
rect 105632 91456 105672 91496
rect 105714 91456 105754 91496
rect 105796 91456 105836 91496
rect 105878 91456 105918 91496
rect 105960 91456 106000 91496
rect 120752 91456 120792 91496
rect 120834 91456 120874 91496
rect 120916 91456 120956 91496
rect 120998 91456 121038 91496
rect 121080 91456 121120 91496
rect 135872 91456 135912 91496
rect 135954 91456 135994 91496
rect 136036 91456 136076 91496
rect 136118 91456 136158 91496
rect 136200 91456 136240 91496
rect 150992 91456 151032 91496
rect 151074 91456 151114 91496
rect 151156 91456 151196 91496
rect 151238 91456 151278 91496
rect 151320 91456 151360 91496
rect 74152 90700 74192 90740
rect 74234 90700 74274 90740
rect 74316 90700 74356 90740
rect 74398 90700 74438 90740
rect 74480 90700 74520 90740
rect 89272 90700 89312 90740
rect 89354 90700 89394 90740
rect 89436 90700 89476 90740
rect 89518 90700 89558 90740
rect 89600 90700 89640 90740
rect 104392 90700 104432 90740
rect 104474 90700 104514 90740
rect 104556 90700 104596 90740
rect 104638 90700 104678 90740
rect 104720 90700 104760 90740
rect 119512 90700 119552 90740
rect 119594 90700 119634 90740
rect 119676 90700 119716 90740
rect 119758 90700 119798 90740
rect 119840 90700 119880 90740
rect 134632 90700 134672 90740
rect 134714 90700 134754 90740
rect 134796 90700 134836 90740
rect 134878 90700 134918 90740
rect 134960 90700 135000 90740
rect 149752 90700 149792 90740
rect 149834 90700 149874 90740
rect 149916 90700 149956 90740
rect 149998 90700 150038 90740
rect 150080 90700 150120 90740
rect 75392 89944 75432 89984
rect 75474 89944 75514 89984
rect 75556 89944 75596 89984
rect 75638 89944 75678 89984
rect 75720 89944 75760 89984
rect 90512 89944 90552 89984
rect 90594 89944 90634 89984
rect 90676 89944 90716 89984
rect 90758 89944 90798 89984
rect 90840 89944 90880 89984
rect 105632 89944 105672 89984
rect 105714 89944 105754 89984
rect 105796 89944 105836 89984
rect 105878 89944 105918 89984
rect 105960 89944 106000 89984
rect 120752 89944 120792 89984
rect 120834 89944 120874 89984
rect 120916 89944 120956 89984
rect 120998 89944 121038 89984
rect 121080 89944 121120 89984
rect 135872 89944 135912 89984
rect 135954 89944 135994 89984
rect 136036 89944 136076 89984
rect 136118 89944 136158 89984
rect 136200 89944 136240 89984
rect 150992 89944 151032 89984
rect 151074 89944 151114 89984
rect 151156 89944 151196 89984
rect 151238 89944 151278 89984
rect 151320 89944 151360 89984
rect 74152 89188 74192 89228
rect 74234 89188 74274 89228
rect 74316 89188 74356 89228
rect 74398 89188 74438 89228
rect 74480 89188 74520 89228
rect 89272 89188 89312 89228
rect 89354 89188 89394 89228
rect 89436 89188 89476 89228
rect 89518 89188 89558 89228
rect 89600 89188 89640 89228
rect 104392 89188 104432 89228
rect 104474 89188 104514 89228
rect 104556 89188 104596 89228
rect 104638 89188 104678 89228
rect 104720 89188 104760 89228
rect 119512 89188 119552 89228
rect 119594 89188 119634 89228
rect 119676 89188 119716 89228
rect 119758 89188 119798 89228
rect 119840 89188 119880 89228
rect 134632 89188 134672 89228
rect 134714 89188 134754 89228
rect 134796 89188 134836 89228
rect 134878 89188 134918 89228
rect 134960 89188 135000 89228
rect 149752 89188 149792 89228
rect 149834 89188 149874 89228
rect 149916 89188 149956 89228
rect 149998 89188 150038 89228
rect 150080 89188 150120 89228
rect 75392 88432 75432 88472
rect 75474 88432 75514 88472
rect 75556 88432 75596 88472
rect 75638 88432 75678 88472
rect 75720 88432 75760 88472
rect 90512 88432 90552 88472
rect 90594 88432 90634 88472
rect 90676 88432 90716 88472
rect 90758 88432 90798 88472
rect 90840 88432 90880 88472
rect 105632 88432 105672 88472
rect 105714 88432 105754 88472
rect 105796 88432 105836 88472
rect 105878 88432 105918 88472
rect 105960 88432 106000 88472
rect 120752 88432 120792 88472
rect 120834 88432 120874 88472
rect 120916 88432 120956 88472
rect 120998 88432 121038 88472
rect 121080 88432 121120 88472
rect 135872 88432 135912 88472
rect 135954 88432 135994 88472
rect 136036 88432 136076 88472
rect 136118 88432 136158 88472
rect 136200 88432 136240 88472
rect 150992 88432 151032 88472
rect 151074 88432 151114 88472
rect 151156 88432 151196 88472
rect 151238 88432 151278 88472
rect 151320 88432 151360 88472
rect 74152 87676 74192 87716
rect 74234 87676 74274 87716
rect 74316 87676 74356 87716
rect 74398 87676 74438 87716
rect 74480 87676 74520 87716
rect 89272 87676 89312 87716
rect 89354 87676 89394 87716
rect 89436 87676 89476 87716
rect 89518 87676 89558 87716
rect 89600 87676 89640 87716
rect 104392 87676 104432 87716
rect 104474 87676 104514 87716
rect 104556 87676 104596 87716
rect 104638 87676 104678 87716
rect 104720 87676 104760 87716
rect 119512 87676 119552 87716
rect 119594 87676 119634 87716
rect 119676 87676 119716 87716
rect 119758 87676 119798 87716
rect 119840 87676 119880 87716
rect 134632 87676 134672 87716
rect 134714 87676 134754 87716
rect 134796 87676 134836 87716
rect 134878 87676 134918 87716
rect 134960 87676 135000 87716
rect 149752 87676 149792 87716
rect 149834 87676 149874 87716
rect 149916 87676 149956 87716
rect 149998 87676 150038 87716
rect 150080 87676 150120 87716
rect 75392 86920 75432 86960
rect 75474 86920 75514 86960
rect 75556 86920 75596 86960
rect 75638 86920 75678 86960
rect 75720 86920 75760 86960
rect 90512 86920 90552 86960
rect 90594 86920 90634 86960
rect 90676 86920 90716 86960
rect 90758 86920 90798 86960
rect 90840 86920 90880 86960
rect 105632 86920 105672 86960
rect 105714 86920 105754 86960
rect 105796 86920 105836 86960
rect 105878 86920 105918 86960
rect 105960 86920 106000 86960
rect 120752 86920 120792 86960
rect 120834 86920 120874 86960
rect 120916 86920 120956 86960
rect 120998 86920 121038 86960
rect 121080 86920 121120 86960
rect 135872 86920 135912 86960
rect 135954 86920 135994 86960
rect 136036 86920 136076 86960
rect 136118 86920 136158 86960
rect 136200 86920 136240 86960
rect 150992 86920 151032 86960
rect 151074 86920 151114 86960
rect 151156 86920 151196 86960
rect 151238 86920 151278 86960
rect 151320 86920 151360 86960
rect 74152 86164 74192 86204
rect 74234 86164 74274 86204
rect 74316 86164 74356 86204
rect 74398 86164 74438 86204
rect 74480 86164 74520 86204
rect 89272 86164 89312 86204
rect 89354 86164 89394 86204
rect 89436 86164 89476 86204
rect 89518 86164 89558 86204
rect 89600 86164 89640 86204
rect 104392 86164 104432 86204
rect 104474 86164 104514 86204
rect 104556 86164 104596 86204
rect 104638 86164 104678 86204
rect 104720 86164 104760 86204
rect 119512 86164 119552 86204
rect 119594 86164 119634 86204
rect 119676 86164 119716 86204
rect 119758 86164 119798 86204
rect 119840 86164 119880 86204
rect 134632 86164 134672 86204
rect 134714 86164 134754 86204
rect 134796 86164 134836 86204
rect 134878 86164 134918 86204
rect 134960 86164 135000 86204
rect 149752 86164 149792 86204
rect 149834 86164 149874 86204
rect 149916 86164 149956 86204
rect 149998 86164 150038 86204
rect 150080 86164 150120 86204
rect 75392 85408 75432 85448
rect 75474 85408 75514 85448
rect 75556 85408 75596 85448
rect 75638 85408 75678 85448
rect 75720 85408 75760 85448
rect 90512 85408 90552 85448
rect 90594 85408 90634 85448
rect 90676 85408 90716 85448
rect 90758 85408 90798 85448
rect 90840 85408 90880 85448
rect 105632 85408 105672 85448
rect 105714 85408 105754 85448
rect 105796 85408 105836 85448
rect 105878 85408 105918 85448
rect 105960 85408 106000 85448
rect 120752 85408 120792 85448
rect 120834 85408 120874 85448
rect 120916 85408 120956 85448
rect 120998 85408 121038 85448
rect 121080 85408 121120 85448
rect 135872 85408 135912 85448
rect 135954 85408 135994 85448
rect 136036 85408 136076 85448
rect 136118 85408 136158 85448
rect 136200 85408 136240 85448
rect 150992 85408 151032 85448
rect 151074 85408 151114 85448
rect 151156 85408 151196 85448
rect 151238 85408 151278 85448
rect 151320 85408 151360 85448
rect 74152 84652 74192 84692
rect 74234 84652 74274 84692
rect 74316 84652 74356 84692
rect 74398 84652 74438 84692
rect 74480 84652 74520 84692
rect 89272 84652 89312 84692
rect 89354 84652 89394 84692
rect 89436 84652 89476 84692
rect 89518 84652 89558 84692
rect 89600 84652 89640 84692
rect 104392 84652 104432 84692
rect 104474 84652 104514 84692
rect 104556 84652 104596 84692
rect 104638 84652 104678 84692
rect 104720 84652 104760 84692
rect 119512 84652 119552 84692
rect 119594 84652 119634 84692
rect 119676 84652 119716 84692
rect 119758 84652 119798 84692
rect 119840 84652 119880 84692
rect 134632 84652 134672 84692
rect 134714 84652 134754 84692
rect 134796 84652 134836 84692
rect 134878 84652 134918 84692
rect 134960 84652 135000 84692
rect 149752 84652 149792 84692
rect 149834 84652 149874 84692
rect 149916 84652 149956 84692
rect 149998 84652 150038 84692
rect 150080 84652 150120 84692
rect 75392 83896 75432 83936
rect 75474 83896 75514 83936
rect 75556 83896 75596 83936
rect 75638 83896 75678 83936
rect 75720 83896 75760 83936
rect 90512 83896 90552 83936
rect 90594 83896 90634 83936
rect 90676 83896 90716 83936
rect 90758 83896 90798 83936
rect 90840 83896 90880 83936
rect 105632 83896 105672 83936
rect 105714 83896 105754 83936
rect 105796 83896 105836 83936
rect 105878 83896 105918 83936
rect 105960 83896 106000 83936
rect 120752 83896 120792 83936
rect 120834 83896 120874 83936
rect 120916 83896 120956 83936
rect 120998 83896 121038 83936
rect 121080 83896 121120 83936
rect 135872 83896 135912 83936
rect 135954 83896 135994 83936
rect 136036 83896 136076 83936
rect 136118 83896 136158 83936
rect 136200 83896 136240 83936
rect 150992 83896 151032 83936
rect 151074 83896 151114 83936
rect 151156 83896 151196 83936
rect 151238 83896 151278 83936
rect 151320 83896 151360 83936
rect 74152 83140 74192 83180
rect 74234 83140 74274 83180
rect 74316 83140 74356 83180
rect 74398 83140 74438 83180
rect 74480 83140 74520 83180
rect 89272 83140 89312 83180
rect 89354 83140 89394 83180
rect 89436 83140 89476 83180
rect 89518 83140 89558 83180
rect 89600 83140 89640 83180
rect 104392 83140 104432 83180
rect 104474 83140 104514 83180
rect 104556 83140 104596 83180
rect 104638 83140 104678 83180
rect 104720 83140 104760 83180
rect 119512 83140 119552 83180
rect 119594 83140 119634 83180
rect 119676 83140 119716 83180
rect 119758 83140 119798 83180
rect 119840 83140 119880 83180
rect 134632 83140 134672 83180
rect 134714 83140 134754 83180
rect 134796 83140 134836 83180
rect 134878 83140 134918 83180
rect 134960 83140 135000 83180
rect 149752 83140 149792 83180
rect 149834 83140 149874 83180
rect 149916 83140 149956 83180
rect 149998 83140 150038 83180
rect 150080 83140 150120 83180
rect 75392 82384 75432 82424
rect 75474 82384 75514 82424
rect 75556 82384 75596 82424
rect 75638 82384 75678 82424
rect 75720 82384 75760 82424
rect 90512 82384 90552 82424
rect 90594 82384 90634 82424
rect 90676 82384 90716 82424
rect 90758 82384 90798 82424
rect 90840 82384 90880 82424
rect 105632 82384 105672 82424
rect 105714 82384 105754 82424
rect 105796 82384 105836 82424
rect 105878 82384 105918 82424
rect 105960 82384 106000 82424
rect 120752 82384 120792 82424
rect 120834 82384 120874 82424
rect 120916 82384 120956 82424
rect 120998 82384 121038 82424
rect 121080 82384 121120 82424
rect 135872 82384 135912 82424
rect 135954 82384 135994 82424
rect 136036 82384 136076 82424
rect 136118 82384 136158 82424
rect 136200 82384 136240 82424
rect 150992 82384 151032 82424
rect 151074 82384 151114 82424
rect 151156 82384 151196 82424
rect 151238 82384 151278 82424
rect 151320 82384 151360 82424
rect 74152 81628 74192 81668
rect 74234 81628 74274 81668
rect 74316 81628 74356 81668
rect 74398 81628 74438 81668
rect 74480 81628 74520 81668
rect 89272 81628 89312 81668
rect 89354 81628 89394 81668
rect 89436 81628 89476 81668
rect 89518 81628 89558 81668
rect 89600 81628 89640 81668
rect 104392 81628 104432 81668
rect 104474 81628 104514 81668
rect 104556 81628 104596 81668
rect 104638 81628 104678 81668
rect 104720 81628 104760 81668
rect 119512 81628 119552 81668
rect 119594 81628 119634 81668
rect 119676 81628 119716 81668
rect 119758 81628 119798 81668
rect 119840 81628 119880 81668
rect 134632 81628 134672 81668
rect 134714 81628 134754 81668
rect 134796 81628 134836 81668
rect 134878 81628 134918 81668
rect 134960 81628 135000 81668
rect 149752 81628 149792 81668
rect 149834 81628 149874 81668
rect 149916 81628 149956 81668
rect 149998 81628 150038 81668
rect 150080 81628 150120 81668
rect 75392 80872 75432 80912
rect 75474 80872 75514 80912
rect 75556 80872 75596 80912
rect 75638 80872 75678 80912
rect 75720 80872 75760 80912
rect 90512 80872 90552 80912
rect 90594 80872 90634 80912
rect 90676 80872 90716 80912
rect 90758 80872 90798 80912
rect 90840 80872 90880 80912
rect 105632 80872 105672 80912
rect 105714 80872 105754 80912
rect 105796 80872 105836 80912
rect 105878 80872 105918 80912
rect 105960 80872 106000 80912
rect 120752 80872 120792 80912
rect 120834 80872 120874 80912
rect 120916 80872 120956 80912
rect 120998 80872 121038 80912
rect 121080 80872 121120 80912
rect 135872 80872 135912 80912
rect 135954 80872 135994 80912
rect 136036 80872 136076 80912
rect 136118 80872 136158 80912
rect 136200 80872 136240 80912
rect 150992 80872 151032 80912
rect 151074 80872 151114 80912
rect 151156 80872 151196 80912
rect 151238 80872 151278 80912
rect 151320 80872 151360 80912
rect 74152 80116 74192 80156
rect 74234 80116 74274 80156
rect 74316 80116 74356 80156
rect 74398 80116 74438 80156
rect 74480 80116 74520 80156
rect 89272 80116 89312 80156
rect 89354 80116 89394 80156
rect 89436 80116 89476 80156
rect 89518 80116 89558 80156
rect 89600 80116 89640 80156
rect 104392 80116 104432 80156
rect 104474 80116 104514 80156
rect 104556 80116 104596 80156
rect 104638 80116 104678 80156
rect 104720 80116 104760 80156
rect 119512 80116 119552 80156
rect 119594 80116 119634 80156
rect 119676 80116 119716 80156
rect 119758 80116 119798 80156
rect 119840 80116 119880 80156
rect 134632 80116 134672 80156
rect 134714 80116 134754 80156
rect 134796 80116 134836 80156
rect 134878 80116 134918 80156
rect 134960 80116 135000 80156
rect 149752 80116 149792 80156
rect 149834 80116 149874 80156
rect 149916 80116 149956 80156
rect 149998 80116 150038 80156
rect 150080 80116 150120 80156
rect 75392 79360 75432 79400
rect 75474 79360 75514 79400
rect 75556 79360 75596 79400
rect 75638 79360 75678 79400
rect 75720 79360 75760 79400
rect 90512 79360 90552 79400
rect 90594 79360 90634 79400
rect 90676 79360 90716 79400
rect 90758 79360 90798 79400
rect 90840 79360 90880 79400
rect 105632 79360 105672 79400
rect 105714 79360 105754 79400
rect 105796 79360 105836 79400
rect 105878 79360 105918 79400
rect 105960 79360 106000 79400
rect 120752 79360 120792 79400
rect 120834 79360 120874 79400
rect 120916 79360 120956 79400
rect 120998 79360 121038 79400
rect 121080 79360 121120 79400
rect 135872 79360 135912 79400
rect 135954 79360 135994 79400
rect 136036 79360 136076 79400
rect 136118 79360 136158 79400
rect 136200 79360 136240 79400
rect 150992 79360 151032 79400
rect 151074 79360 151114 79400
rect 151156 79360 151196 79400
rect 151238 79360 151278 79400
rect 151320 79360 151360 79400
rect 74152 78604 74192 78644
rect 74234 78604 74274 78644
rect 74316 78604 74356 78644
rect 74398 78604 74438 78644
rect 74480 78604 74520 78644
rect 89272 78604 89312 78644
rect 89354 78604 89394 78644
rect 89436 78604 89476 78644
rect 89518 78604 89558 78644
rect 89600 78604 89640 78644
rect 104392 78604 104432 78644
rect 104474 78604 104514 78644
rect 104556 78604 104596 78644
rect 104638 78604 104678 78644
rect 104720 78604 104760 78644
rect 119512 78604 119552 78644
rect 119594 78604 119634 78644
rect 119676 78604 119716 78644
rect 119758 78604 119798 78644
rect 119840 78604 119880 78644
rect 134632 78604 134672 78644
rect 134714 78604 134754 78644
rect 134796 78604 134836 78644
rect 134878 78604 134918 78644
rect 134960 78604 135000 78644
rect 149752 78604 149792 78644
rect 149834 78604 149874 78644
rect 149916 78604 149956 78644
rect 149998 78604 150038 78644
rect 150080 78604 150120 78644
rect 75392 77848 75432 77888
rect 75474 77848 75514 77888
rect 75556 77848 75596 77888
rect 75638 77848 75678 77888
rect 75720 77848 75760 77888
rect 90512 77848 90552 77888
rect 90594 77848 90634 77888
rect 90676 77848 90716 77888
rect 90758 77848 90798 77888
rect 90840 77848 90880 77888
rect 105632 77848 105672 77888
rect 105714 77848 105754 77888
rect 105796 77848 105836 77888
rect 105878 77848 105918 77888
rect 105960 77848 106000 77888
rect 120752 77848 120792 77888
rect 120834 77848 120874 77888
rect 120916 77848 120956 77888
rect 120998 77848 121038 77888
rect 121080 77848 121120 77888
rect 135872 77848 135912 77888
rect 135954 77848 135994 77888
rect 136036 77848 136076 77888
rect 136118 77848 136158 77888
rect 136200 77848 136240 77888
rect 150992 77848 151032 77888
rect 151074 77848 151114 77888
rect 151156 77848 151196 77888
rect 151238 77848 151278 77888
rect 151320 77848 151360 77888
rect 74152 77092 74192 77132
rect 74234 77092 74274 77132
rect 74316 77092 74356 77132
rect 74398 77092 74438 77132
rect 74480 77092 74520 77132
rect 89272 77092 89312 77132
rect 89354 77092 89394 77132
rect 89436 77092 89476 77132
rect 89518 77092 89558 77132
rect 89600 77092 89640 77132
rect 104392 77092 104432 77132
rect 104474 77092 104514 77132
rect 104556 77092 104596 77132
rect 104638 77092 104678 77132
rect 104720 77092 104760 77132
rect 119512 77092 119552 77132
rect 119594 77092 119634 77132
rect 119676 77092 119716 77132
rect 119758 77092 119798 77132
rect 119840 77092 119880 77132
rect 134632 77092 134672 77132
rect 134714 77092 134754 77132
rect 134796 77092 134836 77132
rect 134878 77092 134918 77132
rect 134960 77092 135000 77132
rect 149752 77092 149792 77132
rect 149834 77092 149874 77132
rect 149916 77092 149956 77132
rect 149998 77092 150038 77132
rect 150080 77092 150120 77132
rect 75392 76336 75432 76376
rect 75474 76336 75514 76376
rect 75556 76336 75596 76376
rect 75638 76336 75678 76376
rect 75720 76336 75760 76376
rect 90512 76336 90552 76376
rect 90594 76336 90634 76376
rect 90676 76336 90716 76376
rect 90758 76336 90798 76376
rect 90840 76336 90880 76376
rect 105632 76336 105672 76376
rect 105714 76336 105754 76376
rect 105796 76336 105836 76376
rect 105878 76336 105918 76376
rect 105960 76336 106000 76376
rect 120752 76336 120792 76376
rect 120834 76336 120874 76376
rect 120916 76336 120956 76376
rect 120998 76336 121038 76376
rect 121080 76336 121120 76376
rect 135872 76336 135912 76376
rect 135954 76336 135994 76376
rect 136036 76336 136076 76376
rect 136118 76336 136158 76376
rect 136200 76336 136240 76376
rect 150992 76336 151032 76376
rect 151074 76336 151114 76376
rect 151156 76336 151196 76376
rect 151238 76336 151278 76376
rect 151320 76336 151360 76376
rect 74152 75580 74192 75620
rect 74234 75580 74274 75620
rect 74316 75580 74356 75620
rect 74398 75580 74438 75620
rect 74480 75580 74520 75620
rect 89272 75580 89312 75620
rect 89354 75580 89394 75620
rect 89436 75580 89476 75620
rect 89518 75580 89558 75620
rect 89600 75580 89640 75620
rect 104392 75580 104432 75620
rect 104474 75580 104514 75620
rect 104556 75580 104596 75620
rect 104638 75580 104678 75620
rect 104720 75580 104760 75620
rect 119512 75580 119552 75620
rect 119594 75580 119634 75620
rect 119676 75580 119716 75620
rect 119758 75580 119798 75620
rect 119840 75580 119880 75620
rect 134632 75580 134672 75620
rect 134714 75580 134754 75620
rect 134796 75580 134836 75620
rect 134878 75580 134918 75620
rect 134960 75580 135000 75620
rect 149752 75580 149792 75620
rect 149834 75580 149874 75620
rect 149916 75580 149956 75620
rect 149998 75580 150038 75620
rect 150080 75580 150120 75620
rect 75392 74824 75432 74864
rect 75474 74824 75514 74864
rect 75556 74824 75596 74864
rect 75638 74824 75678 74864
rect 75720 74824 75760 74864
rect 90512 74824 90552 74864
rect 90594 74824 90634 74864
rect 90676 74824 90716 74864
rect 90758 74824 90798 74864
rect 90840 74824 90880 74864
rect 105632 74824 105672 74864
rect 105714 74824 105754 74864
rect 105796 74824 105836 74864
rect 105878 74824 105918 74864
rect 105960 74824 106000 74864
rect 120752 74824 120792 74864
rect 120834 74824 120874 74864
rect 120916 74824 120956 74864
rect 120998 74824 121038 74864
rect 121080 74824 121120 74864
rect 135872 74824 135912 74864
rect 135954 74824 135994 74864
rect 136036 74824 136076 74864
rect 136118 74824 136158 74864
rect 136200 74824 136240 74864
rect 150992 74824 151032 74864
rect 151074 74824 151114 74864
rect 151156 74824 151196 74864
rect 151238 74824 151278 74864
rect 151320 74824 151360 74864
rect 74152 74068 74192 74108
rect 74234 74068 74274 74108
rect 74316 74068 74356 74108
rect 74398 74068 74438 74108
rect 74480 74068 74520 74108
rect 89272 74068 89312 74108
rect 89354 74068 89394 74108
rect 89436 74068 89476 74108
rect 89518 74068 89558 74108
rect 89600 74068 89640 74108
rect 104392 74068 104432 74108
rect 104474 74068 104514 74108
rect 104556 74068 104596 74108
rect 104638 74068 104678 74108
rect 104720 74068 104760 74108
rect 119512 74068 119552 74108
rect 119594 74068 119634 74108
rect 119676 74068 119716 74108
rect 119758 74068 119798 74108
rect 119840 74068 119880 74108
rect 134632 74068 134672 74108
rect 134714 74068 134754 74108
rect 134796 74068 134836 74108
rect 134878 74068 134918 74108
rect 134960 74068 135000 74108
rect 149752 74068 149792 74108
rect 149834 74068 149874 74108
rect 149916 74068 149956 74108
rect 149998 74068 150038 74108
rect 150080 74068 150120 74108
rect 75392 73312 75432 73352
rect 75474 73312 75514 73352
rect 75556 73312 75596 73352
rect 75638 73312 75678 73352
rect 75720 73312 75760 73352
rect 90512 73312 90552 73352
rect 90594 73312 90634 73352
rect 90676 73312 90716 73352
rect 90758 73312 90798 73352
rect 90840 73312 90880 73352
rect 105632 73312 105672 73352
rect 105714 73312 105754 73352
rect 105796 73312 105836 73352
rect 105878 73312 105918 73352
rect 105960 73312 106000 73352
rect 120752 73312 120792 73352
rect 120834 73312 120874 73352
rect 120916 73312 120956 73352
rect 120998 73312 121038 73352
rect 121080 73312 121120 73352
rect 135872 73312 135912 73352
rect 135954 73312 135994 73352
rect 136036 73312 136076 73352
rect 136118 73312 136158 73352
rect 136200 73312 136240 73352
rect 150992 73312 151032 73352
rect 151074 73312 151114 73352
rect 151156 73312 151196 73352
rect 151238 73312 151278 73352
rect 151320 73312 151360 73352
rect 74152 72556 74192 72596
rect 74234 72556 74274 72596
rect 74316 72556 74356 72596
rect 74398 72556 74438 72596
rect 74480 72556 74520 72596
rect 89272 72556 89312 72596
rect 89354 72556 89394 72596
rect 89436 72556 89476 72596
rect 89518 72556 89558 72596
rect 89600 72556 89640 72596
rect 104392 72556 104432 72596
rect 104474 72556 104514 72596
rect 104556 72556 104596 72596
rect 104638 72556 104678 72596
rect 104720 72556 104760 72596
rect 119512 72556 119552 72596
rect 119594 72556 119634 72596
rect 119676 72556 119716 72596
rect 119758 72556 119798 72596
rect 119840 72556 119880 72596
rect 134632 72556 134672 72596
rect 134714 72556 134754 72596
rect 134796 72556 134836 72596
rect 134878 72556 134918 72596
rect 134960 72556 135000 72596
rect 149752 72556 149792 72596
rect 149834 72556 149874 72596
rect 149916 72556 149956 72596
rect 149998 72556 150038 72596
rect 150080 72556 150120 72596
rect 75392 71800 75432 71840
rect 75474 71800 75514 71840
rect 75556 71800 75596 71840
rect 75638 71800 75678 71840
rect 75720 71800 75760 71840
rect 90512 71800 90552 71840
rect 90594 71800 90634 71840
rect 90676 71800 90716 71840
rect 90758 71800 90798 71840
rect 90840 71800 90880 71840
rect 105632 71800 105672 71840
rect 105714 71800 105754 71840
rect 105796 71800 105836 71840
rect 105878 71800 105918 71840
rect 105960 71800 106000 71840
rect 120752 71800 120792 71840
rect 120834 71800 120874 71840
rect 120916 71800 120956 71840
rect 120998 71800 121038 71840
rect 121080 71800 121120 71840
rect 135872 71800 135912 71840
rect 135954 71800 135994 71840
rect 136036 71800 136076 71840
rect 136118 71800 136158 71840
rect 136200 71800 136240 71840
rect 150992 71800 151032 71840
rect 151074 71800 151114 71840
rect 151156 71800 151196 71840
rect 151238 71800 151278 71840
rect 151320 71800 151360 71840
<< metal4 >>
rect 75392 151976 75760 151985
rect 75432 151936 75474 151976
rect 75514 151936 75556 151976
rect 75596 151936 75638 151976
rect 75678 151936 75720 151976
rect 75392 151927 75760 151936
rect 90512 151976 90880 151985
rect 90552 151936 90594 151976
rect 90634 151936 90676 151976
rect 90716 151936 90758 151976
rect 90798 151936 90840 151976
rect 90512 151927 90880 151936
rect 105632 151976 106000 151985
rect 105672 151936 105714 151976
rect 105754 151936 105796 151976
rect 105836 151936 105878 151976
rect 105918 151936 105960 151976
rect 105632 151927 106000 151936
rect 120752 151976 121120 151985
rect 120792 151936 120834 151976
rect 120874 151936 120916 151976
rect 120956 151936 120998 151976
rect 121038 151936 121080 151976
rect 120752 151927 121120 151936
rect 135872 151976 136240 151985
rect 135912 151936 135954 151976
rect 135994 151936 136036 151976
rect 136076 151936 136118 151976
rect 136158 151936 136200 151976
rect 135872 151927 136240 151936
rect 150992 151976 151360 151985
rect 151032 151936 151074 151976
rect 151114 151936 151156 151976
rect 151196 151936 151238 151976
rect 151278 151936 151320 151976
rect 150992 151927 151360 151936
rect 74152 151220 74520 151229
rect 74192 151180 74234 151220
rect 74274 151180 74316 151220
rect 74356 151180 74398 151220
rect 74438 151180 74480 151220
rect 74152 151171 74520 151180
rect 89272 151220 89640 151229
rect 89312 151180 89354 151220
rect 89394 151180 89436 151220
rect 89476 151180 89518 151220
rect 89558 151180 89600 151220
rect 89272 151171 89640 151180
rect 104392 151220 104760 151229
rect 104432 151180 104474 151220
rect 104514 151180 104556 151220
rect 104596 151180 104638 151220
rect 104678 151180 104720 151220
rect 104392 151171 104760 151180
rect 119512 151220 119880 151229
rect 119552 151180 119594 151220
rect 119634 151180 119676 151220
rect 119716 151180 119758 151220
rect 119798 151180 119840 151220
rect 119512 151171 119880 151180
rect 134632 151220 135000 151229
rect 134672 151180 134714 151220
rect 134754 151180 134796 151220
rect 134836 151180 134878 151220
rect 134918 151180 134960 151220
rect 134632 151171 135000 151180
rect 149752 151220 150120 151229
rect 149792 151180 149834 151220
rect 149874 151180 149916 151220
rect 149956 151180 149998 151220
rect 150038 151180 150080 151220
rect 149752 151171 150120 151180
rect 75392 150464 75760 150473
rect 75432 150424 75474 150464
rect 75514 150424 75556 150464
rect 75596 150424 75638 150464
rect 75678 150424 75720 150464
rect 75392 150415 75760 150424
rect 90512 150464 90880 150473
rect 90552 150424 90594 150464
rect 90634 150424 90676 150464
rect 90716 150424 90758 150464
rect 90798 150424 90840 150464
rect 90512 150415 90880 150424
rect 105632 150464 106000 150473
rect 105672 150424 105714 150464
rect 105754 150424 105796 150464
rect 105836 150424 105878 150464
rect 105918 150424 105960 150464
rect 105632 150415 106000 150424
rect 120752 150464 121120 150473
rect 120792 150424 120834 150464
rect 120874 150424 120916 150464
rect 120956 150424 120998 150464
rect 121038 150424 121080 150464
rect 120752 150415 121120 150424
rect 135872 150464 136240 150473
rect 135912 150424 135954 150464
rect 135994 150424 136036 150464
rect 136076 150424 136118 150464
rect 136158 150424 136200 150464
rect 135872 150415 136240 150424
rect 150992 150464 151360 150473
rect 151032 150424 151074 150464
rect 151114 150424 151156 150464
rect 151196 150424 151238 150464
rect 151278 150424 151320 150464
rect 150992 150415 151360 150424
rect 74152 149708 74520 149717
rect 74192 149668 74234 149708
rect 74274 149668 74316 149708
rect 74356 149668 74398 149708
rect 74438 149668 74480 149708
rect 74152 149659 74520 149668
rect 89272 149708 89640 149717
rect 89312 149668 89354 149708
rect 89394 149668 89436 149708
rect 89476 149668 89518 149708
rect 89558 149668 89600 149708
rect 89272 149659 89640 149668
rect 104392 149708 104760 149717
rect 104432 149668 104474 149708
rect 104514 149668 104556 149708
rect 104596 149668 104638 149708
rect 104678 149668 104720 149708
rect 104392 149659 104760 149668
rect 119512 149708 119880 149717
rect 119552 149668 119594 149708
rect 119634 149668 119676 149708
rect 119716 149668 119758 149708
rect 119798 149668 119840 149708
rect 119512 149659 119880 149668
rect 134632 149708 135000 149717
rect 134672 149668 134714 149708
rect 134754 149668 134796 149708
rect 134836 149668 134878 149708
rect 134918 149668 134960 149708
rect 134632 149659 135000 149668
rect 149752 149708 150120 149717
rect 149792 149668 149834 149708
rect 149874 149668 149916 149708
rect 149956 149668 149998 149708
rect 150038 149668 150080 149708
rect 149752 149659 150120 149668
rect 75392 148952 75760 148961
rect 75432 148912 75474 148952
rect 75514 148912 75556 148952
rect 75596 148912 75638 148952
rect 75678 148912 75720 148952
rect 75392 148903 75760 148912
rect 90512 148952 90880 148961
rect 90552 148912 90594 148952
rect 90634 148912 90676 148952
rect 90716 148912 90758 148952
rect 90798 148912 90840 148952
rect 90512 148903 90880 148912
rect 105632 148952 106000 148961
rect 105672 148912 105714 148952
rect 105754 148912 105796 148952
rect 105836 148912 105878 148952
rect 105918 148912 105960 148952
rect 105632 148903 106000 148912
rect 120752 148952 121120 148961
rect 120792 148912 120834 148952
rect 120874 148912 120916 148952
rect 120956 148912 120998 148952
rect 121038 148912 121080 148952
rect 120752 148903 121120 148912
rect 135872 148952 136240 148961
rect 135912 148912 135954 148952
rect 135994 148912 136036 148952
rect 136076 148912 136118 148952
rect 136158 148912 136200 148952
rect 135872 148903 136240 148912
rect 150992 148952 151360 148961
rect 151032 148912 151074 148952
rect 151114 148912 151156 148952
rect 151196 148912 151238 148952
rect 151278 148912 151320 148952
rect 150992 148903 151360 148912
rect 74152 148196 74520 148205
rect 74192 148156 74234 148196
rect 74274 148156 74316 148196
rect 74356 148156 74398 148196
rect 74438 148156 74480 148196
rect 74152 148147 74520 148156
rect 89272 148196 89640 148205
rect 89312 148156 89354 148196
rect 89394 148156 89436 148196
rect 89476 148156 89518 148196
rect 89558 148156 89600 148196
rect 89272 148147 89640 148156
rect 104392 148196 104760 148205
rect 104432 148156 104474 148196
rect 104514 148156 104556 148196
rect 104596 148156 104638 148196
rect 104678 148156 104720 148196
rect 104392 148147 104760 148156
rect 119512 148196 119880 148205
rect 119552 148156 119594 148196
rect 119634 148156 119676 148196
rect 119716 148156 119758 148196
rect 119798 148156 119840 148196
rect 119512 148147 119880 148156
rect 134632 148196 135000 148205
rect 134672 148156 134714 148196
rect 134754 148156 134796 148196
rect 134836 148156 134878 148196
rect 134918 148156 134960 148196
rect 134632 148147 135000 148156
rect 149752 148196 150120 148205
rect 149792 148156 149834 148196
rect 149874 148156 149916 148196
rect 149956 148156 149998 148196
rect 150038 148156 150080 148196
rect 149752 148147 150120 148156
rect 75392 147440 75760 147449
rect 75432 147400 75474 147440
rect 75514 147400 75556 147440
rect 75596 147400 75638 147440
rect 75678 147400 75720 147440
rect 75392 147391 75760 147400
rect 90512 147440 90880 147449
rect 90552 147400 90594 147440
rect 90634 147400 90676 147440
rect 90716 147400 90758 147440
rect 90798 147400 90840 147440
rect 90512 147391 90880 147400
rect 105632 147440 106000 147449
rect 105672 147400 105714 147440
rect 105754 147400 105796 147440
rect 105836 147400 105878 147440
rect 105918 147400 105960 147440
rect 105632 147391 106000 147400
rect 120752 147440 121120 147449
rect 120792 147400 120834 147440
rect 120874 147400 120916 147440
rect 120956 147400 120998 147440
rect 121038 147400 121080 147440
rect 120752 147391 121120 147400
rect 135872 147440 136240 147449
rect 135912 147400 135954 147440
rect 135994 147400 136036 147440
rect 136076 147400 136118 147440
rect 136158 147400 136200 147440
rect 135872 147391 136240 147400
rect 150992 147440 151360 147449
rect 151032 147400 151074 147440
rect 151114 147400 151156 147440
rect 151196 147400 151238 147440
rect 151278 147400 151320 147440
rect 150992 147391 151360 147400
rect 74152 146684 74520 146693
rect 74192 146644 74234 146684
rect 74274 146644 74316 146684
rect 74356 146644 74398 146684
rect 74438 146644 74480 146684
rect 74152 146635 74520 146644
rect 89272 146684 89640 146693
rect 89312 146644 89354 146684
rect 89394 146644 89436 146684
rect 89476 146644 89518 146684
rect 89558 146644 89600 146684
rect 89272 146635 89640 146644
rect 104392 146684 104760 146693
rect 104432 146644 104474 146684
rect 104514 146644 104556 146684
rect 104596 146644 104638 146684
rect 104678 146644 104720 146684
rect 104392 146635 104760 146644
rect 119512 146684 119880 146693
rect 119552 146644 119594 146684
rect 119634 146644 119676 146684
rect 119716 146644 119758 146684
rect 119798 146644 119840 146684
rect 119512 146635 119880 146644
rect 134632 146684 135000 146693
rect 134672 146644 134714 146684
rect 134754 146644 134796 146684
rect 134836 146644 134878 146684
rect 134918 146644 134960 146684
rect 134632 146635 135000 146644
rect 149752 146684 150120 146693
rect 149792 146644 149834 146684
rect 149874 146644 149916 146684
rect 149956 146644 149998 146684
rect 150038 146644 150080 146684
rect 149752 146635 150120 146644
rect 75392 145928 75760 145937
rect 75432 145888 75474 145928
rect 75514 145888 75556 145928
rect 75596 145888 75638 145928
rect 75678 145888 75720 145928
rect 75392 145879 75760 145888
rect 90512 145928 90880 145937
rect 90552 145888 90594 145928
rect 90634 145888 90676 145928
rect 90716 145888 90758 145928
rect 90798 145888 90840 145928
rect 90512 145879 90880 145888
rect 105632 145928 106000 145937
rect 105672 145888 105714 145928
rect 105754 145888 105796 145928
rect 105836 145888 105878 145928
rect 105918 145888 105960 145928
rect 105632 145879 106000 145888
rect 120752 145928 121120 145937
rect 120792 145888 120834 145928
rect 120874 145888 120916 145928
rect 120956 145888 120998 145928
rect 121038 145888 121080 145928
rect 120752 145879 121120 145888
rect 135872 145928 136240 145937
rect 135912 145888 135954 145928
rect 135994 145888 136036 145928
rect 136076 145888 136118 145928
rect 136158 145888 136200 145928
rect 135872 145879 136240 145888
rect 150992 145928 151360 145937
rect 151032 145888 151074 145928
rect 151114 145888 151156 145928
rect 151196 145888 151238 145928
rect 151278 145888 151320 145928
rect 150992 145879 151360 145888
rect 74152 145172 74520 145181
rect 74192 145132 74234 145172
rect 74274 145132 74316 145172
rect 74356 145132 74398 145172
rect 74438 145132 74480 145172
rect 74152 145123 74520 145132
rect 89272 145172 89640 145181
rect 89312 145132 89354 145172
rect 89394 145132 89436 145172
rect 89476 145132 89518 145172
rect 89558 145132 89600 145172
rect 89272 145123 89640 145132
rect 104392 145172 104760 145181
rect 104432 145132 104474 145172
rect 104514 145132 104556 145172
rect 104596 145132 104638 145172
rect 104678 145132 104720 145172
rect 104392 145123 104760 145132
rect 119512 145172 119880 145181
rect 119552 145132 119594 145172
rect 119634 145132 119676 145172
rect 119716 145132 119758 145172
rect 119798 145132 119840 145172
rect 119512 145123 119880 145132
rect 134632 145172 135000 145181
rect 134672 145132 134714 145172
rect 134754 145132 134796 145172
rect 134836 145132 134878 145172
rect 134918 145132 134960 145172
rect 134632 145123 135000 145132
rect 149752 145172 150120 145181
rect 149792 145132 149834 145172
rect 149874 145132 149916 145172
rect 149956 145132 149998 145172
rect 150038 145132 150080 145172
rect 149752 145123 150120 145132
rect 75392 144416 75760 144425
rect 75432 144376 75474 144416
rect 75514 144376 75556 144416
rect 75596 144376 75638 144416
rect 75678 144376 75720 144416
rect 75392 144367 75760 144376
rect 90512 144416 90880 144425
rect 90552 144376 90594 144416
rect 90634 144376 90676 144416
rect 90716 144376 90758 144416
rect 90798 144376 90840 144416
rect 90512 144367 90880 144376
rect 105632 144416 106000 144425
rect 105672 144376 105714 144416
rect 105754 144376 105796 144416
rect 105836 144376 105878 144416
rect 105918 144376 105960 144416
rect 105632 144367 106000 144376
rect 120752 144416 121120 144425
rect 120792 144376 120834 144416
rect 120874 144376 120916 144416
rect 120956 144376 120998 144416
rect 121038 144376 121080 144416
rect 120752 144367 121120 144376
rect 135872 144416 136240 144425
rect 135912 144376 135954 144416
rect 135994 144376 136036 144416
rect 136076 144376 136118 144416
rect 136158 144376 136200 144416
rect 135872 144367 136240 144376
rect 150992 144416 151360 144425
rect 151032 144376 151074 144416
rect 151114 144376 151156 144416
rect 151196 144376 151238 144416
rect 151278 144376 151320 144416
rect 150992 144367 151360 144376
rect 74152 143660 74520 143669
rect 74192 143620 74234 143660
rect 74274 143620 74316 143660
rect 74356 143620 74398 143660
rect 74438 143620 74480 143660
rect 74152 143611 74520 143620
rect 89272 143660 89640 143669
rect 89312 143620 89354 143660
rect 89394 143620 89436 143660
rect 89476 143620 89518 143660
rect 89558 143620 89600 143660
rect 89272 143611 89640 143620
rect 104392 143660 104760 143669
rect 104432 143620 104474 143660
rect 104514 143620 104556 143660
rect 104596 143620 104638 143660
rect 104678 143620 104720 143660
rect 104392 143611 104760 143620
rect 119512 143660 119880 143669
rect 119552 143620 119594 143660
rect 119634 143620 119676 143660
rect 119716 143620 119758 143660
rect 119798 143620 119840 143660
rect 119512 143611 119880 143620
rect 134632 143660 135000 143669
rect 134672 143620 134714 143660
rect 134754 143620 134796 143660
rect 134836 143620 134878 143660
rect 134918 143620 134960 143660
rect 134632 143611 135000 143620
rect 149752 143660 150120 143669
rect 149792 143620 149834 143660
rect 149874 143620 149916 143660
rect 149956 143620 149998 143660
rect 150038 143620 150080 143660
rect 149752 143611 150120 143620
rect 75392 142904 75760 142913
rect 75432 142864 75474 142904
rect 75514 142864 75556 142904
rect 75596 142864 75638 142904
rect 75678 142864 75720 142904
rect 75392 142855 75760 142864
rect 90512 142904 90880 142913
rect 90552 142864 90594 142904
rect 90634 142864 90676 142904
rect 90716 142864 90758 142904
rect 90798 142864 90840 142904
rect 90512 142855 90880 142864
rect 105632 142904 106000 142913
rect 105672 142864 105714 142904
rect 105754 142864 105796 142904
rect 105836 142864 105878 142904
rect 105918 142864 105960 142904
rect 105632 142855 106000 142864
rect 120752 142904 121120 142913
rect 120792 142864 120834 142904
rect 120874 142864 120916 142904
rect 120956 142864 120998 142904
rect 121038 142864 121080 142904
rect 120752 142855 121120 142864
rect 135872 142904 136240 142913
rect 135912 142864 135954 142904
rect 135994 142864 136036 142904
rect 136076 142864 136118 142904
rect 136158 142864 136200 142904
rect 135872 142855 136240 142864
rect 150992 142904 151360 142913
rect 151032 142864 151074 142904
rect 151114 142864 151156 142904
rect 151196 142864 151238 142904
rect 151278 142864 151320 142904
rect 150992 142855 151360 142864
rect 74152 142148 74520 142157
rect 74192 142108 74234 142148
rect 74274 142108 74316 142148
rect 74356 142108 74398 142148
rect 74438 142108 74480 142148
rect 74152 142099 74520 142108
rect 89272 142148 89640 142157
rect 89312 142108 89354 142148
rect 89394 142108 89436 142148
rect 89476 142108 89518 142148
rect 89558 142108 89600 142148
rect 89272 142099 89640 142108
rect 104392 142148 104760 142157
rect 104432 142108 104474 142148
rect 104514 142108 104556 142148
rect 104596 142108 104638 142148
rect 104678 142108 104720 142148
rect 104392 142099 104760 142108
rect 119512 142148 119880 142157
rect 119552 142108 119594 142148
rect 119634 142108 119676 142148
rect 119716 142108 119758 142148
rect 119798 142108 119840 142148
rect 119512 142099 119880 142108
rect 134632 142148 135000 142157
rect 134672 142108 134714 142148
rect 134754 142108 134796 142148
rect 134836 142108 134878 142148
rect 134918 142108 134960 142148
rect 134632 142099 135000 142108
rect 149752 142148 150120 142157
rect 149792 142108 149834 142148
rect 149874 142108 149916 142148
rect 149956 142108 149998 142148
rect 150038 142108 150080 142148
rect 149752 142099 150120 142108
rect 75392 141392 75760 141401
rect 75432 141352 75474 141392
rect 75514 141352 75556 141392
rect 75596 141352 75638 141392
rect 75678 141352 75720 141392
rect 75392 141343 75760 141352
rect 90512 141392 90880 141401
rect 90552 141352 90594 141392
rect 90634 141352 90676 141392
rect 90716 141352 90758 141392
rect 90798 141352 90840 141392
rect 90512 141343 90880 141352
rect 105632 141392 106000 141401
rect 105672 141352 105714 141392
rect 105754 141352 105796 141392
rect 105836 141352 105878 141392
rect 105918 141352 105960 141392
rect 105632 141343 106000 141352
rect 120752 141392 121120 141401
rect 120792 141352 120834 141392
rect 120874 141352 120916 141392
rect 120956 141352 120998 141392
rect 121038 141352 121080 141392
rect 120752 141343 121120 141352
rect 135872 141392 136240 141401
rect 135912 141352 135954 141392
rect 135994 141352 136036 141392
rect 136076 141352 136118 141392
rect 136158 141352 136200 141392
rect 135872 141343 136240 141352
rect 150992 141392 151360 141401
rect 151032 141352 151074 141392
rect 151114 141352 151156 141392
rect 151196 141352 151238 141392
rect 151278 141352 151320 141392
rect 150992 141343 151360 141352
rect 74152 140636 74520 140645
rect 74192 140596 74234 140636
rect 74274 140596 74316 140636
rect 74356 140596 74398 140636
rect 74438 140596 74480 140636
rect 74152 140587 74520 140596
rect 89272 140636 89640 140645
rect 89312 140596 89354 140636
rect 89394 140596 89436 140636
rect 89476 140596 89518 140636
rect 89558 140596 89600 140636
rect 89272 140587 89640 140596
rect 104392 140636 104760 140645
rect 104432 140596 104474 140636
rect 104514 140596 104556 140636
rect 104596 140596 104638 140636
rect 104678 140596 104720 140636
rect 104392 140587 104760 140596
rect 119512 140636 119880 140645
rect 119552 140596 119594 140636
rect 119634 140596 119676 140636
rect 119716 140596 119758 140636
rect 119798 140596 119840 140636
rect 119512 140587 119880 140596
rect 134632 140636 135000 140645
rect 134672 140596 134714 140636
rect 134754 140596 134796 140636
rect 134836 140596 134878 140636
rect 134918 140596 134960 140636
rect 134632 140587 135000 140596
rect 149752 140636 150120 140645
rect 149792 140596 149834 140636
rect 149874 140596 149916 140636
rect 149956 140596 149998 140636
rect 150038 140596 150080 140636
rect 149752 140587 150120 140596
rect 75392 139880 75760 139889
rect 75432 139840 75474 139880
rect 75514 139840 75556 139880
rect 75596 139840 75638 139880
rect 75678 139840 75720 139880
rect 75392 139831 75760 139840
rect 90512 139880 90880 139889
rect 90552 139840 90594 139880
rect 90634 139840 90676 139880
rect 90716 139840 90758 139880
rect 90798 139840 90840 139880
rect 90512 139831 90880 139840
rect 105632 139880 106000 139889
rect 105672 139840 105714 139880
rect 105754 139840 105796 139880
rect 105836 139840 105878 139880
rect 105918 139840 105960 139880
rect 105632 139831 106000 139840
rect 120752 139880 121120 139889
rect 120792 139840 120834 139880
rect 120874 139840 120916 139880
rect 120956 139840 120998 139880
rect 121038 139840 121080 139880
rect 120752 139831 121120 139840
rect 135872 139880 136240 139889
rect 135912 139840 135954 139880
rect 135994 139840 136036 139880
rect 136076 139840 136118 139880
rect 136158 139840 136200 139880
rect 135872 139831 136240 139840
rect 150992 139880 151360 139889
rect 151032 139840 151074 139880
rect 151114 139840 151156 139880
rect 151196 139840 151238 139880
rect 151278 139840 151320 139880
rect 150992 139831 151360 139840
rect 74152 139124 74520 139133
rect 74192 139084 74234 139124
rect 74274 139084 74316 139124
rect 74356 139084 74398 139124
rect 74438 139084 74480 139124
rect 74152 139075 74520 139084
rect 89272 139124 89640 139133
rect 89312 139084 89354 139124
rect 89394 139084 89436 139124
rect 89476 139084 89518 139124
rect 89558 139084 89600 139124
rect 89272 139075 89640 139084
rect 104392 139124 104760 139133
rect 104432 139084 104474 139124
rect 104514 139084 104556 139124
rect 104596 139084 104638 139124
rect 104678 139084 104720 139124
rect 104392 139075 104760 139084
rect 119512 139124 119880 139133
rect 119552 139084 119594 139124
rect 119634 139084 119676 139124
rect 119716 139084 119758 139124
rect 119798 139084 119840 139124
rect 119512 139075 119880 139084
rect 134632 139124 135000 139133
rect 134672 139084 134714 139124
rect 134754 139084 134796 139124
rect 134836 139084 134878 139124
rect 134918 139084 134960 139124
rect 134632 139075 135000 139084
rect 149752 139124 150120 139133
rect 149792 139084 149834 139124
rect 149874 139084 149916 139124
rect 149956 139084 149998 139124
rect 150038 139084 150080 139124
rect 149752 139075 150120 139084
rect 75392 138368 75760 138377
rect 75432 138328 75474 138368
rect 75514 138328 75556 138368
rect 75596 138328 75638 138368
rect 75678 138328 75720 138368
rect 75392 138319 75760 138328
rect 90512 138368 90880 138377
rect 90552 138328 90594 138368
rect 90634 138328 90676 138368
rect 90716 138328 90758 138368
rect 90798 138328 90840 138368
rect 90512 138319 90880 138328
rect 105632 138368 106000 138377
rect 105672 138328 105714 138368
rect 105754 138328 105796 138368
rect 105836 138328 105878 138368
rect 105918 138328 105960 138368
rect 105632 138319 106000 138328
rect 120752 138368 121120 138377
rect 120792 138328 120834 138368
rect 120874 138328 120916 138368
rect 120956 138328 120998 138368
rect 121038 138328 121080 138368
rect 120752 138319 121120 138328
rect 135872 138368 136240 138377
rect 135912 138328 135954 138368
rect 135994 138328 136036 138368
rect 136076 138328 136118 138368
rect 136158 138328 136200 138368
rect 135872 138319 136240 138328
rect 150992 138368 151360 138377
rect 151032 138328 151074 138368
rect 151114 138328 151156 138368
rect 151196 138328 151238 138368
rect 151278 138328 151320 138368
rect 150992 138319 151360 138328
rect 74152 137612 74520 137621
rect 74192 137572 74234 137612
rect 74274 137572 74316 137612
rect 74356 137572 74398 137612
rect 74438 137572 74480 137612
rect 74152 137563 74520 137572
rect 89272 137612 89640 137621
rect 89312 137572 89354 137612
rect 89394 137572 89436 137612
rect 89476 137572 89518 137612
rect 89558 137572 89600 137612
rect 89272 137563 89640 137572
rect 104392 137612 104760 137621
rect 104432 137572 104474 137612
rect 104514 137572 104556 137612
rect 104596 137572 104638 137612
rect 104678 137572 104720 137612
rect 104392 137563 104760 137572
rect 119512 137612 119880 137621
rect 119552 137572 119594 137612
rect 119634 137572 119676 137612
rect 119716 137572 119758 137612
rect 119798 137572 119840 137612
rect 119512 137563 119880 137572
rect 134632 137612 135000 137621
rect 134672 137572 134714 137612
rect 134754 137572 134796 137612
rect 134836 137572 134878 137612
rect 134918 137572 134960 137612
rect 134632 137563 135000 137572
rect 149752 137612 150120 137621
rect 149792 137572 149834 137612
rect 149874 137572 149916 137612
rect 149956 137572 149998 137612
rect 150038 137572 150080 137612
rect 149752 137563 150120 137572
rect 75392 136856 75760 136865
rect 75432 136816 75474 136856
rect 75514 136816 75556 136856
rect 75596 136816 75638 136856
rect 75678 136816 75720 136856
rect 75392 136807 75760 136816
rect 90512 136856 90880 136865
rect 90552 136816 90594 136856
rect 90634 136816 90676 136856
rect 90716 136816 90758 136856
rect 90798 136816 90840 136856
rect 90512 136807 90880 136816
rect 105632 136856 106000 136865
rect 105672 136816 105714 136856
rect 105754 136816 105796 136856
rect 105836 136816 105878 136856
rect 105918 136816 105960 136856
rect 105632 136807 106000 136816
rect 120752 136856 121120 136865
rect 120792 136816 120834 136856
rect 120874 136816 120916 136856
rect 120956 136816 120998 136856
rect 121038 136816 121080 136856
rect 120752 136807 121120 136816
rect 135872 136856 136240 136865
rect 135912 136816 135954 136856
rect 135994 136816 136036 136856
rect 136076 136816 136118 136856
rect 136158 136816 136200 136856
rect 135872 136807 136240 136816
rect 150992 136856 151360 136865
rect 151032 136816 151074 136856
rect 151114 136816 151156 136856
rect 151196 136816 151238 136856
rect 151278 136816 151320 136856
rect 150992 136807 151360 136816
rect 74152 136100 74520 136109
rect 74192 136060 74234 136100
rect 74274 136060 74316 136100
rect 74356 136060 74398 136100
rect 74438 136060 74480 136100
rect 74152 136051 74520 136060
rect 89272 136100 89640 136109
rect 89312 136060 89354 136100
rect 89394 136060 89436 136100
rect 89476 136060 89518 136100
rect 89558 136060 89600 136100
rect 89272 136051 89640 136060
rect 104392 136100 104760 136109
rect 104432 136060 104474 136100
rect 104514 136060 104556 136100
rect 104596 136060 104638 136100
rect 104678 136060 104720 136100
rect 104392 136051 104760 136060
rect 119512 136100 119880 136109
rect 119552 136060 119594 136100
rect 119634 136060 119676 136100
rect 119716 136060 119758 136100
rect 119798 136060 119840 136100
rect 119512 136051 119880 136060
rect 134632 136100 135000 136109
rect 134672 136060 134714 136100
rect 134754 136060 134796 136100
rect 134836 136060 134878 136100
rect 134918 136060 134960 136100
rect 134632 136051 135000 136060
rect 149752 136100 150120 136109
rect 149792 136060 149834 136100
rect 149874 136060 149916 136100
rect 149956 136060 149998 136100
rect 150038 136060 150080 136100
rect 149752 136051 150120 136060
rect 75392 135344 75760 135353
rect 75432 135304 75474 135344
rect 75514 135304 75556 135344
rect 75596 135304 75638 135344
rect 75678 135304 75720 135344
rect 75392 135295 75760 135304
rect 90512 135344 90880 135353
rect 90552 135304 90594 135344
rect 90634 135304 90676 135344
rect 90716 135304 90758 135344
rect 90798 135304 90840 135344
rect 90512 135295 90880 135304
rect 105632 135344 106000 135353
rect 105672 135304 105714 135344
rect 105754 135304 105796 135344
rect 105836 135304 105878 135344
rect 105918 135304 105960 135344
rect 105632 135295 106000 135304
rect 120752 135344 121120 135353
rect 120792 135304 120834 135344
rect 120874 135304 120916 135344
rect 120956 135304 120998 135344
rect 121038 135304 121080 135344
rect 120752 135295 121120 135304
rect 135872 135344 136240 135353
rect 135912 135304 135954 135344
rect 135994 135304 136036 135344
rect 136076 135304 136118 135344
rect 136158 135304 136200 135344
rect 135872 135295 136240 135304
rect 150992 135344 151360 135353
rect 151032 135304 151074 135344
rect 151114 135304 151156 135344
rect 151196 135304 151238 135344
rect 151278 135304 151320 135344
rect 150992 135295 151360 135304
rect 74152 134588 74520 134597
rect 74192 134548 74234 134588
rect 74274 134548 74316 134588
rect 74356 134548 74398 134588
rect 74438 134548 74480 134588
rect 74152 134539 74520 134548
rect 89272 134588 89640 134597
rect 89312 134548 89354 134588
rect 89394 134548 89436 134588
rect 89476 134548 89518 134588
rect 89558 134548 89600 134588
rect 89272 134539 89640 134548
rect 104392 134588 104760 134597
rect 104432 134548 104474 134588
rect 104514 134548 104556 134588
rect 104596 134548 104638 134588
rect 104678 134548 104720 134588
rect 104392 134539 104760 134548
rect 119512 134588 119880 134597
rect 119552 134548 119594 134588
rect 119634 134548 119676 134588
rect 119716 134548 119758 134588
rect 119798 134548 119840 134588
rect 119512 134539 119880 134548
rect 134632 134588 135000 134597
rect 134672 134548 134714 134588
rect 134754 134548 134796 134588
rect 134836 134548 134878 134588
rect 134918 134548 134960 134588
rect 134632 134539 135000 134548
rect 149752 134588 150120 134597
rect 149792 134548 149834 134588
rect 149874 134548 149916 134588
rect 149956 134548 149998 134588
rect 150038 134548 150080 134588
rect 149752 134539 150120 134548
rect 75392 133832 75760 133841
rect 75432 133792 75474 133832
rect 75514 133792 75556 133832
rect 75596 133792 75638 133832
rect 75678 133792 75720 133832
rect 75392 133783 75760 133792
rect 90512 133832 90880 133841
rect 90552 133792 90594 133832
rect 90634 133792 90676 133832
rect 90716 133792 90758 133832
rect 90798 133792 90840 133832
rect 90512 133783 90880 133792
rect 105632 133832 106000 133841
rect 105672 133792 105714 133832
rect 105754 133792 105796 133832
rect 105836 133792 105878 133832
rect 105918 133792 105960 133832
rect 105632 133783 106000 133792
rect 120752 133832 121120 133841
rect 120792 133792 120834 133832
rect 120874 133792 120916 133832
rect 120956 133792 120998 133832
rect 121038 133792 121080 133832
rect 120752 133783 121120 133792
rect 135872 133832 136240 133841
rect 135912 133792 135954 133832
rect 135994 133792 136036 133832
rect 136076 133792 136118 133832
rect 136158 133792 136200 133832
rect 135872 133783 136240 133792
rect 150992 133832 151360 133841
rect 151032 133792 151074 133832
rect 151114 133792 151156 133832
rect 151196 133792 151238 133832
rect 151278 133792 151320 133832
rect 150992 133783 151360 133792
rect 74152 133076 74520 133085
rect 74192 133036 74234 133076
rect 74274 133036 74316 133076
rect 74356 133036 74398 133076
rect 74438 133036 74480 133076
rect 74152 133027 74520 133036
rect 89272 133076 89640 133085
rect 89312 133036 89354 133076
rect 89394 133036 89436 133076
rect 89476 133036 89518 133076
rect 89558 133036 89600 133076
rect 89272 133027 89640 133036
rect 104392 133076 104760 133085
rect 104432 133036 104474 133076
rect 104514 133036 104556 133076
rect 104596 133036 104638 133076
rect 104678 133036 104720 133076
rect 104392 133027 104760 133036
rect 119512 133076 119880 133085
rect 119552 133036 119594 133076
rect 119634 133036 119676 133076
rect 119716 133036 119758 133076
rect 119798 133036 119840 133076
rect 119512 133027 119880 133036
rect 134632 133076 135000 133085
rect 134672 133036 134714 133076
rect 134754 133036 134796 133076
rect 134836 133036 134878 133076
rect 134918 133036 134960 133076
rect 134632 133027 135000 133036
rect 149752 133076 150120 133085
rect 149792 133036 149834 133076
rect 149874 133036 149916 133076
rect 149956 133036 149998 133076
rect 150038 133036 150080 133076
rect 149752 133027 150120 133036
rect 75392 132320 75760 132329
rect 75432 132280 75474 132320
rect 75514 132280 75556 132320
rect 75596 132280 75638 132320
rect 75678 132280 75720 132320
rect 75392 132271 75760 132280
rect 90512 132320 90880 132329
rect 90552 132280 90594 132320
rect 90634 132280 90676 132320
rect 90716 132280 90758 132320
rect 90798 132280 90840 132320
rect 90512 132271 90880 132280
rect 105632 132320 106000 132329
rect 105672 132280 105714 132320
rect 105754 132280 105796 132320
rect 105836 132280 105878 132320
rect 105918 132280 105960 132320
rect 105632 132271 106000 132280
rect 120752 132320 121120 132329
rect 120792 132280 120834 132320
rect 120874 132280 120916 132320
rect 120956 132280 120998 132320
rect 121038 132280 121080 132320
rect 120752 132271 121120 132280
rect 135872 132320 136240 132329
rect 135912 132280 135954 132320
rect 135994 132280 136036 132320
rect 136076 132280 136118 132320
rect 136158 132280 136200 132320
rect 135872 132271 136240 132280
rect 150992 132320 151360 132329
rect 151032 132280 151074 132320
rect 151114 132280 151156 132320
rect 151196 132280 151238 132320
rect 151278 132280 151320 132320
rect 150992 132271 151360 132280
rect 74152 131564 74520 131573
rect 74192 131524 74234 131564
rect 74274 131524 74316 131564
rect 74356 131524 74398 131564
rect 74438 131524 74480 131564
rect 74152 131515 74520 131524
rect 89272 131564 89640 131573
rect 89312 131524 89354 131564
rect 89394 131524 89436 131564
rect 89476 131524 89518 131564
rect 89558 131524 89600 131564
rect 89272 131515 89640 131524
rect 104392 131564 104760 131573
rect 104432 131524 104474 131564
rect 104514 131524 104556 131564
rect 104596 131524 104638 131564
rect 104678 131524 104720 131564
rect 104392 131515 104760 131524
rect 119512 131564 119880 131573
rect 119552 131524 119594 131564
rect 119634 131524 119676 131564
rect 119716 131524 119758 131564
rect 119798 131524 119840 131564
rect 119512 131515 119880 131524
rect 134632 131564 135000 131573
rect 134672 131524 134714 131564
rect 134754 131524 134796 131564
rect 134836 131524 134878 131564
rect 134918 131524 134960 131564
rect 134632 131515 135000 131524
rect 149752 131564 150120 131573
rect 149792 131524 149834 131564
rect 149874 131524 149916 131564
rect 149956 131524 149998 131564
rect 150038 131524 150080 131564
rect 149752 131515 150120 131524
rect 75392 130808 75760 130817
rect 75432 130768 75474 130808
rect 75514 130768 75556 130808
rect 75596 130768 75638 130808
rect 75678 130768 75720 130808
rect 75392 130759 75760 130768
rect 90512 130808 90880 130817
rect 90552 130768 90594 130808
rect 90634 130768 90676 130808
rect 90716 130768 90758 130808
rect 90798 130768 90840 130808
rect 90512 130759 90880 130768
rect 105632 130808 106000 130817
rect 105672 130768 105714 130808
rect 105754 130768 105796 130808
rect 105836 130768 105878 130808
rect 105918 130768 105960 130808
rect 105632 130759 106000 130768
rect 120752 130808 121120 130817
rect 120792 130768 120834 130808
rect 120874 130768 120916 130808
rect 120956 130768 120998 130808
rect 121038 130768 121080 130808
rect 120752 130759 121120 130768
rect 135872 130808 136240 130817
rect 135912 130768 135954 130808
rect 135994 130768 136036 130808
rect 136076 130768 136118 130808
rect 136158 130768 136200 130808
rect 135872 130759 136240 130768
rect 150992 130808 151360 130817
rect 151032 130768 151074 130808
rect 151114 130768 151156 130808
rect 151196 130768 151238 130808
rect 151278 130768 151320 130808
rect 150992 130759 151360 130768
rect 74152 130052 74520 130061
rect 74192 130012 74234 130052
rect 74274 130012 74316 130052
rect 74356 130012 74398 130052
rect 74438 130012 74480 130052
rect 74152 130003 74520 130012
rect 89272 130052 89640 130061
rect 89312 130012 89354 130052
rect 89394 130012 89436 130052
rect 89476 130012 89518 130052
rect 89558 130012 89600 130052
rect 89272 130003 89640 130012
rect 104392 130052 104760 130061
rect 104432 130012 104474 130052
rect 104514 130012 104556 130052
rect 104596 130012 104638 130052
rect 104678 130012 104720 130052
rect 104392 130003 104760 130012
rect 119512 130052 119880 130061
rect 119552 130012 119594 130052
rect 119634 130012 119676 130052
rect 119716 130012 119758 130052
rect 119798 130012 119840 130052
rect 119512 130003 119880 130012
rect 134632 130052 135000 130061
rect 134672 130012 134714 130052
rect 134754 130012 134796 130052
rect 134836 130012 134878 130052
rect 134918 130012 134960 130052
rect 134632 130003 135000 130012
rect 149752 130052 150120 130061
rect 149792 130012 149834 130052
rect 149874 130012 149916 130052
rect 149956 130012 149998 130052
rect 150038 130012 150080 130052
rect 149752 130003 150120 130012
rect 75392 129296 75760 129305
rect 75432 129256 75474 129296
rect 75514 129256 75556 129296
rect 75596 129256 75638 129296
rect 75678 129256 75720 129296
rect 75392 129247 75760 129256
rect 90512 129296 90880 129305
rect 90552 129256 90594 129296
rect 90634 129256 90676 129296
rect 90716 129256 90758 129296
rect 90798 129256 90840 129296
rect 90512 129247 90880 129256
rect 105632 129296 106000 129305
rect 105672 129256 105714 129296
rect 105754 129256 105796 129296
rect 105836 129256 105878 129296
rect 105918 129256 105960 129296
rect 105632 129247 106000 129256
rect 120752 129296 121120 129305
rect 120792 129256 120834 129296
rect 120874 129256 120916 129296
rect 120956 129256 120998 129296
rect 121038 129256 121080 129296
rect 120752 129247 121120 129256
rect 135872 129296 136240 129305
rect 135912 129256 135954 129296
rect 135994 129256 136036 129296
rect 136076 129256 136118 129296
rect 136158 129256 136200 129296
rect 135872 129247 136240 129256
rect 150992 129296 151360 129305
rect 151032 129256 151074 129296
rect 151114 129256 151156 129296
rect 151196 129256 151238 129296
rect 151278 129256 151320 129296
rect 150992 129247 151360 129256
rect 74152 128540 74520 128549
rect 74192 128500 74234 128540
rect 74274 128500 74316 128540
rect 74356 128500 74398 128540
rect 74438 128500 74480 128540
rect 74152 128491 74520 128500
rect 89272 128540 89640 128549
rect 89312 128500 89354 128540
rect 89394 128500 89436 128540
rect 89476 128500 89518 128540
rect 89558 128500 89600 128540
rect 89272 128491 89640 128500
rect 104392 128540 104760 128549
rect 104432 128500 104474 128540
rect 104514 128500 104556 128540
rect 104596 128500 104638 128540
rect 104678 128500 104720 128540
rect 104392 128491 104760 128500
rect 119512 128540 119880 128549
rect 119552 128500 119594 128540
rect 119634 128500 119676 128540
rect 119716 128500 119758 128540
rect 119798 128500 119840 128540
rect 119512 128491 119880 128500
rect 134632 128540 135000 128549
rect 134672 128500 134714 128540
rect 134754 128500 134796 128540
rect 134836 128500 134878 128540
rect 134918 128500 134960 128540
rect 134632 128491 135000 128500
rect 149752 128540 150120 128549
rect 149792 128500 149834 128540
rect 149874 128500 149916 128540
rect 149956 128500 149998 128540
rect 150038 128500 150080 128540
rect 149752 128491 150120 128500
rect 75392 127784 75760 127793
rect 75432 127744 75474 127784
rect 75514 127744 75556 127784
rect 75596 127744 75638 127784
rect 75678 127744 75720 127784
rect 75392 127735 75760 127744
rect 90512 127784 90880 127793
rect 90552 127744 90594 127784
rect 90634 127744 90676 127784
rect 90716 127744 90758 127784
rect 90798 127744 90840 127784
rect 90512 127735 90880 127744
rect 105632 127784 106000 127793
rect 105672 127744 105714 127784
rect 105754 127744 105796 127784
rect 105836 127744 105878 127784
rect 105918 127744 105960 127784
rect 105632 127735 106000 127744
rect 120752 127784 121120 127793
rect 120792 127744 120834 127784
rect 120874 127744 120916 127784
rect 120956 127744 120998 127784
rect 121038 127744 121080 127784
rect 120752 127735 121120 127744
rect 135872 127784 136240 127793
rect 135912 127744 135954 127784
rect 135994 127744 136036 127784
rect 136076 127744 136118 127784
rect 136158 127744 136200 127784
rect 135872 127735 136240 127744
rect 150992 127784 151360 127793
rect 151032 127744 151074 127784
rect 151114 127744 151156 127784
rect 151196 127744 151238 127784
rect 151278 127744 151320 127784
rect 150992 127735 151360 127744
rect 74152 127028 74520 127037
rect 74192 126988 74234 127028
rect 74274 126988 74316 127028
rect 74356 126988 74398 127028
rect 74438 126988 74480 127028
rect 74152 126979 74520 126988
rect 89272 127028 89640 127037
rect 89312 126988 89354 127028
rect 89394 126988 89436 127028
rect 89476 126988 89518 127028
rect 89558 126988 89600 127028
rect 89272 126979 89640 126988
rect 104392 127028 104760 127037
rect 104432 126988 104474 127028
rect 104514 126988 104556 127028
rect 104596 126988 104638 127028
rect 104678 126988 104720 127028
rect 104392 126979 104760 126988
rect 119512 127028 119880 127037
rect 119552 126988 119594 127028
rect 119634 126988 119676 127028
rect 119716 126988 119758 127028
rect 119798 126988 119840 127028
rect 119512 126979 119880 126988
rect 134632 127028 135000 127037
rect 134672 126988 134714 127028
rect 134754 126988 134796 127028
rect 134836 126988 134878 127028
rect 134918 126988 134960 127028
rect 134632 126979 135000 126988
rect 149752 127028 150120 127037
rect 149792 126988 149834 127028
rect 149874 126988 149916 127028
rect 149956 126988 149998 127028
rect 150038 126988 150080 127028
rect 149752 126979 150120 126988
rect 75392 126272 75760 126281
rect 75432 126232 75474 126272
rect 75514 126232 75556 126272
rect 75596 126232 75638 126272
rect 75678 126232 75720 126272
rect 75392 126223 75760 126232
rect 90512 126272 90880 126281
rect 90552 126232 90594 126272
rect 90634 126232 90676 126272
rect 90716 126232 90758 126272
rect 90798 126232 90840 126272
rect 90512 126223 90880 126232
rect 105632 126272 106000 126281
rect 105672 126232 105714 126272
rect 105754 126232 105796 126272
rect 105836 126232 105878 126272
rect 105918 126232 105960 126272
rect 105632 126223 106000 126232
rect 120752 126272 121120 126281
rect 120792 126232 120834 126272
rect 120874 126232 120916 126272
rect 120956 126232 120998 126272
rect 121038 126232 121080 126272
rect 120752 126223 121120 126232
rect 135872 126272 136240 126281
rect 135912 126232 135954 126272
rect 135994 126232 136036 126272
rect 136076 126232 136118 126272
rect 136158 126232 136200 126272
rect 135872 126223 136240 126232
rect 150992 126272 151360 126281
rect 151032 126232 151074 126272
rect 151114 126232 151156 126272
rect 151196 126232 151238 126272
rect 151278 126232 151320 126272
rect 150992 126223 151360 126232
rect 74152 125516 74520 125525
rect 74192 125476 74234 125516
rect 74274 125476 74316 125516
rect 74356 125476 74398 125516
rect 74438 125476 74480 125516
rect 74152 125467 74520 125476
rect 89272 125516 89640 125525
rect 89312 125476 89354 125516
rect 89394 125476 89436 125516
rect 89476 125476 89518 125516
rect 89558 125476 89600 125516
rect 89272 125467 89640 125476
rect 104392 125516 104760 125525
rect 104432 125476 104474 125516
rect 104514 125476 104556 125516
rect 104596 125476 104638 125516
rect 104678 125476 104720 125516
rect 104392 125467 104760 125476
rect 119512 125516 119880 125525
rect 119552 125476 119594 125516
rect 119634 125476 119676 125516
rect 119716 125476 119758 125516
rect 119798 125476 119840 125516
rect 119512 125467 119880 125476
rect 134632 125516 135000 125525
rect 134672 125476 134714 125516
rect 134754 125476 134796 125516
rect 134836 125476 134878 125516
rect 134918 125476 134960 125516
rect 134632 125467 135000 125476
rect 149752 125516 150120 125525
rect 149792 125476 149834 125516
rect 149874 125476 149916 125516
rect 149956 125476 149998 125516
rect 150038 125476 150080 125516
rect 149752 125467 150120 125476
rect 75392 124760 75760 124769
rect 75432 124720 75474 124760
rect 75514 124720 75556 124760
rect 75596 124720 75638 124760
rect 75678 124720 75720 124760
rect 75392 124711 75760 124720
rect 90512 124760 90880 124769
rect 90552 124720 90594 124760
rect 90634 124720 90676 124760
rect 90716 124720 90758 124760
rect 90798 124720 90840 124760
rect 90512 124711 90880 124720
rect 105632 124760 106000 124769
rect 105672 124720 105714 124760
rect 105754 124720 105796 124760
rect 105836 124720 105878 124760
rect 105918 124720 105960 124760
rect 105632 124711 106000 124720
rect 120752 124760 121120 124769
rect 120792 124720 120834 124760
rect 120874 124720 120916 124760
rect 120956 124720 120998 124760
rect 121038 124720 121080 124760
rect 120752 124711 121120 124720
rect 135872 124760 136240 124769
rect 135912 124720 135954 124760
rect 135994 124720 136036 124760
rect 136076 124720 136118 124760
rect 136158 124720 136200 124760
rect 135872 124711 136240 124720
rect 150992 124760 151360 124769
rect 151032 124720 151074 124760
rect 151114 124720 151156 124760
rect 151196 124720 151238 124760
rect 151278 124720 151320 124760
rect 150992 124711 151360 124720
rect 74152 124004 74520 124013
rect 74192 123964 74234 124004
rect 74274 123964 74316 124004
rect 74356 123964 74398 124004
rect 74438 123964 74480 124004
rect 74152 123955 74520 123964
rect 89272 124004 89640 124013
rect 89312 123964 89354 124004
rect 89394 123964 89436 124004
rect 89476 123964 89518 124004
rect 89558 123964 89600 124004
rect 89272 123955 89640 123964
rect 104392 124004 104760 124013
rect 104432 123964 104474 124004
rect 104514 123964 104556 124004
rect 104596 123964 104638 124004
rect 104678 123964 104720 124004
rect 104392 123955 104760 123964
rect 119512 124004 119880 124013
rect 119552 123964 119594 124004
rect 119634 123964 119676 124004
rect 119716 123964 119758 124004
rect 119798 123964 119840 124004
rect 119512 123955 119880 123964
rect 134632 124004 135000 124013
rect 134672 123964 134714 124004
rect 134754 123964 134796 124004
rect 134836 123964 134878 124004
rect 134918 123964 134960 124004
rect 134632 123955 135000 123964
rect 149752 124004 150120 124013
rect 149792 123964 149834 124004
rect 149874 123964 149916 124004
rect 149956 123964 149998 124004
rect 150038 123964 150080 124004
rect 149752 123955 150120 123964
rect 75392 123248 75760 123257
rect 75432 123208 75474 123248
rect 75514 123208 75556 123248
rect 75596 123208 75638 123248
rect 75678 123208 75720 123248
rect 75392 123199 75760 123208
rect 90512 123248 90880 123257
rect 90552 123208 90594 123248
rect 90634 123208 90676 123248
rect 90716 123208 90758 123248
rect 90798 123208 90840 123248
rect 90512 123199 90880 123208
rect 105632 123248 106000 123257
rect 105672 123208 105714 123248
rect 105754 123208 105796 123248
rect 105836 123208 105878 123248
rect 105918 123208 105960 123248
rect 105632 123199 106000 123208
rect 120752 123248 121120 123257
rect 120792 123208 120834 123248
rect 120874 123208 120916 123248
rect 120956 123208 120998 123248
rect 121038 123208 121080 123248
rect 120752 123199 121120 123208
rect 135872 123248 136240 123257
rect 135912 123208 135954 123248
rect 135994 123208 136036 123248
rect 136076 123208 136118 123248
rect 136158 123208 136200 123248
rect 135872 123199 136240 123208
rect 150992 123248 151360 123257
rect 151032 123208 151074 123248
rect 151114 123208 151156 123248
rect 151196 123208 151238 123248
rect 151278 123208 151320 123248
rect 150992 123199 151360 123208
rect 74152 122492 74520 122501
rect 74192 122452 74234 122492
rect 74274 122452 74316 122492
rect 74356 122452 74398 122492
rect 74438 122452 74480 122492
rect 74152 122443 74520 122452
rect 89272 122492 89640 122501
rect 89312 122452 89354 122492
rect 89394 122452 89436 122492
rect 89476 122452 89518 122492
rect 89558 122452 89600 122492
rect 89272 122443 89640 122452
rect 104392 122492 104760 122501
rect 104432 122452 104474 122492
rect 104514 122452 104556 122492
rect 104596 122452 104638 122492
rect 104678 122452 104720 122492
rect 104392 122443 104760 122452
rect 119512 122492 119880 122501
rect 119552 122452 119594 122492
rect 119634 122452 119676 122492
rect 119716 122452 119758 122492
rect 119798 122452 119840 122492
rect 119512 122443 119880 122452
rect 134632 122492 135000 122501
rect 134672 122452 134714 122492
rect 134754 122452 134796 122492
rect 134836 122452 134878 122492
rect 134918 122452 134960 122492
rect 134632 122443 135000 122452
rect 149752 122492 150120 122501
rect 149792 122452 149834 122492
rect 149874 122452 149916 122492
rect 149956 122452 149998 122492
rect 150038 122452 150080 122492
rect 149752 122443 150120 122452
rect 75392 121736 75760 121745
rect 75432 121696 75474 121736
rect 75514 121696 75556 121736
rect 75596 121696 75638 121736
rect 75678 121696 75720 121736
rect 75392 121687 75760 121696
rect 90512 121736 90880 121745
rect 90552 121696 90594 121736
rect 90634 121696 90676 121736
rect 90716 121696 90758 121736
rect 90798 121696 90840 121736
rect 90512 121687 90880 121696
rect 105632 121736 106000 121745
rect 105672 121696 105714 121736
rect 105754 121696 105796 121736
rect 105836 121696 105878 121736
rect 105918 121696 105960 121736
rect 105632 121687 106000 121696
rect 120752 121736 121120 121745
rect 120792 121696 120834 121736
rect 120874 121696 120916 121736
rect 120956 121696 120998 121736
rect 121038 121696 121080 121736
rect 120752 121687 121120 121696
rect 135872 121736 136240 121745
rect 135912 121696 135954 121736
rect 135994 121696 136036 121736
rect 136076 121696 136118 121736
rect 136158 121696 136200 121736
rect 135872 121687 136240 121696
rect 150992 121736 151360 121745
rect 151032 121696 151074 121736
rect 151114 121696 151156 121736
rect 151196 121696 151238 121736
rect 151278 121696 151320 121736
rect 150992 121687 151360 121696
rect 74152 120980 74520 120989
rect 74192 120940 74234 120980
rect 74274 120940 74316 120980
rect 74356 120940 74398 120980
rect 74438 120940 74480 120980
rect 74152 120931 74520 120940
rect 89272 120980 89640 120989
rect 89312 120940 89354 120980
rect 89394 120940 89436 120980
rect 89476 120940 89518 120980
rect 89558 120940 89600 120980
rect 89272 120931 89640 120940
rect 104392 120980 104760 120989
rect 104432 120940 104474 120980
rect 104514 120940 104556 120980
rect 104596 120940 104638 120980
rect 104678 120940 104720 120980
rect 104392 120931 104760 120940
rect 119512 120980 119880 120989
rect 119552 120940 119594 120980
rect 119634 120940 119676 120980
rect 119716 120940 119758 120980
rect 119798 120940 119840 120980
rect 119512 120931 119880 120940
rect 134632 120980 135000 120989
rect 134672 120940 134714 120980
rect 134754 120940 134796 120980
rect 134836 120940 134878 120980
rect 134918 120940 134960 120980
rect 134632 120931 135000 120940
rect 149752 120980 150120 120989
rect 149792 120940 149834 120980
rect 149874 120940 149916 120980
rect 149956 120940 149998 120980
rect 150038 120940 150080 120980
rect 149752 120931 150120 120940
rect 75392 120224 75760 120233
rect 75432 120184 75474 120224
rect 75514 120184 75556 120224
rect 75596 120184 75638 120224
rect 75678 120184 75720 120224
rect 75392 120175 75760 120184
rect 90512 120224 90880 120233
rect 90552 120184 90594 120224
rect 90634 120184 90676 120224
rect 90716 120184 90758 120224
rect 90798 120184 90840 120224
rect 90512 120175 90880 120184
rect 105632 120224 106000 120233
rect 105672 120184 105714 120224
rect 105754 120184 105796 120224
rect 105836 120184 105878 120224
rect 105918 120184 105960 120224
rect 105632 120175 106000 120184
rect 120752 120224 121120 120233
rect 120792 120184 120834 120224
rect 120874 120184 120916 120224
rect 120956 120184 120998 120224
rect 121038 120184 121080 120224
rect 120752 120175 121120 120184
rect 135872 120224 136240 120233
rect 135912 120184 135954 120224
rect 135994 120184 136036 120224
rect 136076 120184 136118 120224
rect 136158 120184 136200 120224
rect 135872 120175 136240 120184
rect 150992 120224 151360 120233
rect 151032 120184 151074 120224
rect 151114 120184 151156 120224
rect 151196 120184 151238 120224
rect 151278 120184 151320 120224
rect 150992 120175 151360 120184
rect 74152 119468 74520 119477
rect 74192 119428 74234 119468
rect 74274 119428 74316 119468
rect 74356 119428 74398 119468
rect 74438 119428 74480 119468
rect 74152 119419 74520 119428
rect 89272 119468 89640 119477
rect 89312 119428 89354 119468
rect 89394 119428 89436 119468
rect 89476 119428 89518 119468
rect 89558 119428 89600 119468
rect 89272 119419 89640 119428
rect 104392 119468 104760 119477
rect 104432 119428 104474 119468
rect 104514 119428 104556 119468
rect 104596 119428 104638 119468
rect 104678 119428 104720 119468
rect 104392 119419 104760 119428
rect 119512 119468 119880 119477
rect 119552 119428 119594 119468
rect 119634 119428 119676 119468
rect 119716 119428 119758 119468
rect 119798 119428 119840 119468
rect 119512 119419 119880 119428
rect 134632 119468 135000 119477
rect 134672 119428 134714 119468
rect 134754 119428 134796 119468
rect 134836 119428 134878 119468
rect 134918 119428 134960 119468
rect 134632 119419 135000 119428
rect 149752 119468 150120 119477
rect 149792 119428 149834 119468
rect 149874 119428 149916 119468
rect 149956 119428 149998 119468
rect 150038 119428 150080 119468
rect 149752 119419 150120 119428
rect 75392 118712 75760 118721
rect 75432 118672 75474 118712
rect 75514 118672 75556 118712
rect 75596 118672 75638 118712
rect 75678 118672 75720 118712
rect 75392 118663 75760 118672
rect 90512 118712 90880 118721
rect 90552 118672 90594 118712
rect 90634 118672 90676 118712
rect 90716 118672 90758 118712
rect 90798 118672 90840 118712
rect 90512 118663 90880 118672
rect 105632 118712 106000 118721
rect 105672 118672 105714 118712
rect 105754 118672 105796 118712
rect 105836 118672 105878 118712
rect 105918 118672 105960 118712
rect 105632 118663 106000 118672
rect 120752 118712 121120 118721
rect 120792 118672 120834 118712
rect 120874 118672 120916 118712
rect 120956 118672 120998 118712
rect 121038 118672 121080 118712
rect 120752 118663 121120 118672
rect 135872 118712 136240 118721
rect 135912 118672 135954 118712
rect 135994 118672 136036 118712
rect 136076 118672 136118 118712
rect 136158 118672 136200 118712
rect 135872 118663 136240 118672
rect 150992 118712 151360 118721
rect 151032 118672 151074 118712
rect 151114 118672 151156 118712
rect 151196 118672 151238 118712
rect 151278 118672 151320 118712
rect 150992 118663 151360 118672
rect 74152 117956 74520 117965
rect 74192 117916 74234 117956
rect 74274 117916 74316 117956
rect 74356 117916 74398 117956
rect 74438 117916 74480 117956
rect 74152 117907 74520 117916
rect 89272 117956 89640 117965
rect 89312 117916 89354 117956
rect 89394 117916 89436 117956
rect 89476 117916 89518 117956
rect 89558 117916 89600 117956
rect 89272 117907 89640 117916
rect 104392 117956 104760 117965
rect 104432 117916 104474 117956
rect 104514 117916 104556 117956
rect 104596 117916 104638 117956
rect 104678 117916 104720 117956
rect 104392 117907 104760 117916
rect 119512 117956 119880 117965
rect 119552 117916 119594 117956
rect 119634 117916 119676 117956
rect 119716 117916 119758 117956
rect 119798 117916 119840 117956
rect 119512 117907 119880 117916
rect 134632 117956 135000 117965
rect 134672 117916 134714 117956
rect 134754 117916 134796 117956
rect 134836 117916 134878 117956
rect 134918 117916 134960 117956
rect 134632 117907 135000 117916
rect 149752 117956 150120 117965
rect 149792 117916 149834 117956
rect 149874 117916 149916 117956
rect 149956 117916 149998 117956
rect 150038 117916 150080 117956
rect 149752 117907 150120 117916
rect 75392 117200 75760 117209
rect 75432 117160 75474 117200
rect 75514 117160 75556 117200
rect 75596 117160 75638 117200
rect 75678 117160 75720 117200
rect 75392 117151 75760 117160
rect 90512 117200 90880 117209
rect 90552 117160 90594 117200
rect 90634 117160 90676 117200
rect 90716 117160 90758 117200
rect 90798 117160 90840 117200
rect 90512 117151 90880 117160
rect 105632 117200 106000 117209
rect 105672 117160 105714 117200
rect 105754 117160 105796 117200
rect 105836 117160 105878 117200
rect 105918 117160 105960 117200
rect 105632 117151 106000 117160
rect 120752 117200 121120 117209
rect 120792 117160 120834 117200
rect 120874 117160 120916 117200
rect 120956 117160 120998 117200
rect 121038 117160 121080 117200
rect 120752 117151 121120 117160
rect 135872 117200 136240 117209
rect 135912 117160 135954 117200
rect 135994 117160 136036 117200
rect 136076 117160 136118 117200
rect 136158 117160 136200 117200
rect 135872 117151 136240 117160
rect 150992 117200 151360 117209
rect 151032 117160 151074 117200
rect 151114 117160 151156 117200
rect 151196 117160 151238 117200
rect 151278 117160 151320 117200
rect 150992 117151 151360 117160
rect 74152 116444 74520 116453
rect 74192 116404 74234 116444
rect 74274 116404 74316 116444
rect 74356 116404 74398 116444
rect 74438 116404 74480 116444
rect 74152 116395 74520 116404
rect 89272 116444 89640 116453
rect 89312 116404 89354 116444
rect 89394 116404 89436 116444
rect 89476 116404 89518 116444
rect 89558 116404 89600 116444
rect 89272 116395 89640 116404
rect 104392 116444 104760 116453
rect 104432 116404 104474 116444
rect 104514 116404 104556 116444
rect 104596 116404 104638 116444
rect 104678 116404 104720 116444
rect 104392 116395 104760 116404
rect 119512 116444 119880 116453
rect 119552 116404 119594 116444
rect 119634 116404 119676 116444
rect 119716 116404 119758 116444
rect 119798 116404 119840 116444
rect 119512 116395 119880 116404
rect 134632 116444 135000 116453
rect 134672 116404 134714 116444
rect 134754 116404 134796 116444
rect 134836 116404 134878 116444
rect 134918 116404 134960 116444
rect 134632 116395 135000 116404
rect 149752 116444 150120 116453
rect 149792 116404 149834 116444
rect 149874 116404 149916 116444
rect 149956 116404 149998 116444
rect 150038 116404 150080 116444
rect 149752 116395 150120 116404
rect 75392 115688 75760 115697
rect 75432 115648 75474 115688
rect 75514 115648 75556 115688
rect 75596 115648 75638 115688
rect 75678 115648 75720 115688
rect 75392 115639 75760 115648
rect 90512 115688 90880 115697
rect 90552 115648 90594 115688
rect 90634 115648 90676 115688
rect 90716 115648 90758 115688
rect 90798 115648 90840 115688
rect 90512 115639 90880 115648
rect 105632 115688 106000 115697
rect 105672 115648 105714 115688
rect 105754 115648 105796 115688
rect 105836 115648 105878 115688
rect 105918 115648 105960 115688
rect 105632 115639 106000 115648
rect 120752 115688 121120 115697
rect 120792 115648 120834 115688
rect 120874 115648 120916 115688
rect 120956 115648 120998 115688
rect 121038 115648 121080 115688
rect 120752 115639 121120 115648
rect 135872 115688 136240 115697
rect 135912 115648 135954 115688
rect 135994 115648 136036 115688
rect 136076 115648 136118 115688
rect 136158 115648 136200 115688
rect 135872 115639 136240 115648
rect 150992 115688 151360 115697
rect 151032 115648 151074 115688
rect 151114 115648 151156 115688
rect 151196 115648 151238 115688
rect 151278 115648 151320 115688
rect 150992 115639 151360 115648
rect 74152 114932 74520 114941
rect 74192 114892 74234 114932
rect 74274 114892 74316 114932
rect 74356 114892 74398 114932
rect 74438 114892 74480 114932
rect 74152 114883 74520 114892
rect 89272 114932 89640 114941
rect 89312 114892 89354 114932
rect 89394 114892 89436 114932
rect 89476 114892 89518 114932
rect 89558 114892 89600 114932
rect 89272 114883 89640 114892
rect 104392 114932 104760 114941
rect 104432 114892 104474 114932
rect 104514 114892 104556 114932
rect 104596 114892 104638 114932
rect 104678 114892 104720 114932
rect 104392 114883 104760 114892
rect 119512 114932 119880 114941
rect 119552 114892 119594 114932
rect 119634 114892 119676 114932
rect 119716 114892 119758 114932
rect 119798 114892 119840 114932
rect 119512 114883 119880 114892
rect 134632 114932 135000 114941
rect 134672 114892 134714 114932
rect 134754 114892 134796 114932
rect 134836 114892 134878 114932
rect 134918 114892 134960 114932
rect 134632 114883 135000 114892
rect 149752 114932 150120 114941
rect 149792 114892 149834 114932
rect 149874 114892 149916 114932
rect 149956 114892 149998 114932
rect 150038 114892 150080 114932
rect 149752 114883 150120 114892
rect 75392 114176 75760 114185
rect 75432 114136 75474 114176
rect 75514 114136 75556 114176
rect 75596 114136 75638 114176
rect 75678 114136 75720 114176
rect 75392 114127 75760 114136
rect 90512 114176 90880 114185
rect 90552 114136 90594 114176
rect 90634 114136 90676 114176
rect 90716 114136 90758 114176
rect 90798 114136 90840 114176
rect 90512 114127 90880 114136
rect 105632 114176 106000 114185
rect 105672 114136 105714 114176
rect 105754 114136 105796 114176
rect 105836 114136 105878 114176
rect 105918 114136 105960 114176
rect 105632 114127 106000 114136
rect 120752 114176 121120 114185
rect 120792 114136 120834 114176
rect 120874 114136 120916 114176
rect 120956 114136 120998 114176
rect 121038 114136 121080 114176
rect 120752 114127 121120 114136
rect 135872 114176 136240 114185
rect 135912 114136 135954 114176
rect 135994 114136 136036 114176
rect 136076 114136 136118 114176
rect 136158 114136 136200 114176
rect 135872 114127 136240 114136
rect 150992 114176 151360 114185
rect 151032 114136 151074 114176
rect 151114 114136 151156 114176
rect 151196 114136 151238 114176
rect 151278 114136 151320 114176
rect 150992 114127 151360 114136
rect 74152 113420 74520 113429
rect 74192 113380 74234 113420
rect 74274 113380 74316 113420
rect 74356 113380 74398 113420
rect 74438 113380 74480 113420
rect 74152 113371 74520 113380
rect 89272 113420 89640 113429
rect 89312 113380 89354 113420
rect 89394 113380 89436 113420
rect 89476 113380 89518 113420
rect 89558 113380 89600 113420
rect 89272 113371 89640 113380
rect 104392 113420 104760 113429
rect 104432 113380 104474 113420
rect 104514 113380 104556 113420
rect 104596 113380 104638 113420
rect 104678 113380 104720 113420
rect 104392 113371 104760 113380
rect 119512 113420 119880 113429
rect 119552 113380 119594 113420
rect 119634 113380 119676 113420
rect 119716 113380 119758 113420
rect 119798 113380 119840 113420
rect 119512 113371 119880 113380
rect 134632 113420 135000 113429
rect 134672 113380 134714 113420
rect 134754 113380 134796 113420
rect 134836 113380 134878 113420
rect 134918 113380 134960 113420
rect 134632 113371 135000 113380
rect 149752 113420 150120 113429
rect 149792 113380 149834 113420
rect 149874 113380 149916 113420
rect 149956 113380 149998 113420
rect 150038 113380 150080 113420
rect 149752 113371 150120 113380
rect 75392 112664 75760 112673
rect 75432 112624 75474 112664
rect 75514 112624 75556 112664
rect 75596 112624 75638 112664
rect 75678 112624 75720 112664
rect 75392 112615 75760 112624
rect 90512 112664 90880 112673
rect 90552 112624 90594 112664
rect 90634 112624 90676 112664
rect 90716 112624 90758 112664
rect 90798 112624 90840 112664
rect 90512 112615 90880 112624
rect 105632 112664 106000 112673
rect 105672 112624 105714 112664
rect 105754 112624 105796 112664
rect 105836 112624 105878 112664
rect 105918 112624 105960 112664
rect 105632 112615 106000 112624
rect 120752 112664 121120 112673
rect 120792 112624 120834 112664
rect 120874 112624 120916 112664
rect 120956 112624 120998 112664
rect 121038 112624 121080 112664
rect 120752 112615 121120 112624
rect 135872 112664 136240 112673
rect 135912 112624 135954 112664
rect 135994 112624 136036 112664
rect 136076 112624 136118 112664
rect 136158 112624 136200 112664
rect 135872 112615 136240 112624
rect 150992 112664 151360 112673
rect 151032 112624 151074 112664
rect 151114 112624 151156 112664
rect 151196 112624 151238 112664
rect 151278 112624 151320 112664
rect 150992 112615 151360 112624
rect 74152 111908 74520 111917
rect 74192 111868 74234 111908
rect 74274 111868 74316 111908
rect 74356 111868 74398 111908
rect 74438 111868 74480 111908
rect 74152 111859 74520 111868
rect 89272 111908 89640 111917
rect 89312 111868 89354 111908
rect 89394 111868 89436 111908
rect 89476 111868 89518 111908
rect 89558 111868 89600 111908
rect 89272 111859 89640 111868
rect 104392 111908 104760 111917
rect 104432 111868 104474 111908
rect 104514 111868 104556 111908
rect 104596 111868 104638 111908
rect 104678 111868 104720 111908
rect 104392 111859 104760 111868
rect 119512 111908 119880 111917
rect 119552 111868 119594 111908
rect 119634 111868 119676 111908
rect 119716 111868 119758 111908
rect 119798 111868 119840 111908
rect 119512 111859 119880 111868
rect 134632 111908 135000 111917
rect 134672 111868 134714 111908
rect 134754 111868 134796 111908
rect 134836 111868 134878 111908
rect 134918 111868 134960 111908
rect 134632 111859 135000 111868
rect 149752 111908 150120 111917
rect 149792 111868 149834 111908
rect 149874 111868 149916 111908
rect 149956 111868 149998 111908
rect 150038 111868 150080 111908
rect 149752 111859 150120 111868
rect 75392 111152 75760 111161
rect 75432 111112 75474 111152
rect 75514 111112 75556 111152
rect 75596 111112 75638 111152
rect 75678 111112 75720 111152
rect 75392 111103 75760 111112
rect 90512 111152 90880 111161
rect 90552 111112 90594 111152
rect 90634 111112 90676 111152
rect 90716 111112 90758 111152
rect 90798 111112 90840 111152
rect 90512 111103 90880 111112
rect 105632 111152 106000 111161
rect 105672 111112 105714 111152
rect 105754 111112 105796 111152
rect 105836 111112 105878 111152
rect 105918 111112 105960 111152
rect 105632 111103 106000 111112
rect 120752 111152 121120 111161
rect 120792 111112 120834 111152
rect 120874 111112 120916 111152
rect 120956 111112 120998 111152
rect 121038 111112 121080 111152
rect 120752 111103 121120 111112
rect 135872 111152 136240 111161
rect 135912 111112 135954 111152
rect 135994 111112 136036 111152
rect 136076 111112 136118 111152
rect 136158 111112 136200 111152
rect 135872 111103 136240 111112
rect 150992 111152 151360 111161
rect 151032 111112 151074 111152
rect 151114 111112 151156 111152
rect 151196 111112 151238 111152
rect 151278 111112 151320 111152
rect 150992 111103 151360 111112
rect 74152 110396 74520 110405
rect 74192 110356 74234 110396
rect 74274 110356 74316 110396
rect 74356 110356 74398 110396
rect 74438 110356 74480 110396
rect 74152 110347 74520 110356
rect 89272 110396 89640 110405
rect 89312 110356 89354 110396
rect 89394 110356 89436 110396
rect 89476 110356 89518 110396
rect 89558 110356 89600 110396
rect 89272 110347 89640 110356
rect 104392 110396 104760 110405
rect 104432 110356 104474 110396
rect 104514 110356 104556 110396
rect 104596 110356 104638 110396
rect 104678 110356 104720 110396
rect 104392 110347 104760 110356
rect 119512 110396 119880 110405
rect 119552 110356 119594 110396
rect 119634 110356 119676 110396
rect 119716 110356 119758 110396
rect 119798 110356 119840 110396
rect 119512 110347 119880 110356
rect 134632 110396 135000 110405
rect 134672 110356 134714 110396
rect 134754 110356 134796 110396
rect 134836 110356 134878 110396
rect 134918 110356 134960 110396
rect 134632 110347 135000 110356
rect 149752 110396 150120 110405
rect 149792 110356 149834 110396
rect 149874 110356 149916 110396
rect 149956 110356 149998 110396
rect 150038 110356 150080 110396
rect 149752 110347 150120 110356
rect 75392 109640 75760 109649
rect 75432 109600 75474 109640
rect 75514 109600 75556 109640
rect 75596 109600 75638 109640
rect 75678 109600 75720 109640
rect 75392 109591 75760 109600
rect 90512 109640 90880 109649
rect 90552 109600 90594 109640
rect 90634 109600 90676 109640
rect 90716 109600 90758 109640
rect 90798 109600 90840 109640
rect 90512 109591 90880 109600
rect 105632 109640 106000 109649
rect 105672 109600 105714 109640
rect 105754 109600 105796 109640
rect 105836 109600 105878 109640
rect 105918 109600 105960 109640
rect 105632 109591 106000 109600
rect 120752 109640 121120 109649
rect 120792 109600 120834 109640
rect 120874 109600 120916 109640
rect 120956 109600 120998 109640
rect 121038 109600 121080 109640
rect 120752 109591 121120 109600
rect 135872 109640 136240 109649
rect 135912 109600 135954 109640
rect 135994 109600 136036 109640
rect 136076 109600 136118 109640
rect 136158 109600 136200 109640
rect 135872 109591 136240 109600
rect 150992 109640 151360 109649
rect 151032 109600 151074 109640
rect 151114 109600 151156 109640
rect 151196 109600 151238 109640
rect 151278 109600 151320 109640
rect 150992 109591 151360 109600
rect 74152 108884 74520 108893
rect 74192 108844 74234 108884
rect 74274 108844 74316 108884
rect 74356 108844 74398 108884
rect 74438 108844 74480 108884
rect 74152 108835 74520 108844
rect 89272 108884 89640 108893
rect 89312 108844 89354 108884
rect 89394 108844 89436 108884
rect 89476 108844 89518 108884
rect 89558 108844 89600 108884
rect 89272 108835 89640 108844
rect 104392 108884 104760 108893
rect 104432 108844 104474 108884
rect 104514 108844 104556 108884
rect 104596 108844 104638 108884
rect 104678 108844 104720 108884
rect 104392 108835 104760 108844
rect 119512 108884 119880 108893
rect 119552 108844 119594 108884
rect 119634 108844 119676 108884
rect 119716 108844 119758 108884
rect 119798 108844 119840 108884
rect 119512 108835 119880 108844
rect 134632 108884 135000 108893
rect 134672 108844 134714 108884
rect 134754 108844 134796 108884
rect 134836 108844 134878 108884
rect 134918 108844 134960 108884
rect 134632 108835 135000 108844
rect 149752 108884 150120 108893
rect 149792 108844 149834 108884
rect 149874 108844 149916 108884
rect 149956 108844 149998 108884
rect 150038 108844 150080 108884
rect 149752 108835 150120 108844
rect 75392 108128 75760 108137
rect 75432 108088 75474 108128
rect 75514 108088 75556 108128
rect 75596 108088 75638 108128
rect 75678 108088 75720 108128
rect 75392 108079 75760 108088
rect 90512 108128 90880 108137
rect 90552 108088 90594 108128
rect 90634 108088 90676 108128
rect 90716 108088 90758 108128
rect 90798 108088 90840 108128
rect 90512 108079 90880 108088
rect 105632 108128 106000 108137
rect 105672 108088 105714 108128
rect 105754 108088 105796 108128
rect 105836 108088 105878 108128
rect 105918 108088 105960 108128
rect 105632 108079 106000 108088
rect 120752 108128 121120 108137
rect 120792 108088 120834 108128
rect 120874 108088 120916 108128
rect 120956 108088 120998 108128
rect 121038 108088 121080 108128
rect 120752 108079 121120 108088
rect 135872 108128 136240 108137
rect 135912 108088 135954 108128
rect 135994 108088 136036 108128
rect 136076 108088 136118 108128
rect 136158 108088 136200 108128
rect 135872 108079 136240 108088
rect 150992 108128 151360 108137
rect 151032 108088 151074 108128
rect 151114 108088 151156 108128
rect 151196 108088 151238 108128
rect 151278 108088 151320 108128
rect 150992 108079 151360 108088
rect 74152 107372 74520 107381
rect 74192 107332 74234 107372
rect 74274 107332 74316 107372
rect 74356 107332 74398 107372
rect 74438 107332 74480 107372
rect 74152 107323 74520 107332
rect 89272 107372 89640 107381
rect 89312 107332 89354 107372
rect 89394 107332 89436 107372
rect 89476 107332 89518 107372
rect 89558 107332 89600 107372
rect 89272 107323 89640 107332
rect 104392 107372 104760 107381
rect 104432 107332 104474 107372
rect 104514 107332 104556 107372
rect 104596 107332 104638 107372
rect 104678 107332 104720 107372
rect 104392 107323 104760 107332
rect 119512 107372 119880 107381
rect 119552 107332 119594 107372
rect 119634 107332 119676 107372
rect 119716 107332 119758 107372
rect 119798 107332 119840 107372
rect 119512 107323 119880 107332
rect 134632 107372 135000 107381
rect 134672 107332 134714 107372
rect 134754 107332 134796 107372
rect 134836 107332 134878 107372
rect 134918 107332 134960 107372
rect 134632 107323 135000 107332
rect 149752 107372 150120 107381
rect 149792 107332 149834 107372
rect 149874 107332 149916 107372
rect 149956 107332 149998 107372
rect 150038 107332 150080 107372
rect 149752 107323 150120 107332
rect 75392 106616 75760 106625
rect 75432 106576 75474 106616
rect 75514 106576 75556 106616
rect 75596 106576 75638 106616
rect 75678 106576 75720 106616
rect 75392 106567 75760 106576
rect 90512 106616 90880 106625
rect 90552 106576 90594 106616
rect 90634 106576 90676 106616
rect 90716 106576 90758 106616
rect 90798 106576 90840 106616
rect 90512 106567 90880 106576
rect 105632 106616 106000 106625
rect 105672 106576 105714 106616
rect 105754 106576 105796 106616
rect 105836 106576 105878 106616
rect 105918 106576 105960 106616
rect 105632 106567 106000 106576
rect 120752 106616 121120 106625
rect 120792 106576 120834 106616
rect 120874 106576 120916 106616
rect 120956 106576 120998 106616
rect 121038 106576 121080 106616
rect 120752 106567 121120 106576
rect 135872 106616 136240 106625
rect 135912 106576 135954 106616
rect 135994 106576 136036 106616
rect 136076 106576 136118 106616
rect 136158 106576 136200 106616
rect 135872 106567 136240 106576
rect 150992 106616 151360 106625
rect 151032 106576 151074 106616
rect 151114 106576 151156 106616
rect 151196 106576 151238 106616
rect 151278 106576 151320 106616
rect 150992 106567 151360 106576
rect 74152 105860 74520 105869
rect 74192 105820 74234 105860
rect 74274 105820 74316 105860
rect 74356 105820 74398 105860
rect 74438 105820 74480 105860
rect 74152 105811 74520 105820
rect 89272 105860 89640 105869
rect 89312 105820 89354 105860
rect 89394 105820 89436 105860
rect 89476 105820 89518 105860
rect 89558 105820 89600 105860
rect 89272 105811 89640 105820
rect 104392 105860 104760 105869
rect 104432 105820 104474 105860
rect 104514 105820 104556 105860
rect 104596 105820 104638 105860
rect 104678 105820 104720 105860
rect 104392 105811 104760 105820
rect 119512 105860 119880 105869
rect 119552 105820 119594 105860
rect 119634 105820 119676 105860
rect 119716 105820 119758 105860
rect 119798 105820 119840 105860
rect 119512 105811 119880 105820
rect 134632 105860 135000 105869
rect 134672 105820 134714 105860
rect 134754 105820 134796 105860
rect 134836 105820 134878 105860
rect 134918 105820 134960 105860
rect 134632 105811 135000 105820
rect 149752 105860 150120 105869
rect 149792 105820 149834 105860
rect 149874 105820 149916 105860
rect 149956 105820 149998 105860
rect 150038 105820 150080 105860
rect 149752 105811 150120 105820
rect 75392 105104 75760 105113
rect 75432 105064 75474 105104
rect 75514 105064 75556 105104
rect 75596 105064 75638 105104
rect 75678 105064 75720 105104
rect 75392 105055 75760 105064
rect 90512 105104 90880 105113
rect 90552 105064 90594 105104
rect 90634 105064 90676 105104
rect 90716 105064 90758 105104
rect 90798 105064 90840 105104
rect 90512 105055 90880 105064
rect 105632 105104 106000 105113
rect 105672 105064 105714 105104
rect 105754 105064 105796 105104
rect 105836 105064 105878 105104
rect 105918 105064 105960 105104
rect 105632 105055 106000 105064
rect 120752 105104 121120 105113
rect 120792 105064 120834 105104
rect 120874 105064 120916 105104
rect 120956 105064 120998 105104
rect 121038 105064 121080 105104
rect 120752 105055 121120 105064
rect 135872 105104 136240 105113
rect 135912 105064 135954 105104
rect 135994 105064 136036 105104
rect 136076 105064 136118 105104
rect 136158 105064 136200 105104
rect 135872 105055 136240 105064
rect 150992 105104 151360 105113
rect 151032 105064 151074 105104
rect 151114 105064 151156 105104
rect 151196 105064 151238 105104
rect 151278 105064 151320 105104
rect 150992 105055 151360 105064
rect 74152 104348 74520 104357
rect 74192 104308 74234 104348
rect 74274 104308 74316 104348
rect 74356 104308 74398 104348
rect 74438 104308 74480 104348
rect 74152 104299 74520 104308
rect 89272 104348 89640 104357
rect 89312 104308 89354 104348
rect 89394 104308 89436 104348
rect 89476 104308 89518 104348
rect 89558 104308 89600 104348
rect 89272 104299 89640 104308
rect 104392 104348 104760 104357
rect 104432 104308 104474 104348
rect 104514 104308 104556 104348
rect 104596 104308 104638 104348
rect 104678 104308 104720 104348
rect 104392 104299 104760 104308
rect 119512 104348 119880 104357
rect 119552 104308 119594 104348
rect 119634 104308 119676 104348
rect 119716 104308 119758 104348
rect 119798 104308 119840 104348
rect 119512 104299 119880 104308
rect 134632 104348 135000 104357
rect 134672 104308 134714 104348
rect 134754 104308 134796 104348
rect 134836 104308 134878 104348
rect 134918 104308 134960 104348
rect 134632 104299 135000 104308
rect 149752 104348 150120 104357
rect 149792 104308 149834 104348
rect 149874 104308 149916 104348
rect 149956 104308 149998 104348
rect 150038 104308 150080 104348
rect 149752 104299 150120 104308
rect 75392 103592 75760 103601
rect 75432 103552 75474 103592
rect 75514 103552 75556 103592
rect 75596 103552 75638 103592
rect 75678 103552 75720 103592
rect 75392 103543 75760 103552
rect 90512 103592 90880 103601
rect 90552 103552 90594 103592
rect 90634 103552 90676 103592
rect 90716 103552 90758 103592
rect 90798 103552 90840 103592
rect 90512 103543 90880 103552
rect 105632 103592 106000 103601
rect 105672 103552 105714 103592
rect 105754 103552 105796 103592
rect 105836 103552 105878 103592
rect 105918 103552 105960 103592
rect 105632 103543 106000 103552
rect 120752 103592 121120 103601
rect 120792 103552 120834 103592
rect 120874 103552 120916 103592
rect 120956 103552 120998 103592
rect 121038 103552 121080 103592
rect 120752 103543 121120 103552
rect 135872 103592 136240 103601
rect 135912 103552 135954 103592
rect 135994 103552 136036 103592
rect 136076 103552 136118 103592
rect 136158 103552 136200 103592
rect 135872 103543 136240 103552
rect 150992 103592 151360 103601
rect 151032 103552 151074 103592
rect 151114 103552 151156 103592
rect 151196 103552 151238 103592
rect 151278 103552 151320 103592
rect 150992 103543 151360 103552
rect 74152 102836 74520 102845
rect 74192 102796 74234 102836
rect 74274 102796 74316 102836
rect 74356 102796 74398 102836
rect 74438 102796 74480 102836
rect 74152 102787 74520 102796
rect 89272 102836 89640 102845
rect 89312 102796 89354 102836
rect 89394 102796 89436 102836
rect 89476 102796 89518 102836
rect 89558 102796 89600 102836
rect 89272 102787 89640 102796
rect 104392 102836 104760 102845
rect 104432 102796 104474 102836
rect 104514 102796 104556 102836
rect 104596 102796 104638 102836
rect 104678 102796 104720 102836
rect 104392 102787 104760 102796
rect 119512 102836 119880 102845
rect 119552 102796 119594 102836
rect 119634 102796 119676 102836
rect 119716 102796 119758 102836
rect 119798 102796 119840 102836
rect 119512 102787 119880 102796
rect 134632 102836 135000 102845
rect 134672 102796 134714 102836
rect 134754 102796 134796 102836
rect 134836 102796 134878 102836
rect 134918 102796 134960 102836
rect 134632 102787 135000 102796
rect 149752 102836 150120 102845
rect 149792 102796 149834 102836
rect 149874 102796 149916 102836
rect 149956 102796 149998 102836
rect 150038 102796 150080 102836
rect 149752 102787 150120 102796
rect 75392 102080 75760 102089
rect 75432 102040 75474 102080
rect 75514 102040 75556 102080
rect 75596 102040 75638 102080
rect 75678 102040 75720 102080
rect 75392 102031 75760 102040
rect 90512 102080 90880 102089
rect 90552 102040 90594 102080
rect 90634 102040 90676 102080
rect 90716 102040 90758 102080
rect 90798 102040 90840 102080
rect 90512 102031 90880 102040
rect 105632 102080 106000 102089
rect 105672 102040 105714 102080
rect 105754 102040 105796 102080
rect 105836 102040 105878 102080
rect 105918 102040 105960 102080
rect 105632 102031 106000 102040
rect 120752 102080 121120 102089
rect 120792 102040 120834 102080
rect 120874 102040 120916 102080
rect 120956 102040 120998 102080
rect 121038 102040 121080 102080
rect 120752 102031 121120 102040
rect 135872 102080 136240 102089
rect 135912 102040 135954 102080
rect 135994 102040 136036 102080
rect 136076 102040 136118 102080
rect 136158 102040 136200 102080
rect 135872 102031 136240 102040
rect 150992 102080 151360 102089
rect 151032 102040 151074 102080
rect 151114 102040 151156 102080
rect 151196 102040 151238 102080
rect 151278 102040 151320 102080
rect 150992 102031 151360 102040
rect 74152 101324 74520 101333
rect 74192 101284 74234 101324
rect 74274 101284 74316 101324
rect 74356 101284 74398 101324
rect 74438 101284 74480 101324
rect 74152 101275 74520 101284
rect 89272 101324 89640 101333
rect 89312 101284 89354 101324
rect 89394 101284 89436 101324
rect 89476 101284 89518 101324
rect 89558 101284 89600 101324
rect 89272 101275 89640 101284
rect 104392 101324 104760 101333
rect 104432 101284 104474 101324
rect 104514 101284 104556 101324
rect 104596 101284 104638 101324
rect 104678 101284 104720 101324
rect 104392 101275 104760 101284
rect 119512 101324 119880 101333
rect 119552 101284 119594 101324
rect 119634 101284 119676 101324
rect 119716 101284 119758 101324
rect 119798 101284 119840 101324
rect 119512 101275 119880 101284
rect 134632 101324 135000 101333
rect 134672 101284 134714 101324
rect 134754 101284 134796 101324
rect 134836 101284 134878 101324
rect 134918 101284 134960 101324
rect 134632 101275 135000 101284
rect 149752 101324 150120 101333
rect 149792 101284 149834 101324
rect 149874 101284 149916 101324
rect 149956 101284 149998 101324
rect 150038 101284 150080 101324
rect 149752 101275 150120 101284
rect 75392 100568 75760 100577
rect 75432 100528 75474 100568
rect 75514 100528 75556 100568
rect 75596 100528 75638 100568
rect 75678 100528 75720 100568
rect 75392 100519 75760 100528
rect 90512 100568 90880 100577
rect 90552 100528 90594 100568
rect 90634 100528 90676 100568
rect 90716 100528 90758 100568
rect 90798 100528 90840 100568
rect 90512 100519 90880 100528
rect 105632 100568 106000 100577
rect 105672 100528 105714 100568
rect 105754 100528 105796 100568
rect 105836 100528 105878 100568
rect 105918 100528 105960 100568
rect 105632 100519 106000 100528
rect 120752 100568 121120 100577
rect 120792 100528 120834 100568
rect 120874 100528 120916 100568
rect 120956 100528 120998 100568
rect 121038 100528 121080 100568
rect 120752 100519 121120 100528
rect 135872 100568 136240 100577
rect 135912 100528 135954 100568
rect 135994 100528 136036 100568
rect 136076 100528 136118 100568
rect 136158 100528 136200 100568
rect 135872 100519 136240 100528
rect 150992 100568 151360 100577
rect 151032 100528 151074 100568
rect 151114 100528 151156 100568
rect 151196 100528 151238 100568
rect 151278 100528 151320 100568
rect 150992 100519 151360 100528
rect 74152 99812 74520 99821
rect 74192 99772 74234 99812
rect 74274 99772 74316 99812
rect 74356 99772 74398 99812
rect 74438 99772 74480 99812
rect 74152 99763 74520 99772
rect 89272 99812 89640 99821
rect 89312 99772 89354 99812
rect 89394 99772 89436 99812
rect 89476 99772 89518 99812
rect 89558 99772 89600 99812
rect 89272 99763 89640 99772
rect 104392 99812 104760 99821
rect 104432 99772 104474 99812
rect 104514 99772 104556 99812
rect 104596 99772 104638 99812
rect 104678 99772 104720 99812
rect 104392 99763 104760 99772
rect 119512 99812 119880 99821
rect 119552 99772 119594 99812
rect 119634 99772 119676 99812
rect 119716 99772 119758 99812
rect 119798 99772 119840 99812
rect 119512 99763 119880 99772
rect 134632 99812 135000 99821
rect 134672 99772 134714 99812
rect 134754 99772 134796 99812
rect 134836 99772 134878 99812
rect 134918 99772 134960 99812
rect 134632 99763 135000 99772
rect 149752 99812 150120 99821
rect 149792 99772 149834 99812
rect 149874 99772 149916 99812
rect 149956 99772 149998 99812
rect 150038 99772 150080 99812
rect 149752 99763 150120 99772
rect 75392 99056 75760 99065
rect 75432 99016 75474 99056
rect 75514 99016 75556 99056
rect 75596 99016 75638 99056
rect 75678 99016 75720 99056
rect 75392 99007 75760 99016
rect 90512 99056 90880 99065
rect 90552 99016 90594 99056
rect 90634 99016 90676 99056
rect 90716 99016 90758 99056
rect 90798 99016 90840 99056
rect 90512 99007 90880 99016
rect 105632 99056 106000 99065
rect 105672 99016 105714 99056
rect 105754 99016 105796 99056
rect 105836 99016 105878 99056
rect 105918 99016 105960 99056
rect 105632 99007 106000 99016
rect 120752 99056 121120 99065
rect 120792 99016 120834 99056
rect 120874 99016 120916 99056
rect 120956 99016 120998 99056
rect 121038 99016 121080 99056
rect 120752 99007 121120 99016
rect 135872 99056 136240 99065
rect 135912 99016 135954 99056
rect 135994 99016 136036 99056
rect 136076 99016 136118 99056
rect 136158 99016 136200 99056
rect 135872 99007 136240 99016
rect 150992 99056 151360 99065
rect 151032 99016 151074 99056
rect 151114 99016 151156 99056
rect 151196 99016 151238 99056
rect 151278 99016 151320 99056
rect 150992 99007 151360 99016
rect 74152 98300 74520 98309
rect 74192 98260 74234 98300
rect 74274 98260 74316 98300
rect 74356 98260 74398 98300
rect 74438 98260 74480 98300
rect 74152 98251 74520 98260
rect 89272 98300 89640 98309
rect 89312 98260 89354 98300
rect 89394 98260 89436 98300
rect 89476 98260 89518 98300
rect 89558 98260 89600 98300
rect 89272 98251 89640 98260
rect 104392 98300 104760 98309
rect 104432 98260 104474 98300
rect 104514 98260 104556 98300
rect 104596 98260 104638 98300
rect 104678 98260 104720 98300
rect 104392 98251 104760 98260
rect 119512 98300 119880 98309
rect 119552 98260 119594 98300
rect 119634 98260 119676 98300
rect 119716 98260 119758 98300
rect 119798 98260 119840 98300
rect 119512 98251 119880 98260
rect 134632 98300 135000 98309
rect 134672 98260 134714 98300
rect 134754 98260 134796 98300
rect 134836 98260 134878 98300
rect 134918 98260 134960 98300
rect 134632 98251 135000 98260
rect 149752 98300 150120 98309
rect 149792 98260 149834 98300
rect 149874 98260 149916 98300
rect 149956 98260 149998 98300
rect 150038 98260 150080 98300
rect 149752 98251 150120 98260
rect 75392 97544 75760 97553
rect 75432 97504 75474 97544
rect 75514 97504 75556 97544
rect 75596 97504 75638 97544
rect 75678 97504 75720 97544
rect 75392 97495 75760 97504
rect 90512 97544 90880 97553
rect 90552 97504 90594 97544
rect 90634 97504 90676 97544
rect 90716 97504 90758 97544
rect 90798 97504 90840 97544
rect 90512 97495 90880 97504
rect 105632 97544 106000 97553
rect 105672 97504 105714 97544
rect 105754 97504 105796 97544
rect 105836 97504 105878 97544
rect 105918 97504 105960 97544
rect 105632 97495 106000 97504
rect 120752 97544 121120 97553
rect 120792 97504 120834 97544
rect 120874 97504 120916 97544
rect 120956 97504 120998 97544
rect 121038 97504 121080 97544
rect 120752 97495 121120 97504
rect 135872 97544 136240 97553
rect 135912 97504 135954 97544
rect 135994 97504 136036 97544
rect 136076 97504 136118 97544
rect 136158 97504 136200 97544
rect 135872 97495 136240 97504
rect 150992 97544 151360 97553
rect 151032 97504 151074 97544
rect 151114 97504 151156 97544
rect 151196 97504 151238 97544
rect 151278 97504 151320 97544
rect 150992 97495 151360 97504
rect 74152 96788 74520 96797
rect 74192 96748 74234 96788
rect 74274 96748 74316 96788
rect 74356 96748 74398 96788
rect 74438 96748 74480 96788
rect 74152 96739 74520 96748
rect 89272 96788 89640 96797
rect 89312 96748 89354 96788
rect 89394 96748 89436 96788
rect 89476 96748 89518 96788
rect 89558 96748 89600 96788
rect 89272 96739 89640 96748
rect 104392 96788 104760 96797
rect 104432 96748 104474 96788
rect 104514 96748 104556 96788
rect 104596 96748 104638 96788
rect 104678 96748 104720 96788
rect 104392 96739 104760 96748
rect 119512 96788 119880 96797
rect 119552 96748 119594 96788
rect 119634 96748 119676 96788
rect 119716 96748 119758 96788
rect 119798 96748 119840 96788
rect 119512 96739 119880 96748
rect 134632 96788 135000 96797
rect 134672 96748 134714 96788
rect 134754 96748 134796 96788
rect 134836 96748 134878 96788
rect 134918 96748 134960 96788
rect 134632 96739 135000 96748
rect 149752 96788 150120 96797
rect 149792 96748 149834 96788
rect 149874 96748 149916 96788
rect 149956 96748 149998 96788
rect 150038 96748 150080 96788
rect 149752 96739 150120 96748
rect 75392 96032 75760 96041
rect 75432 95992 75474 96032
rect 75514 95992 75556 96032
rect 75596 95992 75638 96032
rect 75678 95992 75720 96032
rect 75392 95983 75760 95992
rect 90512 96032 90880 96041
rect 90552 95992 90594 96032
rect 90634 95992 90676 96032
rect 90716 95992 90758 96032
rect 90798 95992 90840 96032
rect 90512 95983 90880 95992
rect 105632 96032 106000 96041
rect 105672 95992 105714 96032
rect 105754 95992 105796 96032
rect 105836 95992 105878 96032
rect 105918 95992 105960 96032
rect 105632 95983 106000 95992
rect 120752 96032 121120 96041
rect 120792 95992 120834 96032
rect 120874 95992 120916 96032
rect 120956 95992 120998 96032
rect 121038 95992 121080 96032
rect 120752 95983 121120 95992
rect 135872 96032 136240 96041
rect 135912 95992 135954 96032
rect 135994 95992 136036 96032
rect 136076 95992 136118 96032
rect 136158 95992 136200 96032
rect 135872 95983 136240 95992
rect 150992 96032 151360 96041
rect 151032 95992 151074 96032
rect 151114 95992 151156 96032
rect 151196 95992 151238 96032
rect 151278 95992 151320 96032
rect 150992 95983 151360 95992
rect 74152 95276 74520 95285
rect 74192 95236 74234 95276
rect 74274 95236 74316 95276
rect 74356 95236 74398 95276
rect 74438 95236 74480 95276
rect 74152 95227 74520 95236
rect 89272 95276 89640 95285
rect 89312 95236 89354 95276
rect 89394 95236 89436 95276
rect 89476 95236 89518 95276
rect 89558 95236 89600 95276
rect 89272 95227 89640 95236
rect 104392 95276 104760 95285
rect 104432 95236 104474 95276
rect 104514 95236 104556 95276
rect 104596 95236 104638 95276
rect 104678 95236 104720 95276
rect 104392 95227 104760 95236
rect 119512 95276 119880 95285
rect 119552 95236 119594 95276
rect 119634 95236 119676 95276
rect 119716 95236 119758 95276
rect 119798 95236 119840 95276
rect 119512 95227 119880 95236
rect 134632 95276 135000 95285
rect 134672 95236 134714 95276
rect 134754 95236 134796 95276
rect 134836 95236 134878 95276
rect 134918 95236 134960 95276
rect 134632 95227 135000 95236
rect 149752 95276 150120 95285
rect 149792 95236 149834 95276
rect 149874 95236 149916 95276
rect 149956 95236 149998 95276
rect 150038 95236 150080 95276
rect 149752 95227 150120 95236
rect 75392 94520 75760 94529
rect 75432 94480 75474 94520
rect 75514 94480 75556 94520
rect 75596 94480 75638 94520
rect 75678 94480 75720 94520
rect 75392 94471 75760 94480
rect 90512 94520 90880 94529
rect 90552 94480 90594 94520
rect 90634 94480 90676 94520
rect 90716 94480 90758 94520
rect 90798 94480 90840 94520
rect 90512 94471 90880 94480
rect 105632 94520 106000 94529
rect 105672 94480 105714 94520
rect 105754 94480 105796 94520
rect 105836 94480 105878 94520
rect 105918 94480 105960 94520
rect 105632 94471 106000 94480
rect 120752 94520 121120 94529
rect 120792 94480 120834 94520
rect 120874 94480 120916 94520
rect 120956 94480 120998 94520
rect 121038 94480 121080 94520
rect 120752 94471 121120 94480
rect 135872 94520 136240 94529
rect 135912 94480 135954 94520
rect 135994 94480 136036 94520
rect 136076 94480 136118 94520
rect 136158 94480 136200 94520
rect 135872 94471 136240 94480
rect 150992 94520 151360 94529
rect 151032 94480 151074 94520
rect 151114 94480 151156 94520
rect 151196 94480 151238 94520
rect 151278 94480 151320 94520
rect 150992 94471 151360 94480
rect 74152 93764 74520 93773
rect 74192 93724 74234 93764
rect 74274 93724 74316 93764
rect 74356 93724 74398 93764
rect 74438 93724 74480 93764
rect 74152 93715 74520 93724
rect 89272 93764 89640 93773
rect 89312 93724 89354 93764
rect 89394 93724 89436 93764
rect 89476 93724 89518 93764
rect 89558 93724 89600 93764
rect 89272 93715 89640 93724
rect 104392 93764 104760 93773
rect 104432 93724 104474 93764
rect 104514 93724 104556 93764
rect 104596 93724 104638 93764
rect 104678 93724 104720 93764
rect 104392 93715 104760 93724
rect 119512 93764 119880 93773
rect 119552 93724 119594 93764
rect 119634 93724 119676 93764
rect 119716 93724 119758 93764
rect 119798 93724 119840 93764
rect 119512 93715 119880 93724
rect 134632 93764 135000 93773
rect 134672 93724 134714 93764
rect 134754 93724 134796 93764
rect 134836 93724 134878 93764
rect 134918 93724 134960 93764
rect 134632 93715 135000 93724
rect 149752 93764 150120 93773
rect 149792 93724 149834 93764
rect 149874 93724 149916 93764
rect 149956 93724 149998 93764
rect 150038 93724 150080 93764
rect 149752 93715 150120 93724
rect 75392 93008 75760 93017
rect 75432 92968 75474 93008
rect 75514 92968 75556 93008
rect 75596 92968 75638 93008
rect 75678 92968 75720 93008
rect 75392 92959 75760 92968
rect 90512 93008 90880 93017
rect 90552 92968 90594 93008
rect 90634 92968 90676 93008
rect 90716 92968 90758 93008
rect 90798 92968 90840 93008
rect 90512 92959 90880 92968
rect 105632 93008 106000 93017
rect 105672 92968 105714 93008
rect 105754 92968 105796 93008
rect 105836 92968 105878 93008
rect 105918 92968 105960 93008
rect 105632 92959 106000 92968
rect 120752 93008 121120 93017
rect 120792 92968 120834 93008
rect 120874 92968 120916 93008
rect 120956 92968 120998 93008
rect 121038 92968 121080 93008
rect 120752 92959 121120 92968
rect 135872 93008 136240 93017
rect 135912 92968 135954 93008
rect 135994 92968 136036 93008
rect 136076 92968 136118 93008
rect 136158 92968 136200 93008
rect 135872 92959 136240 92968
rect 150992 93008 151360 93017
rect 151032 92968 151074 93008
rect 151114 92968 151156 93008
rect 151196 92968 151238 93008
rect 151278 92968 151320 93008
rect 150992 92959 151360 92968
rect 74152 92252 74520 92261
rect 74192 92212 74234 92252
rect 74274 92212 74316 92252
rect 74356 92212 74398 92252
rect 74438 92212 74480 92252
rect 74152 92203 74520 92212
rect 89272 92252 89640 92261
rect 89312 92212 89354 92252
rect 89394 92212 89436 92252
rect 89476 92212 89518 92252
rect 89558 92212 89600 92252
rect 89272 92203 89640 92212
rect 104392 92252 104760 92261
rect 104432 92212 104474 92252
rect 104514 92212 104556 92252
rect 104596 92212 104638 92252
rect 104678 92212 104720 92252
rect 104392 92203 104760 92212
rect 119512 92252 119880 92261
rect 119552 92212 119594 92252
rect 119634 92212 119676 92252
rect 119716 92212 119758 92252
rect 119798 92212 119840 92252
rect 119512 92203 119880 92212
rect 134632 92252 135000 92261
rect 134672 92212 134714 92252
rect 134754 92212 134796 92252
rect 134836 92212 134878 92252
rect 134918 92212 134960 92252
rect 134632 92203 135000 92212
rect 149752 92252 150120 92261
rect 149792 92212 149834 92252
rect 149874 92212 149916 92252
rect 149956 92212 149998 92252
rect 150038 92212 150080 92252
rect 149752 92203 150120 92212
rect 75392 91496 75760 91505
rect 75432 91456 75474 91496
rect 75514 91456 75556 91496
rect 75596 91456 75638 91496
rect 75678 91456 75720 91496
rect 75392 91447 75760 91456
rect 90512 91496 90880 91505
rect 90552 91456 90594 91496
rect 90634 91456 90676 91496
rect 90716 91456 90758 91496
rect 90798 91456 90840 91496
rect 90512 91447 90880 91456
rect 105632 91496 106000 91505
rect 105672 91456 105714 91496
rect 105754 91456 105796 91496
rect 105836 91456 105878 91496
rect 105918 91456 105960 91496
rect 105632 91447 106000 91456
rect 120752 91496 121120 91505
rect 120792 91456 120834 91496
rect 120874 91456 120916 91496
rect 120956 91456 120998 91496
rect 121038 91456 121080 91496
rect 120752 91447 121120 91456
rect 135872 91496 136240 91505
rect 135912 91456 135954 91496
rect 135994 91456 136036 91496
rect 136076 91456 136118 91496
rect 136158 91456 136200 91496
rect 135872 91447 136240 91456
rect 150992 91496 151360 91505
rect 151032 91456 151074 91496
rect 151114 91456 151156 91496
rect 151196 91456 151238 91496
rect 151278 91456 151320 91496
rect 150992 91447 151360 91456
rect 74152 90740 74520 90749
rect 74192 90700 74234 90740
rect 74274 90700 74316 90740
rect 74356 90700 74398 90740
rect 74438 90700 74480 90740
rect 74152 90691 74520 90700
rect 89272 90740 89640 90749
rect 89312 90700 89354 90740
rect 89394 90700 89436 90740
rect 89476 90700 89518 90740
rect 89558 90700 89600 90740
rect 89272 90691 89640 90700
rect 104392 90740 104760 90749
rect 104432 90700 104474 90740
rect 104514 90700 104556 90740
rect 104596 90700 104638 90740
rect 104678 90700 104720 90740
rect 104392 90691 104760 90700
rect 119512 90740 119880 90749
rect 119552 90700 119594 90740
rect 119634 90700 119676 90740
rect 119716 90700 119758 90740
rect 119798 90700 119840 90740
rect 119512 90691 119880 90700
rect 134632 90740 135000 90749
rect 134672 90700 134714 90740
rect 134754 90700 134796 90740
rect 134836 90700 134878 90740
rect 134918 90700 134960 90740
rect 134632 90691 135000 90700
rect 149752 90740 150120 90749
rect 149792 90700 149834 90740
rect 149874 90700 149916 90740
rect 149956 90700 149998 90740
rect 150038 90700 150080 90740
rect 149752 90691 150120 90700
rect 75392 89984 75760 89993
rect 75432 89944 75474 89984
rect 75514 89944 75556 89984
rect 75596 89944 75638 89984
rect 75678 89944 75720 89984
rect 75392 89935 75760 89944
rect 90512 89984 90880 89993
rect 90552 89944 90594 89984
rect 90634 89944 90676 89984
rect 90716 89944 90758 89984
rect 90798 89944 90840 89984
rect 90512 89935 90880 89944
rect 105632 89984 106000 89993
rect 105672 89944 105714 89984
rect 105754 89944 105796 89984
rect 105836 89944 105878 89984
rect 105918 89944 105960 89984
rect 105632 89935 106000 89944
rect 120752 89984 121120 89993
rect 120792 89944 120834 89984
rect 120874 89944 120916 89984
rect 120956 89944 120998 89984
rect 121038 89944 121080 89984
rect 120752 89935 121120 89944
rect 135872 89984 136240 89993
rect 135912 89944 135954 89984
rect 135994 89944 136036 89984
rect 136076 89944 136118 89984
rect 136158 89944 136200 89984
rect 135872 89935 136240 89944
rect 150992 89984 151360 89993
rect 151032 89944 151074 89984
rect 151114 89944 151156 89984
rect 151196 89944 151238 89984
rect 151278 89944 151320 89984
rect 150992 89935 151360 89944
rect 74152 89228 74520 89237
rect 74192 89188 74234 89228
rect 74274 89188 74316 89228
rect 74356 89188 74398 89228
rect 74438 89188 74480 89228
rect 74152 89179 74520 89188
rect 89272 89228 89640 89237
rect 89312 89188 89354 89228
rect 89394 89188 89436 89228
rect 89476 89188 89518 89228
rect 89558 89188 89600 89228
rect 89272 89179 89640 89188
rect 104392 89228 104760 89237
rect 104432 89188 104474 89228
rect 104514 89188 104556 89228
rect 104596 89188 104638 89228
rect 104678 89188 104720 89228
rect 104392 89179 104760 89188
rect 119512 89228 119880 89237
rect 119552 89188 119594 89228
rect 119634 89188 119676 89228
rect 119716 89188 119758 89228
rect 119798 89188 119840 89228
rect 119512 89179 119880 89188
rect 134632 89228 135000 89237
rect 134672 89188 134714 89228
rect 134754 89188 134796 89228
rect 134836 89188 134878 89228
rect 134918 89188 134960 89228
rect 134632 89179 135000 89188
rect 149752 89228 150120 89237
rect 149792 89188 149834 89228
rect 149874 89188 149916 89228
rect 149956 89188 149998 89228
rect 150038 89188 150080 89228
rect 149752 89179 150120 89188
rect 75392 88472 75760 88481
rect 75432 88432 75474 88472
rect 75514 88432 75556 88472
rect 75596 88432 75638 88472
rect 75678 88432 75720 88472
rect 75392 88423 75760 88432
rect 90512 88472 90880 88481
rect 90552 88432 90594 88472
rect 90634 88432 90676 88472
rect 90716 88432 90758 88472
rect 90798 88432 90840 88472
rect 90512 88423 90880 88432
rect 105632 88472 106000 88481
rect 105672 88432 105714 88472
rect 105754 88432 105796 88472
rect 105836 88432 105878 88472
rect 105918 88432 105960 88472
rect 105632 88423 106000 88432
rect 120752 88472 121120 88481
rect 120792 88432 120834 88472
rect 120874 88432 120916 88472
rect 120956 88432 120998 88472
rect 121038 88432 121080 88472
rect 120752 88423 121120 88432
rect 135872 88472 136240 88481
rect 135912 88432 135954 88472
rect 135994 88432 136036 88472
rect 136076 88432 136118 88472
rect 136158 88432 136200 88472
rect 135872 88423 136240 88432
rect 150992 88472 151360 88481
rect 151032 88432 151074 88472
rect 151114 88432 151156 88472
rect 151196 88432 151238 88472
rect 151278 88432 151320 88472
rect 150992 88423 151360 88432
rect 74152 87716 74520 87725
rect 74192 87676 74234 87716
rect 74274 87676 74316 87716
rect 74356 87676 74398 87716
rect 74438 87676 74480 87716
rect 74152 87667 74520 87676
rect 89272 87716 89640 87725
rect 89312 87676 89354 87716
rect 89394 87676 89436 87716
rect 89476 87676 89518 87716
rect 89558 87676 89600 87716
rect 89272 87667 89640 87676
rect 104392 87716 104760 87725
rect 104432 87676 104474 87716
rect 104514 87676 104556 87716
rect 104596 87676 104638 87716
rect 104678 87676 104720 87716
rect 104392 87667 104760 87676
rect 119512 87716 119880 87725
rect 119552 87676 119594 87716
rect 119634 87676 119676 87716
rect 119716 87676 119758 87716
rect 119798 87676 119840 87716
rect 119512 87667 119880 87676
rect 134632 87716 135000 87725
rect 134672 87676 134714 87716
rect 134754 87676 134796 87716
rect 134836 87676 134878 87716
rect 134918 87676 134960 87716
rect 134632 87667 135000 87676
rect 149752 87716 150120 87725
rect 149792 87676 149834 87716
rect 149874 87676 149916 87716
rect 149956 87676 149998 87716
rect 150038 87676 150080 87716
rect 149752 87667 150120 87676
rect 75392 86960 75760 86969
rect 75432 86920 75474 86960
rect 75514 86920 75556 86960
rect 75596 86920 75638 86960
rect 75678 86920 75720 86960
rect 75392 86911 75760 86920
rect 90512 86960 90880 86969
rect 90552 86920 90594 86960
rect 90634 86920 90676 86960
rect 90716 86920 90758 86960
rect 90798 86920 90840 86960
rect 90512 86911 90880 86920
rect 105632 86960 106000 86969
rect 105672 86920 105714 86960
rect 105754 86920 105796 86960
rect 105836 86920 105878 86960
rect 105918 86920 105960 86960
rect 105632 86911 106000 86920
rect 120752 86960 121120 86969
rect 120792 86920 120834 86960
rect 120874 86920 120916 86960
rect 120956 86920 120998 86960
rect 121038 86920 121080 86960
rect 120752 86911 121120 86920
rect 135872 86960 136240 86969
rect 135912 86920 135954 86960
rect 135994 86920 136036 86960
rect 136076 86920 136118 86960
rect 136158 86920 136200 86960
rect 135872 86911 136240 86920
rect 150992 86960 151360 86969
rect 151032 86920 151074 86960
rect 151114 86920 151156 86960
rect 151196 86920 151238 86960
rect 151278 86920 151320 86960
rect 150992 86911 151360 86920
rect 74152 86204 74520 86213
rect 74192 86164 74234 86204
rect 74274 86164 74316 86204
rect 74356 86164 74398 86204
rect 74438 86164 74480 86204
rect 74152 86155 74520 86164
rect 89272 86204 89640 86213
rect 89312 86164 89354 86204
rect 89394 86164 89436 86204
rect 89476 86164 89518 86204
rect 89558 86164 89600 86204
rect 89272 86155 89640 86164
rect 104392 86204 104760 86213
rect 104432 86164 104474 86204
rect 104514 86164 104556 86204
rect 104596 86164 104638 86204
rect 104678 86164 104720 86204
rect 104392 86155 104760 86164
rect 119512 86204 119880 86213
rect 119552 86164 119594 86204
rect 119634 86164 119676 86204
rect 119716 86164 119758 86204
rect 119798 86164 119840 86204
rect 119512 86155 119880 86164
rect 134632 86204 135000 86213
rect 134672 86164 134714 86204
rect 134754 86164 134796 86204
rect 134836 86164 134878 86204
rect 134918 86164 134960 86204
rect 134632 86155 135000 86164
rect 149752 86204 150120 86213
rect 149792 86164 149834 86204
rect 149874 86164 149916 86204
rect 149956 86164 149998 86204
rect 150038 86164 150080 86204
rect 149752 86155 150120 86164
rect 75392 85448 75760 85457
rect 75432 85408 75474 85448
rect 75514 85408 75556 85448
rect 75596 85408 75638 85448
rect 75678 85408 75720 85448
rect 75392 85399 75760 85408
rect 90512 85448 90880 85457
rect 90552 85408 90594 85448
rect 90634 85408 90676 85448
rect 90716 85408 90758 85448
rect 90798 85408 90840 85448
rect 90512 85399 90880 85408
rect 105632 85448 106000 85457
rect 105672 85408 105714 85448
rect 105754 85408 105796 85448
rect 105836 85408 105878 85448
rect 105918 85408 105960 85448
rect 105632 85399 106000 85408
rect 120752 85448 121120 85457
rect 120792 85408 120834 85448
rect 120874 85408 120916 85448
rect 120956 85408 120998 85448
rect 121038 85408 121080 85448
rect 120752 85399 121120 85408
rect 135872 85448 136240 85457
rect 135912 85408 135954 85448
rect 135994 85408 136036 85448
rect 136076 85408 136118 85448
rect 136158 85408 136200 85448
rect 135872 85399 136240 85408
rect 150992 85448 151360 85457
rect 151032 85408 151074 85448
rect 151114 85408 151156 85448
rect 151196 85408 151238 85448
rect 151278 85408 151320 85448
rect 150992 85399 151360 85408
rect 74152 84692 74520 84701
rect 74192 84652 74234 84692
rect 74274 84652 74316 84692
rect 74356 84652 74398 84692
rect 74438 84652 74480 84692
rect 74152 84643 74520 84652
rect 89272 84692 89640 84701
rect 89312 84652 89354 84692
rect 89394 84652 89436 84692
rect 89476 84652 89518 84692
rect 89558 84652 89600 84692
rect 89272 84643 89640 84652
rect 104392 84692 104760 84701
rect 104432 84652 104474 84692
rect 104514 84652 104556 84692
rect 104596 84652 104638 84692
rect 104678 84652 104720 84692
rect 104392 84643 104760 84652
rect 119512 84692 119880 84701
rect 119552 84652 119594 84692
rect 119634 84652 119676 84692
rect 119716 84652 119758 84692
rect 119798 84652 119840 84692
rect 119512 84643 119880 84652
rect 134632 84692 135000 84701
rect 134672 84652 134714 84692
rect 134754 84652 134796 84692
rect 134836 84652 134878 84692
rect 134918 84652 134960 84692
rect 134632 84643 135000 84652
rect 149752 84692 150120 84701
rect 149792 84652 149834 84692
rect 149874 84652 149916 84692
rect 149956 84652 149998 84692
rect 150038 84652 150080 84692
rect 149752 84643 150120 84652
rect 75392 83936 75760 83945
rect 75432 83896 75474 83936
rect 75514 83896 75556 83936
rect 75596 83896 75638 83936
rect 75678 83896 75720 83936
rect 75392 83887 75760 83896
rect 90512 83936 90880 83945
rect 90552 83896 90594 83936
rect 90634 83896 90676 83936
rect 90716 83896 90758 83936
rect 90798 83896 90840 83936
rect 90512 83887 90880 83896
rect 105632 83936 106000 83945
rect 105672 83896 105714 83936
rect 105754 83896 105796 83936
rect 105836 83896 105878 83936
rect 105918 83896 105960 83936
rect 105632 83887 106000 83896
rect 120752 83936 121120 83945
rect 120792 83896 120834 83936
rect 120874 83896 120916 83936
rect 120956 83896 120998 83936
rect 121038 83896 121080 83936
rect 120752 83887 121120 83896
rect 135872 83936 136240 83945
rect 135912 83896 135954 83936
rect 135994 83896 136036 83936
rect 136076 83896 136118 83936
rect 136158 83896 136200 83936
rect 135872 83887 136240 83896
rect 150992 83936 151360 83945
rect 151032 83896 151074 83936
rect 151114 83896 151156 83936
rect 151196 83896 151238 83936
rect 151278 83896 151320 83936
rect 150992 83887 151360 83896
rect 74152 83180 74520 83189
rect 74192 83140 74234 83180
rect 74274 83140 74316 83180
rect 74356 83140 74398 83180
rect 74438 83140 74480 83180
rect 74152 83131 74520 83140
rect 89272 83180 89640 83189
rect 89312 83140 89354 83180
rect 89394 83140 89436 83180
rect 89476 83140 89518 83180
rect 89558 83140 89600 83180
rect 89272 83131 89640 83140
rect 104392 83180 104760 83189
rect 104432 83140 104474 83180
rect 104514 83140 104556 83180
rect 104596 83140 104638 83180
rect 104678 83140 104720 83180
rect 104392 83131 104760 83140
rect 119512 83180 119880 83189
rect 119552 83140 119594 83180
rect 119634 83140 119676 83180
rect 119716 83140 119758 83180
rect 119798 83140 119840 83180
rect 119512 83131 119880 83140
rect 134632 83180 135000 83189
rect 134672 83140 134714 83180
rect 134754 83140 134796 83180
rect 134836 83140 134878 83180
rect 134918 83140 134960 83180
rect 134632 83131 135000 83140
rect 149752 83180 150120 83189
rect 149792 83140 149834 83180
rect 149874 83140 149916 83180
rect 149956 83140 149998 83180
rect 150038 83140 150080 83180
rect 149752 83131 150120 83140
rect 75392 82424 75760 82433
rect 75432 82384 75474 82424
rect 75514 82384 75556 82424
rect 75596 82384 75638 82424
rect 75678 82384 75720 82424
rect 75392 82375 75760 82384
rect 90512 82424 90880 82433
rect 90552 82384 90594 82424
rect 90634 82384 90676 82424
rect 90716 82384 90758 82424
rect 90798 82384 90840 82424
rect 90512 82375 90880 82384
rect 105632 82424 106000 82433
rect 105672 82384 105714 82424
rect 105754 82384 105796 82424
rect 105836 82384 105878 82424
rect 105918 82384 105960 82424
rect 105632 82375 106000 82384
rect 120752 82424 121120 82433
rect 120792 82384 120834 82424
rect 120874 82384 120916 82424
rect 120956 82384 120998 82424
rect 121038 82384 121080 82424
rect 120752 82375 121120 82384
rect 135872 82424 136240 82433
rect 135912 82384 135954 82424
rect 135994 82384 136036 82424
rect 136076 82384 136118 82424
rect 136158 82384 136200 82424
rect 135872 82375 136240 82384
rect 150992 82424 151360 82433
rect 151032 82384 151074 82424
rect 151114 82384 151156 82424
rect 151196 82384 151238 82424
rect 151278 82384 151320 82424
rect 150992 82375 151360 82384
rect 74152 81668 74520 81677
rect 74192 81628 74234 81668
rect 74274 81628 74316 81668
rect 74356 81628 74398 81668
rect 74438 81628 74480 81668
rect 74152 81619 74520 81628
rect 89272 81668 89640 81677
rect 89312 81628 89354 81668
rect 89394 81628 89436 81668
rect 89476 81628 89518 81668
rect 89558 81628 89600 81668
rect 89272 81619 89640 81628
rect 104392 81668 104760 81677
rect 104432 81628 104474 81668
rect 104514 81628 104556 81668
rect 104596 81628 104638 81668
rect 104678 81628 104720 81668
rect 104392 81619 104760 81628
rect 119512 81668 119880 81677
rect 119552 81628 119594 81668
rect 119634 81628 119676 81668
rect 119716 81628 119758 81668
rect 119798 81628 119840 81668
rect 119512 81619 119880 81628
rect 134632 81668 135000 81677
rect 134672 81628 134714 81668
rect 134754 81628 134796 81668
rect 134836 81628 134878 81668
rect 134918 81628 134960 81668
rect 134632 81619 135000 81628
rect 149752 81668 150120 81677
rect 149792 81628 149834 81668
rect 149874 81628 149916 81668
rect 149956 81628 149998 81668
rect 150038 81628 150080 81668
rect 149752 81619 150120 81628
rect 75392 80912 75760 80921
rect 75432 80872 75474 80912
rect 75514 80872 75556 80912
rect 75596 80872 75638 80912
rect 75678 80872 75720 80912
rect 75392 80863 75760 80872
rect 90512 80912 90880 80921
rect 90552 80872 90594 80912
rect 90634 80872 90676 80912
rect 90716 80872 90758 80912
rect 90798 80872 90840 80912
rect 90512 80863 90880 80872
rect 105632 80912 106000 80921
rect 105672 80872 105714 80912
rect 105754 80872 105796 80912
rect 105836 80872 105878 80912
rect 105918 80872 105960 80912
rect 105632 80863 106000 80872
rect 120752 80912 121120 80921
rect 120792 80872 120834 80912
rect 120874 80872 120916 80912
rect 120956 80872 120998 80912
rect 121038 80872 121080 80912
rect 120752 80863 121120 80872
rect 135872 80912 136240 80921
rect 135912 80872 135954 80912
rect 135994 80872 136036 80912
rect 136076 80872 136118 80912
rect 136158 80872 136200 80912
rect 135872 80863 136240 80872
rect 150992 80912 151360 80921
rect 151032 80872 151074 80912
rect 151114 80872 151156 80912
rect 151196 80872 151238 80912
rect 151278 80872 151320 80912
rect 150992 80863 151360 80872
rect 74152 80156 74520 80165
rect 74192 80116 74234 80156
rect 74274 80116 74316 80156
rect 74356 80116 74398 80156
rect 74438 80116 74480 80156
rect 74152 80107 74520 80116
rect 89272 80156 89640 80165
rect 89312 80116 89354 80156
rect 89394 80116 89436 80156
rect 89476 80116 89518 80156
rect 89558 80116 89600 80156
rect 89272 80107 89640 80116
rect 104392 80156 104760 80165
rect 104432 80116 104474 80156
rect 104514 80116 104556 80156
rect 104596 80116 104638 80156
rect 104678 80116 104720 80156
rect 104392 80107 104760 80116
rect 119512 80156 119880 80165
rect 119552 80116 119594 80156
rect 119634 80116 119676 80156
rect 119716 80116 119758 80156
rect 119798 80116 119840 80156
rect 119512 80107 119880 80116
rect 134632 80156 135000 80165
rect 134672 80116 134714 80156
rect 134754 80116 134796 80156
rect 134836 80116 134878 80156
rect 134918 80116 134960 80156
rect 134632 80107 135000 80116
rect 149752 80156 150120 80165
rect 149792 80116 149834 80156
rect 149874 80116 149916 80156
rect 149956 80116 149998 80156
rect 150038 80116 150080 80156
rect 149752 80107 150120 80116
rect 75392 79400 75760 79409
rect 75432 79360 75474 79400
rect 75514 79360 75556 79400
rect 75596 79360 75638 79400
rect 75678 79360 75720 79400
rect 75392 79351 75760 79360
rect 90512 79400 90880 79409
rect 90552 79360 90594 79400
rect 90634 79360 90676 79400
rect 90716 79360 90758 79400
rect 90798 79360 90840 79400
rect 90512 79351 90880 79360
rect 105632 79400 106000 79409
rect 105672 79360 105714 79400
rect 105754 79360 105796 79400
rect 105836 79360 105878 79400
rect 105918 79360 105960 79400
rect 105632 79351 106000 79360
rect 120752 79400 121120 79409
rect 120792 79360 120834 79400
rect 120874 79360 120916 79400
rect 120956 79360 120998 79400
rect 121038 79360 121080 79400
rect 120752 79351 121120 79360
rect 135872 79400 136240 79409
rect 135912 79360 135954 79400
rect 135994 79360 136036 79400
rect 136076 79360 136118 79400
rect 136158 79360 136200 79400
rect 135872 79351 136240 79360
rect 150992 79400 151360 79409
rect 151032 79360 151074 79400
rect 151114 79360 151156 79400
rect 151196 79360 151238 79400
rect 151278 79360 151320 79400
rect 150992 79351 151360 79360
rect 74152 78644 74520 78653
rect 74192 78604 74234 78644
rect 74274 78604 74316 78644
rect 74356 78604 74398 78644
rect 74438 78604 74480 78644
rect 74152 78595 74520 78604
rect 89272 78644 89640 78653
rect 89312 78604 89354 78644
rect 89394 78604 89436 78644
rect 89476 78604 89518 78644
rect 89558 78604 89600 78644
rect 89272 78595 89640 78604
rect 104392 78644 104760 78653
rect 104432 78604 104474 78644
rect 104514 78604 104556 78644
rect 104596 78604 104638 78644
rect 104678 78604 104720 78644
rect 104392 78595 104760 78604
rect 119512 78644 119880 78653
rect 119552 78604 119594 78644
rect 119634 78604 119676 78644
rect 119716 78604 119758 78644
rect 119798 78604 119840 78644
rect 119512 78595 119880 78604
rect 134632 78644 135000 78653
rect 134672 78604 134714 78644
rect 134754 78604 134796 78644
rect 134836 78604 134878 78644
rect 134918 78604 134960 78644
rect 134632 78595 135000 78604
rect 149752 78644 150120 78653
rect 149792 78604 149834 78644
rect 149874 78604 149916 78644
rect 149956 78604 149998 78644
rect 150038 78604 150080 78644
rect 149752 78595 150120 78604
rect 75392 77888 75760 77897
rect 75432 77848 75474 77888
rect 75514 77848 75556 77888
rect 75596 77848 75638 77888
rect 75678 77848 75720 77888
rect 75392 77839 75760 77848
rect 90512 77888 90880 77897
rect 90552 77848 90594 77888
rect 90634 77848 90676 77888
rect 90716 77848 90758 77888
rect 90798 77848 90840 77888
rect 90512 77839 90880 77848
rect 105632 77888 106000 77897
rect 105672 77848 105714 77888
rect 105754 77848 105796 77888
rect 105836 77848 105878 77888
rect 105918 77848 105960 77888
rect 105632 77839 106000 77848
rect 120752 77888 121120 77897
rect 120792 77848 120834 77888
rect 120874 77848 120916 77888
rect 120956 77848 120998 77888
rect 121038 77848 121080 77888
rect 120752 77839 121120 77848
rect 135872 77888 136240 77897
rect 135912 77848 135954 77888
rect 135994 77848 136036 77888
rect 136076 77848 136118 77888
rect 136158 77848 136200 77888
rect 135872 77839 136240 77848
rect 150992 77888 151360 77897
rect 151032 77848 151074 77888
rect 151114 77848 151156 77888
rect 151196 77848 151238 77888
rect 151278 77848 151320 77888
rect 150992 77839 151360 77848
rect 74152 77132 74520 77141
rect 74192 77092 74234 77132
rect 74274 77092 74316 77132
rect 74356 77092 74398 77132
rect 74438 77092 74480 77132
rect 74152 77083 74520 77092
rect 89272 77132 89640 77141
rect 89312 77092 89354 77132
rect 89394 77092 89436 77132
rect 89476 77092 89518 77132
rect 89558 77092 89600 77132
rect 89272 77083 89640 77092
rect 104392 77132 104760 77141
rect 104432 77092 104474 77132
rect 104514 77092 104556 77132
rect 104596 77092 104638 77132
rect 104678 77092 104720 77132
rect 104392 77083 104760 77092
rect 119512 77132 119880 77141
rect 119552 77092 119594 77132
rect 119634 77092 119676 77132
rect 119716 77092 119758 77132
rect 119798 77092 119840 77132
rect 119512 77083 119880 77092
rect 134632 77132 135000 77141
rect 134672 77092 134714 77132
rect 134754 77092 134796 77132
rect 134836 77092 134878 77132
rect 134918 77092 134960 77132
rect 134632 77083 135000 77092
rect 149752 77132 150120 77141
rect 149792 77092 149834 77132
rect 149874 77092 149916 77132
rect 149956 77092 149998 77132
rect 150038 77092 150080 77132
rect 149752 77083 150120 77092
rect 75392 76376 75760 76385
rect 75432 76336 75474 76376
rect 75514 76336 75556 76376
rect 75596 76336 75638 76376
rect 75678 76336 75720 76376
rect 75392 76327 75760 76336
rect 90512 76376 90880 76385
rect 90552 76336 90594 76376
rect 90634 76336 90676 76376
rect 90716 76336 90758 76376
rect 90798 76336 90840 76376
rect 90512 76327 90880 76336
rect 105632 76376 106000 76385
rect 105672 76336 105714 76376
rect 105754 76336 105796 76376
rect 105836 76336 105878 76376
rect 105918 76336 105960 76376
rect 105632 76327 106000 76336
rect 120752 76376 121120 76385
rect 120792 76336 120834 76376
rect 120874 76336 120916 76376
rect 120956 76336 120998 76376
rect 121038 76336 121080 76376
rect 120752 76327 121120 76336
rect 135872 76376 136240 76385
rect 135912 76336 135954 76376
rect 135994 76336 136036 76376
rect 136076 76336 136118 76376
rect 136158 76336 136200 76376
rect 135872 76327 136240 76336
rect 150992 76376 151360 76385
rect 151032 76336 151074 76376
rect 151114 76336 151156 76376
rect 151196 76336 151238 76376
rect 151278 76336 151320 76376
rect 150992 76327 151360 76336
rect 74152 75620 74520 75629
rect 74192 75580 74234 75620
rect 74274 75580 74316 75620
rect 74356 75580 74398 75620
rect 74438 75580 74480 75620
rect 74152 75571 74520 75580
rect 89272 75620 89640 75629
rect 89312 75580 89354 75620
rect 89394 75580 89436 75620
rect 89476 75580 89518 75620
rect 89558 75580 89600 75620
rect 89272 75571 89640 75580
rect 104392 75620 104760 75629
rect 104432 75580 104474 75620
rect 104514 75580 104556 75620
rect 104596 75580 104638 75620
rect 104678 75580 104720 75620
rect 104392 75571 104760 75580
rect 119512 75620 119880 75629
rect 119552 75580 119594 75620
rect 119634 75580 119676 75620
rect 119716 75580 119758 75620
rect 119798 75580 119840 75620
rect 119512 75571 119880 75580
rect 134632 75620 135000 75629
rect 134672 75580 134714 75620
rect 134754 75580 134796 75620
rect 134836 75580 134878 75620
rect 134918 75580 134960 75620
rect 134632 75571 135000 75580
rect 149752 75620 150120 75629
rect 149792 75580 149834 75620
rect 149874 75580 149916 75620
rect 149956 75580 149998 75620
rect 150038 75580 150080 75620
rect 149752 75571 150120 75580
rect 75392 74864 75760 74873
rect 75432 74824 75474 74864
rect 75514 74824 75556 74864
rect 75596 74824 75638 74864
rect 75678 74824 75720 74864
rect 75392 74815 75760 74824
rect 90512 74864 90880 74873
rect 90552 74824 90594 74864
rect 90634 74824 90676 74864
rect 90716 74824 90758 74864
rect 90798 74824 90840 74864
rect 90512 74815 90880 74824
rect 105632 74864 106000 74873
rect 105672 74824 105714 74864
rect 105754 74824 105796 74864
rect 105836 74824 105878 74864
rect 105918 74824 105960 74864
rect 105632 74815 106000 74824
rect 120752 74864 121120 74873
rect 120792 74824 120834 74864
rect 120874 74824 120916 74864
rect 120956 74824 120998 74864
rect 121038 74824 121080 74864
rect 120752 74815 121120 74824
rect 135872 74864 136240 74873
rect 135912 74824 135954 74864
rect 135994 74824 136036 74864
rect 136076 74824 136118 74864
rect 136158 74824 136200 74864
rect 135872 74815 136240 74824
rect 150992 74864 151360 74873
rect 151032 74824 151074 74864
rect 151114 74824 151156 74864
rect 151196 74824 151238 74864
rect 151278 74824 151320 74864
rect 150992 74815 151360 74824
rect 74152 74108 74520 74117
rect 74192 74068 74234 74108
rect 74274 74068 74316 74108
rect 74356 74068 74398 74108
rect 74438 74068 74480 74108
rect 74152 74059 74520 74068
rect 89272 74108 89640 74117
rect 89312 74068 89354 74108
rect 89394 74068 89436 74108
rect 89476 74068 89518 74108
rect 89558 74068 89600 74108
rect 89272 74059 89640 74068
rect 104392 74108 104760 74117
rect 104432 74068 104474 74108
rect 104514 74068 104556 74108
rect 104596 74068 104638 74108
rect 104678 74068 104720 74108
rect 104392 74059 104760 74068
rect 119512 74108 119880 74117
rect 119552 74068 119594 74108
rect 119634 74068 119676 74108
rect 119716 74068 119758 74108
rect 119798 74068 119840 74108
rect 119512 74059 119880 74068
rect 134632 74108 135000 74117
rect 134672 74068 134714 74108
rect 134754 74068 134796 74108
rect 134836 74068 134878 74108
rect 134918 74068 134960 74108
rect 134632 74059 135000 74068
rect 149752 74108 150120 74117
rect 149792 74068 149834 74108
rect 149874 74068 149916 74108
rect 149956 74068 149998 74108
rect 150038 74068 150080 74108
rect 149752 74059 150120 74068
rect 75392 73352 75760 73361
rect 75432 73312 75474 73352
rect 75514 73312 75556 73352
rect 75596 73312 75638 73352
rect 75678 73312 75720 73352
rect 75392 73303 75760 73312
rect 90512 73352 90880 73361
rect 90552 73312 90594 73352
rect 90634 73312 90676 73352
rect 90716 73312 90758 73352
rect 90798 73312 90840 73352
rect 90512 73303 90880 73312
rect 105632 73352 106000 73361
rect 105672 73312 105714 73352
rect 105754 73312 105796 73352
rect 105836 73312 105878 73352
rect 105918 73312 105960 73352
rect 105632 73303 106000 73312
rect 120752 73352 121120 73361
rect 120792 73312 120834 73352
rect 120874 73312 120916 73352
rect 120956 73312 120998 73352
rect 121038 73312 121080 73352
rect 120752 73303 121120 73312
rect 135872 73352 136240 73361
rect 135912 73312 135954 73352
rect 135994 73312 136036 73352
rect 136076 73312 136118 73352
rect 136158 73312 136200 73352
rect 135872 73303 136240 73312
rect 150992 73352 151360 73361
rect 151032 73312 151074 73352
rect 151114 73312 151156 73352
rect 151196 73312 151238 73352
rect 151278 73312 151320 73352
rect 150992 73303 151360 73312
rect 74152 72596 74520 72605
rect 74192 72556 74234 72596
rect 74274 72556 74316 72596
rect 74356 72556 74398 72596
rect 74438 72556 74480 72596
rect 74152 72547 74520 72556
rect 89272 72596 89640 72605
rect 89312 72556 89354 72596
rect 89394 72556 89436 72596
rect 89476 72556 89518 72596
rect 89558 72556 89600 72596
rect 89272 72547 89640 72556
rect 104392 72596 104760 72605
rect 104432 72556 104474 72596
rect 104514 72556 104556 72596
rect 104596 72556 104638 72596
rect 104678 72556 104720 72596
rect 104392 72547 104760 72556
rect 119512 72596 119880 72605
rect 119552 72556 119594 72596
rect 119634 72556 119676 72596
rect 119716 72556 119758 72596
rect 119798 72556 119840 72596
rect 119512 72547 119880 72556
rect 134632 72596 135000 72605
rect 134672 72556 134714 72596
rect 134754 72556 134796 72596
rect 134836 72556 134878 72596
rect 134918 72556 134960 72596
rect 134632 72547 135000 72556
rect 149752 72596 150120 72605
rect 149792 72556 149834 72596
rect 149874 72556 149916 72596
rect 149956 72556 149998 72596
rect 150038 72556 150080 72596
rect 149752 72547 150120 72556
rect 75392 71840 75760 71849
rect 75432 71800 75474 71840
rect 75514 71800 75556 71840
rect 75596 71800 75638 71840
rect 75678 71800 75720 71840
rect 75392 71791 75760 71800
rect 90512 71840 90880 71849
rect 90552 71800 90594 71840
rect 90634 71800 90676 71840
rect 90716 71800 90758 71840
rect 90798 71800 90840 71840
rect 90512 71791 90880 71800
rect 105632 71840 106000 71849
rect 105672 71800 105714 71840
rect 105754 71800 105796 71840
rect 105836 71800 105878 71840
rect 105918 71800 105960 71840
rect 105632 71791 106000 71800
rect 120752 71840 121120 71849
rect 120792 71800 120834 71840
rect 120874 71800 120916 71840
rect 120956 71800 120998 71840
rect 121038 71800 121080 71840
rect 120752 71791 121120 71800
rect 135872 71840 136240 71849
rect 135912 71800 135954 71840
rect 135994 71800 136036 71840
rect 136076 71800 136118 71840
rect 136158 71800 136200 71840
rect 135872 71791 136240 71800
rect 150992 71840 151360 71849
rect 151032 71800 151074 71840
rect 151114 71800 151156 71840
rect 151196 71800 151238 71840
rect 151278 71800 151320 71840
rect 150992 71791 151360 71800
<< via4 >>
rect 75392 151936 75432 151976
rect 75474 151936 75514 151976
rect 75556 151936 75596 151976
rect 75638 151936 75678 151976
rect 75720 151936 75760 151976
rect 90512 151936 90552 151976
rect 90594 151936 90634 151976
rect 90676 151936 90716 151976
rect 90758 151936 90798 151976
rect 90840 151936 90880 151976
rect 105632 151936 105672 151976
rect 105714 151936 105754 151976
rect 105796 151936 105836 151976
rect 105878 151936 105918 151976
rect 105960 151936 106000 151976
rect 120752 151936 120792 151976
rect 120834 151936 120874 151976
rect 120916 151936 120956 151976
rect 120998 151936 121038 151976
rect 121080 151936 121120 151976
rect 135872 151936 135912 151976
rect 135954 151936 135994 151976
rect 136036 151936 136076 151976
rect 136118 151936 136158 151976
rect 136200 151936 136240 151976
rect 150992 151936 151032 151976
rect 151074 151936 151114 151976
rect 151156 151936 151196 151976
rect 151238 151936 151278 151976
rect 151320 151936 151360 151976
rect 74152 151180 74192 151220
rect 74234 151180 74274 151220
rect 74316 151180 74356 151220
rect 74398 151180 74438 151220
rect 74480 151180 74520 151220
rect 89272 151180 89312 151220
rect 89354 151180 89394 151220
rect 89436 151180 89476 151220
rect 89518 151180 89558 151220
rect 89600 151180 89640 151220
rect 104392 151180 104432 151220
rect 104474 151180 104514 151220
rect 104556 151180 104596 151220
rect 104638 151180 104678 151220
rect 104720 151180 104760 151220
rect 119512 151180 119552 151220
rect 119594 151180 119634 151220
rect 119676 151180 119716 151220
rect 119758 151180 119798 151220
rect 119840 151180 119880 151220
rect 134632 151180 134672 151220
rect 134714 151180 134754 151220
rect 134796 151180 134836 151220
rect 134878 151180 134918 151220
rect 134960 151180 135000 151220
rect 149752 151180 149792 151220
rect 149834 151180 149874 151220
rect 149916 151180 149956 151220
rect 149998 151180 150038 151220
rect 150080 151180 150120 151220
rect 75392 150424 75432 150464
rect 75474 150424 75514 150464
rect 75556 150424 75596 150464
rect 75638 150424 75678 150464
rect 75720 150424 75760 150464
rect 90512 150424 90552 150464
rect 90594 150424 90634 150464
rect 90676 150424 90716 150464
rect 90758 150424 90798 150464
rect 90840 150424 90880 150464
rect 105632 150424 105672 150464
rect 105714 150424 105754 150464
rect 105796 150424 105836 150464
rect 105878 150424 105918 150464
rect 105960 150424 106000 150464
rect 120752 150424 120792 150464
rect 120834 150424 120874 150464
rect 120916 150424 120956 150464
rect 120998 150424 121038 150464
rect 121080 150424 121120 150464
rect 135872 150424 135912 150464
rect 135954 150424 135994 150464
rect 136036 150424 136076 150464
rect 136118 150424 136158 150464
rect 136200 150424 136240 150464
rect 150992 150424 151032 150464
rect 151074 150424 151114 150464
rect 151156 150424 151196 150464
rect 151238 150424 151278 150464
rect 151320 150424 151360 150464
rect 74152 149668 74192 149708
rect 74234 149668 74274 149708
rect 74316 149668 74356 149708
rect 74398 149668 74438 149708
rect 74480 149668 74520 149708
rect 89272 149668 89312 149708
rect 89354 149668 89394 149708
rect 89436 149668 89476 149708
rect 89518 149668 89558 149708
rect 89600 149668 89640 149708
rect 104392 149668 104432 149708
rect 104474 149668 104514 149708
rect 104556 149668 104596 149708
rect 104638 149668 104678 149708
rect 104720 149668 104760 149708
rect 119512 149668 119552 149708
rect 119594 149668 119634 149708
rect 119676 149668 119716 149708
rect 119758 149668 119798 149708
rect 119840 149668 119880 149708
rect 134632 149668 134672 149708
rect 134714 149668 134754 149708
rect 134796 149668 134836 149708
rect 134878 149668 134918 149708
rect 134960 149668 135000 149708
rect 149752 149668 149792 149708
rect 149834 149668 149874 149708
rect 149916 149668 149956 149708
rect 149998 149668 150038 149708
rect 150080 149668 150120 149708
rect 75392 148912 75432 148952
rect 75474 148912 75514 148952
rect 75556 148912 75596 148952
rect 75638 148912 75678 148952
rect 75720 148912 75760 148952
rect 90512 148912 90552 148952
rect 90594 148912 90634 148952
rect 90676 148912 90716 148952
rect 90758 148912 90798 148952
rect 90840 148912 90880 148952
rect 105632 148912 105672 148952
rect 105714 148912 105754 148952
rect 105796 148912 105836 148952
rect 105878 148912 105918 148952
rect 105960 148912 106000 148952
rect 120752 148912 120792 148952
rect 120834 148912 120874 148952
rect 120916 148912 120956 148952
rect 120998 148912 121038 148952
rect 121080 148912 121120 148952
rect 135872 148912 135912 148952
rect 135954 148912 135994 148952
rect 136036 148912 136076 148952
rect 136118 148912 136158 148952
rect 136200 148912 136240 148952
rect 150992 148912 151032 148952
rect 151074 148912 151114 148952
rect 151156 148912 151196 148952
rect 151238 148912 151278 148952
rect 151320 148912 151360 148952
rect 74152 148156 74192 148196
rect 74234 148156 74274 148196
rect 74316 148156 74356 148196
rect 74398 148156 74438 148196
rect 74480 148156 74520 148196
rect 89272 148156 89312 148196
rect 89354 148156 89394 148196
rect 89436 148156 89476 148196
rect 89518 148156 89558 148196
rect 89600 148156 89640 148196
rect 104392 148156 104432 148196
rect 104474 148156 104514 148196
rect 104556 148156 104596 148196
rect 104638 148156 104678 148196
rect 104720 148156 104760 148196
rect 119512 148156 119552 148196
rect 119594 148156 119634 148196
rect 119676 148156 119716 148196
rect 119758 148156 119798 148196
rect 119840 148156 119880 148196
rect 134632 148156 134672 148196
rect 134714 148156 134754 148196
rect 134796 148156 134836 148196
rect 134878 148156 134918 148196
rect 134960 148156 135000 148196
rect 149752 148156 149792 148196
rect 149834 148156 149874 148196
rect 149916 148156 149956 148196
rect 149998 148156 150038 148196
rect 150080 148156 150120 148196
rect 75392 147400 75432 147440
rect 75474 147400 75514 147440
rect 75556 147400 75596 147440
rect 75638 147400 75678 147440
rect 75720 147400 75760 147440
rect 90512 147400 90552 147440
rect 90594 147400 90634 147440
rect 90676 147400 90716 147440
rect 90758 147400 90798 147440
rect 90840 147400 90880 147440
rect 105632 147400 105672 147440
rect 105714 147400 105754 147440
rect 105796 147400 105836 147440
rect 105878 147400 105918 147440
rect 105960 147400 106000 147440
rect 120752 147400 120792 147440
rect 120834 147400 120874 147440
rect 120916 147400 120956 147440
rect 120998 147400 121038 147440
rect 121080 147400 121120 147440
rect 135872 147400 135912 147440
rect 135954 147400 135994 147440
rect 136036 147400 136076 147440
rect 136118 147400 136158 147440
rect 136200 147400 136240 147440
rect 150992 147400 151032 147440
rect 151074 147400 151114 147440
rect 151156 147400 151196 147440
rect 151238 147400 151278 147440
rect 151320 147400 151360 147440
rect 74152 146644 74192 146684
rect 74234 146644 74274 146684
rect 74316 146644 74356 146684
rect 74398 146644 74438 146684
rect 74480 146644 74520 146684
rect 89272 146644 89312 146684
rect 89354 146644 89394 146684
rect 89436 146644 89476 146684
rect 89518 146644 89558 146684
rect 89600 146644 89640 146684
rect 104392 146644 104432 146684
rect 104474 146644 104514 146684
rect 104556 146644 104596 146684
rect 104638 146644 104678 146684
rect 104720 146644 104760 146684
rect 119512 146644 119552 146684
rect 119594 146644 119634 146684
rect 119676 146644 119716 146684
rect 119758 146644 119798 146684
rect 119840 146644 119880 146684
rect 134632 146644 134672 146684
rect 134714 146644 134754 146684
rect 134796 146644 134836 146684
rect 134878 146644 134918 146684
rect 134960 146644 135000 146684
rect 149752 146644 149792 146684
rect 149834 146644 149874 146684
rect 149916 146644 149956 146684
rect 149998 146644 150038 146684
rect 150080 146644 150120 146684
rect 75392 145888 75432 145928
rect 75474 145888 75514 145928
rect 75556 145888 75596 145928
rect 75638 145888 75678 145928
rect 75720 145888 75760 145928
rect 90512 145888 90552 145928
rect 90594 145888 90634 145928
rect 90676 145888 90716 145928
rect 90758 145888 90798 145928
rect 90840 145888 90880 145928
rect 105632 145888 105672 145928
rect 105714 145888 105754 145928
rect 105796 145888 105836 145928
rect 105878 145888 105918 145928
rect 105960 145888 106000 145928
rect 120752 145888 120792 145928
rect 120834 145888 120874 145928
rect 120916 145888 120956 145928
rect 120998 145888 121038 145928
rect 121080 145888 121120 145928
rect 135872 145888 135912 145928
rect 135954 145888 135994 145928
rect 136036 145888 136076 145928
rect 136118 145888 136158 145928
rect 136200 145888 136240 145928
rect 150992 145888 151032 145928
rect 151074 145888 151114 145928
rect 151156 145888 151196 145928
rect 151238 145888 151278 145928
rect 151320 145888 151360 145928
rect 74152 145132 74192 145172
rect 74234 145132 74274 145172
rect 74316 145132 74356 145172
rect 74398 145132 74438 145172
rect 74480 145132 74520 145172
rect 89272 145132 89312 145172
rect 89354 145132 89394 145172
rect 89436 145132 89476 145172
rect 89518 145132 89558 145172
rect 89600 145132 89640 145172
rect 104392 145132 104432 145172
rect 104474 145132 104514 145172
rect 104556 145132 104596 145172
rect 104638 145132 104678 145172
rect 104720 145132 104760 145172
rect 119512 145132 119552 145172
rect 119594 145132 119634 145172
rect 119676 145132 119716 145172
rect 119758 145132 119798 145172
rect 119840 145132 119880 145172
rect 134632 145132 134672 145172
rect 134714 145132 134754 145172
rect 134796 145132 134836 145172
rect 134878 145132 134918 145172
rect 134960 145132 135000 145172
rect 149752 145132 149792 145172
rect 149834 145132 149874 145172
rect 149916 145132 149956 145172
rect 149998 145132 150038 145172
rect 150080 145132 150120 145172
rect 75392 144376 75432 144416
rect 75474 144376 75514 144416
rect 75556 144376 75596 144416
rect 75638 144376 75678 144416
rect 75720 144376 75760 144416
rect 90512 144376 90552 144416
rect 90594 144376 90634 144416
rect 90676 144376 90716 144416
rect 90758 144376 90798 144416
rect 90840 144376 90880 144416
rect 105632 144376 105672 144416
rect 105714 144376 105754 144416
rect 105796 144376 105836 144416
rect 105878 144376 105918 144416
rect 105960 144376 106000 144416
rect 120752 144376 120792 144416
rect 120834 144376 120874 144416
rect 120916 144376 120956 144416
rect 120998 144376 121038 144416
rect 121080 144376 121120 144416
rect 135872 144376 135912 144416
rect 135954 144376 135994 144416
rect 136036 144376 136076 144416
rect 136118 144376 136158 144416
rect 136200 144376 136240 144416
rect 150992 144376 151032 144416
rect 151074 144376 151114 144416
rect 151156 144376 151196 144416
rect 151238 144376 151278 144416
rect 151320 144376 151360 144416
rect 74152 143620 74192 143660
rect 74234 143620 74274 143660
rect 74316 143620 74356 143660
rect 74398 143620 74438 143660
rect 74480 143620 74520 143660
rect 89272 143620 89312 143660
rect 89354 143620 89394 143660
rect 89436 143620 89476 143660
rect 89518 143620 89558 143660
rect 89600 143620 89640 143660
rect 104392 143620 104432 143660
rect 104474 143620 104514 143660
rect 104556 143620 104596 143660
rect 104638 143620 104678 143660
rect 104720 143620 104760 143660
rect 119512 143620 119552 143660
rect 119594 143620 119634 143660
rect 119676 143620 119716 143660
rect 119758 143620 119798 143660
rect 119840 143620 119880 143660
rect 134632 143620 134672 143660
rect 134714 143620 134754 143660
rect 134796 143620 134836 143660
rect 134878 143620 134918 143660
rect 134960 143620 135000 143660
rect 149752 143620 149792 143660
rect 149834 143620 149874 143660
rect 149916 143620 149956 143660
rect 149998 143620 150038 143660
rect 150080 143620 150120 143660
rect 75392 142864 75432 142904
rect 75474 142864 75514 142904
rect 75556 142864 75596 142904
rect 75638 142864 75678 142904
rect 75720 142864 75760 142904
rect 90512 142864 90552 142904
rect 90594 142864 90634 142904
rect 90676 142864 90716 142904
rect 90758 142864 90798 142904
rect 90840 142864 90880 142904
rect 105632 142864 105672 142904
rect 105714 142864 105754 142904
rect 105796 142864 105836 142904
rect 105878 142864 105918 142904
rect 105960 142864 106000 142904
rect 120752 142864 120792 142904
rect 120834 142864 120874 142904
rect 120916 142864 120956 142904
rect 120998 142864 121038 142904
rect 121080 142864 121120 142904
rect 135872 142864 135912 142904
rect 135954 142864 135994 142904
rect 136036 142864 136076 142904
rect 136118 142864 136158 142904
rect 136200 142864 136240 142904
rect 150992 142864 151032 142904
rect 151074 142864 151114 142904
rect 151156 142864 151196 142904
rect 151238 142864 151278 142904
rect 151320 142864 151360 142904
rect 74152 142108 74192 142148
rect 74234 142108 74274 142148
rect 74316 142108 74356 142148
rect 74398 142108 74438 142148
rect 74480 142108 74520 142148
rect 89272 142108 89312 142148
rect 89354 142108 89394 142148
rect 89436 142108 89476 142148
rect 89518 142108 89558 142148
rect 89600 142108 89640 142148
rect 104392 142108 104432 142148
rect 104474 142108 104514 142148
rect 104556 142108 104596 142148
rect 104638 142108 104678 142148
rect 104720 142108 104760 142148
rect 119512 142108 119552 142148
rect 119594 142108 119634 142148
rect 119676 142108 119716 142148
rect 119758 142108 119798 142148
rect 119840 142108 119880 142148
rect 134632 142108 134672 142148
rect 134714 142108 134754 142148
rect 134796 142108 134836 142148
rect 134878 142108 134918 142148
rect 134960 142108 135000 142148
rect 149752 142108 149792 142148
rect 149834 142108 149874 142148
rect 149916 142108 149956 142148
rect 149998 142108 150038 142148
rect 150080 142108 150120 142148
rect 75392 141352 75432 141392
rect 75474 141352 75514 141392
rect 75556 141352 75596 141392
rect 75638 141352 75678 141392
rect 75720 141352 75760 141392
rect 90512 141352 90552 141392
rect 90594 141352 90634 141392
rect 90676 141352 90716 141392
rect 90758 141352 90798 141392
rect 90840 141352 90880 141392
rect 105632 141352 105672 141392
rect 105714 141352 105754 141392
rect 105796 141352 105836 141392
rect 105878 141352 105918 141392
rect 105960 141352 106000 141392
rect 120752 141352 120792 141392
rect 120834 141352 120874 141392
rect 120916 141352 120956 141392
rect 120998 141352 121038 141392
rect 121080 141352 121120 141392
rect 135872 141352 135912 141392
rect 135954 141352 135994 141392
rect 136036 141352 136076 141392
rect 136118 141352 136158 141392
rect 136200 141352 136240 141392
rect 150992 141352 151032 141392
rect 151074 141352 151114 141392
rect 151156 141352 151196 141392
rect 151238 141352 151278 141392
rect 151320 141352 151360 141392
rect 74152 140596 74192 140636
rect 74234 140596 74274 140636
rect 74316 140596 74356 140636
rect 74398 140596 74438 140636
rect 74480 140596 74520 140636
rect 89272 140596 89312 140636
rect 89354 140596 89394 140636
rect 89436 140596 89476 140636
rect 89518 140596 89558 140636
rect 89600 140596 89640 140636
rect 104392 140596 104432 140636
rect 104474 140596 104514 140636
rect 104556 140596 104596 140636
rect 104638 140596 104678 140636
rect 104720 140596 104760 140636
rect 119512 140596 119552 140636
rect 119594 140596 119634 140636
rect 119676 140596 119716 140636
rect 119758 140596 119798 140636
rect 119840 140596 119880 140636
rect 134632 140596 134672 140636
rect 134714 140596 134754 140636
rect 134796 140596 134836 140636
rect 134878 140596 134918 140636
rect 134960 140596 135000 140636
rect 149752 140596 149792 140636
rect 149834 140596 149874 140636
rect 149916 140596 149956 140636
rect 149998 140596 150038 140636
rect 150080 140596 150120 140636
rect 75392 139840 75432 139880
rect 75474 139840 75514 139880
rect 75556 139840 75596 139880
rect 75638 139840 75678 139880
rect 75720 139840 75760 139880
rect 90512 139840 90552 139880
rect 90594 139840 90634 139880
rect 90676 139840 90716 139880
rect 90758 139840 90798 139880
rect 90840 139840 90880 139880
rect 105632 139840 105672 139880
rect 105714 139840 105754 139880
rect 105796 139840 105836 139880
rect 105878 139840 105918 139880
rect 105960 139840 106000 139880
rect 120752 139840 120792 139880
rect 120834 139840 120874 139880
rect 120916 139840 120956 139880
rect 120998 139840 121038 139880
rect 121080 139840 121120 139880
rect 135872 139840 135912 139880
rect 135954 139840 135994 139880
rect 136036 139840 136076 139880
rect 136118 139840 136158 139880
rect 136200 139840 136240 139880
rect 150992 139840 151032 139880
rect 151074 139840 151114 139880
rect 151156 139840 151196 139880
rect 151238 139840 151278 139880
rect 151320 139840 151360 139880
rect 74152 139084 74192 139124
rect 74234 139084 74274 139124
rect 74316 139084 74356 139124
rect 74398 139084 74438 139124
rect 74480 139084 74520 139124
rect 89272 139084 89312 139124
rect 89354 139084 89394 139124
rect 89436 139084 89476 139124
rect 89518 139084 89558 139124
rect 89600 139084 89640 139124
rect 104392 139084 104432 139124
rect 104474 139084 104514 139124
rect 104556 139084 104596 139124
rect 104638 139084 104678 139124
rect 104720 139084 104760 139124
rect 119512 139084 119552 139124
rect 119594 139084 119634 139124
rect 119676 139084 119716 139124
rect 119758 139084 119798 139124
rect 119840 139084 119880 139124
rect 134632 139084 134672 139124
rect 134714 139084 134754 139124
rect 134796 139084 134836 139124
rect 134878 139084 134918 139124
rect 134960 139084 135000 139124
rect 149752 139084 149792 139124
rect 149834 139084 149874 139124
rect 149916 139084 149956 139124
rect 149998 139084 150038 139124
rect 150080 139084 150120 139124
rect 75392 138328 75432 138368
rect 75474 138328 75514 138368
rect 75556 138328 75596 138368
rect 75638 138328 75678 138368
rect 75720 138328 75760 138368
rect 90512 138328 90552 138368
rect 90594 138328 90634 138368
rect 90676 138328 90716 138368
rect 90758 138328 90798 138368
rect 90840 138328 90880 138368
rect 105632 138328 105672 138368
rect 105714 138328 105754 138368
rect 105796 138328 105836 138368
rect 105878 138328 105918 138368
rect 105960 138328 106000 138368
rect 120752 138328 120792 138368
rect 120834 138328 120874 138368
rect 120916 138328 120956 138368
rect 120998 138328 121038 138368
rect 121080 138328 121120 138368
rect 135872 138328 135912 138368
rect 135954 138328 135994 138368
rect 136036 138328 136076 138368
rect 136118 138328 136158 138368
rect 136200 138328 136240 138368
rect 150992 138328 151032 138368
rect 151074 138328 151114 138368
rect 151156 138328 151196 138368
rect 151238 138328 151278 138368
rect 151320 138328 151360 138368
rect 74152 137572 74192 137612
rect 74234 137572 74274 137612
rect 74316 137572 74356 137612
rect 74398 137572 74438 137612
rect 74480 137572 74520 137612
rect 89272 137572 89312 137612
rect 89354 137572 89394 137612
rect 89436 137572 89476 137612
rect 89518 137572 89558 137612
rect 89600 137572 89640 137612
rect 104392 137572 104432 137612
rect 104474 137572 104514 137612
rect 104556 137572 104596 137612
rect 104638 137572 104678 137612
rect 104720 137572 104760 137612
rect 119512 137572 119552 137612
rect 119594 137572 119634 137612
rect 119676 137572 119716 137612
rect 119758 137572 119798 137612
rect 119840 137572 119880 137612
rect 134632 137572 134672 137612
rect 134714 137572 134754 137612
rect 134796 137572 134836 137612
rect 134878 137572 134918 137612
rect 134960 137572 135000 137612
rect 149752 137572 149792 137612
rect 149834 137572 149874 137612
rect 149916 137572 149956 137612
rect 149998 137572 150038 137612
rect 150080 137572 150120 137612
rect 75392 136816 75432 136856
rect 75474 136816 75514 136856
rect 75556 136816 75596 136856
rect 75638 136816 75678 136856
rect 75720 136816 75760 136856
rect 90512 136816 90552 136856
rect 90594 136816 90634 136856
rect 90676 136816 90716 136856
rect 90758 136816 90798 136856
rect 90840 136816 90880 136856
rect 105632 136816 105672 136856
rect 105714 136816 105754 136856
rect 105796 136816 105836 136856
rect 105878 136816 105918 136856
rect 105960 136816 106000 136856
rect 120752 136816 120792 136856
rect 120834 136816 120874 136856
rect 120916 136816 120956 136856
rect 120998 136816 121038 136856
rect 121080 136816 121120 136856
rect 135872 136816 135912 136856
rect 135954 136816 135994 136856
rect 136036 136816 136076 136856
rect 136118 136816 136158 136856
rect 136200 136816 136240 136856
rect 150992 136816 151032 136856
rect 151074 136816 151114 136856
rect 151156 136816 151196 136856
rect 151238 136816 151278 136856
rect 151320 136816 151360 136856
rect 74152 136060 74192 136100
rect 74234 136060 74274 136100
rect 74316 136060 74356 136100
rect 74398 136060 74438 136100
rect 74480 136060 74520 136100
rect 89272 136060 89312 136100
rect 89354 136060 89394 136100
rect 89436 136060 89476 136100
rect 89518 136060 89558 136100
rect 89600 136060 89640 136100
rect 104392 136060 104432 136100
rect 104474 136060 104514 136100
rect 104556 136060 104596 136100
rect 104638 136060 104678 136100
rect 104720 136060 104760 136100
rect 119512 136060 119552 136100
rect 119594 136060 119634 136100
rect 119676 136060 119716 136100
rect 119758 136060 119798 136100
rect 119840 136060 119880 136100
rect 134632 136060 134672 136100
rect 134714 136060 134754 136100
rect 134796 136060 134836 136100
rect 134878 136060 134918 136100
rect 134960 136060 135000 136100
rect 149752 136060 149792 136100
rect 149834 136060 149874 136100
rect 149916 136060 149956 136100
rect 149998 136060 150038 136100
rect 150080 136060 150120 136100
rect 75392 135304 75432 135344
rect 75474 135304 75514 135344
rect 75556 135304 75596 135344
rect 75638 135304 75678 135344
rect 75720 135304 75760 135344
rect 90512 135304 90552 135344
rect 90594 135304 90634 135344
rect 90676 135304 90716 135344
rect 90758 135304 90798 135344
rect 90840 135304 90880 135344
rect 105632 135304 105672 135344
rect 105714 135304 105754 135344
rect 105796 135304 105836 135344
rect 105878 135304 105918 135344
rect 105960 135304 106000 135344
rect 120752 135304 120792 135344
rect 120834 135304 120874 135344
rect 120916 135304 120956 135344
rect 120998 135304 121038 135344
rect 121080 135304 121120 135344
rect 135872 135304 135912 135344
rect 135954 135304 135994 135344
rect 136036 135304 136076 135344
rect 136118 135304 136158 135344
rect 136200 135304 136240 135344
rect 150992 135304 151032 135344
rect 151074 135304 151114 135344
rect 151156 135304 151196 135344
rect 151238 135304 151278 135344
rect 151320 135304 151360 135344
rect 74152 134548 74192 134588
rect 74234 134548 74274 134588
rect 74316 134548 74356 134588
rect 74398 134548 74438 134588
rect 74480 134548 74520 134588
rect 89272 134548 89312 134588
rect 89354 134548 89394 134588
rect 89436 134548 89476 134588
rect 89518 134548 89558 134588
rect 89600 134548 89640 134588
rect 104392 134548 104432 134588
rect 104474 134548 104514 134588
rect 104556 134548 104596 134588
rect 104638 134548 104678 134588
rect 104720 134548 104760 134588
rect 119512 134548 119552 134588
rect 119594 134548 119634 134588
rect 119676 134548 119716 134588
rect 119758 134548 119798 134588
rect 119840 134548 119880 134588
rect 134632 134548 134672 134588
rect 134714 134548 134754 134588
rect 134796 134548 134836 134588
rect 134878 134548 134918 134588
rect 134960 134548 135000 134588
rect 149752 134548 149792 134588
rect 149834 134548 149874 134588
rect 149916 134548 149956 134588
rect 149998 134548 150038 134588
rect 150080 134548 150120 134588
rect 75392 133792 75432 133832
rect 75474 133792 75514 133832
rect 75556 133792 75596 133832
rect 75638 133792 75678 133832
rect 75720 133792 75760 133832
rect 90512 133792 90552 133832
rect 90594 133792 90634 133832
rect 90676 133792 90716 133832
rect 90758 133792 90798 133832
rect 90840 133792 90880 133832
rect 105632 133792 105672 133832
rect 105714 133792 105754 133832
rect 105796 133792 105836 133832
rect 105878 133792 105918 133832
rect 105960 133792 106000 133832
rect 120752 133792 120792 133832
rect 120834 133792 120874 133832
rect 120916 133792 120956 133832
rect 120998 133792 121038 133832
rect 121080 133792 121120 133832
rect 135872 133792 135912 133832
rect 135954 133792 135994 133832
rect 136036 133792 136076 133832
rect 136118 133792 136158 133832
rect 136200 133792 136240 133832
rect 150992 133792 151032 133832
rect 151074 133792 151114 133832
rect 151156 133792 151196 133832
rect 151238 133792 151278 133832
rect 151320 133792 151360 133832
rect 74152 133036 74192 133076
rect 74234 133036 74274 133076
rect 74316 133036 74356 133076
rect 74398 133036 74438 133076
rect 74480 133036 74520 133076
rect 89272 133036 89312 133076
rect 89354 133036 89394 133076
rect 89436 133036 89476 133076
rect 89518 133036 89558 133076
rect 89600 133036 89640 133076
rect 104392 133036 104432 133076
rect 104474 133036 104514 133076
rect 104556 133036 104596 133076
rect 104638 133036 104678 133076
rect 104720 133036 104760 133076
rect 119512 133036 119552 133076
rect 119594 133036 119634 133076
rect 119676 133036 119716 133076
rect 119758 133036 119798 133076
rect 119840 133036 119880 133076
rect 134632 133036 134672 133076
rect 134714 133036 134754 133076
rect 134796 133036 134836 133076
rect 134878 133036 134918 133076
rect 134960 133036 135000 133076
rect 149752 133036 149792 133076
rect 149834 133036 149874 133076
rect 149916 133036 149956 133076
rect 149998 133036 150038 133076
rect 150080 133036 150120 133076
rect 75392 132280 75432 132320
rect 75474 132280 75514 132320
rect 75556 132280 75596 132320
rect 75638 132280 75678 132320
rect 75720 132280 75760 132320
rect 90512 132280 90552 132320
rect 90594 132280 90634 132320
rect 90676 132280 90716 132320
rect 90758 132280 90798 132320
rect 90840 132280 90880 132320
rect 105632 132280 105672 132320
rect 105714 132280 105754 132320
rect 105796 132280 105836 132320
rect 105878 132280 105918 132320
rect 105960 132280 106000 132320
rect 120752 132280 120792 132320
rect 120834 132280 120874 132320
rect 120916 132280 120956 132320
rect 120998 132280 121038 132320
rect 121080 132280 121120 132320
rect 135872 132280 135912 132320
rect 135954 132280 135994 132320
rect 136036 132280 136076 132320
rect 136118 132280 136158 132320
rect 136200 132280 136240 132320
rect 150992 132280 151032 132320
rect 151074 132280 151114 132320
rect 151156 132280 151196 132320
rect 151238 132280 151278 132320
rect 151320 132280 151360 132320
rect 74152 131524 74192 131564
rect 74234 131524 74274 131564
rect 74316 131524 74356 131564
rect 74398 131524 74438 131564
rect 74480 131524 74520 131564
rect 89272 131524 89312 131564
rect 89354 131524 89394 131564
rect 89436 131524 89476 131564
rect 89518 131524 89558 131564
rect 89600 131524 89640 131564
rect 104392 131524 104432 131564
rect 104474 131524 104514 131564
rect 104556 131524 104596 131564
rect 104638 131524 104678 131564
rect 104720 131524 104760 131564
rect 119512 131524 119552 131564
rect 119594 131524 119634 131564
rect 119676 131524 119716 131564
rect 119758 131524 119798 131564
rect 119840 131524 119880 131564
rect 134632 131524 134672 131564
rect 134714 131524 134754 131564
rect 134796 131524 134836 131564
rect 134878 131524 134918 131564
rect 134960 131524 135000 131564
rect 149752 131524 149792 131564
rect 149834 131524 149874 131564
rect 149916 131524 149956 131564
rect 149998 131524 150038 131564
rect 150080 131524 150120 131564
rect 75392 130768 75432 130808
rect 75474 130768 75514 130808
rect 75556 130768 75596 130808
rect 75638 130768 75678 130808
rect 75720 130768 75760 130808
rect 90512 130768 90552 130808
rect 90594 130768 90634 130808
rect 90676 130768 90716 130808
rect 90758 130768 90798 130808
rect 90840 130768 90880 130808
rect 105632 130768 105672 130808
rect 105714 130768 105754 130808
rect 105796 130768 105836 130808
rect 105878 130768 105918 130808
rect 105960 130768 106000 130808
rect 120752 130768 120792 130808
rect 120834 130768 120874 130808
rect 120916 130768 120956 130808
rect 120998 130768 121038 130808
rect 121080 130768 121120 130808
rect 135872 130768 135912 130808
rect 135954 130768 135994 130808
rect 136036 130768 136076 130808
rect 136118 130768 136158 130808
rect 136200 130768 136240 130808
rect 150992 130768 151032 130808
rect 151074 130768 151114 130808
rect 151156 130768 151196 130808
rect 151238 130768 151278 130808
rect 151320 130768 151360 130808
rect 74152 130012 74192 130052
rect 74234 130012 74274 130052
rect 74316 130012 74356 130052
rect 74398 130012 74438 130052
rect 74480 130012 74520 130052
rect 89272 130012 89312 130052
rect 89354 130012 89394 130052
rect 89436 130012 89476 130052
rect 89518 130012 89558 130052
rect 89600 130012 89640 130052
rect 104392 130012 104432 130052
rect 104474 130012 104514 130052
rect 104556 130012 104596 130052
rect 104638 130012 104678 130052
rect 104720 130012 104760 130052
rect 119512 130012 119552 130052
rect 119594 130012 119634 130052
rect 119676 130012 119716 130052
rect 119758 130012 119798 130052
rect 119840 130012 119880 130052
rect 134632 130012 134672 130052
rect 134714 130012 134754 130052
rect 134796 130012 134836 130052
rect 134878 130012 134918 130052
rect 134960 130012 135000 130052
rect 149752 130012 149792 130052
rect 149834 130012 149874 130052
rect 149916 130012 149956 130052
rect 149998 130012 150038 130052
rect 150080 130012 150120 130052
rect 75392 129256 75432 129296
rect 75474 129256 75514 129296
rect 75556 129256 75596 129296
rect 75638 129256 75678 129296
rect 75720 129256 75760 129296
rect 90512 129256 90552 129296
rect 90594 129256 90634 129296
rect 90676 129256 90716 129296
rect 90758 129256 90798 129296
rect 90840 129256 90880 129296
rect 105632 129256 105672 129296
rect 105714 129256 105754 129296
rect 105796 129256 105836 129296
rect 105878 129256 105918 129296
rect 105960 129256 106000 129296
rect 120752 129256 120792 129296
rect 120834 129256 120874 129296
rect 120916 129256 120956 129296
rect 120998 129256 121038 129296
rect 121080 129256 121120 129296
rect 135872 129256 135912 129296
rect 135954 129256 135994 129296
rect 136036 129256 136076 129296
rect 136118 129256 136158 129296
rect 136200 129256 136240 129296
rect 150992 129256 151032 129296
rect 151074 129256 151114 129296
rect 151156 129256 151196 129296
rect 151238 129256 151278 129296
rect 151320 129256 151360 129296
rect 74152 128500 74192 128540
rect 74234 128500 74274 128540
rect 74316 128500 74356 128540
rect 74398 128500 74438 128540
rect 74480 128500 74520 128540
rect 89272 128500 89312 128540
rect 89354 128500 89394 128540
rect 89436 128500 89476 128540
rect 89518 128500 89558 128540
rect 89600 128500 89640 128540
rect 104392 128500 104432 128540
rect 104474 128500 104514 128540
rect 104556 128500 104596 128540
rect 104638 128500 104678 128540
rect 104720 128500 104760 128540
rect 119512 128500 119552 128540
rect 119594 128500 119634 128540
rect 119676 128500 119716 128540
rect 119758 128500 119798 128540
rect 119840 128500 119880 128540
rect 134632 128500 134672 128540
rect 134714 128500 134754 128540
rect 134796 128500 134836 128540
rect 134878 128500 134918 128540
rect 134960 128500 135000 128540
rect 149752 128500 149792 128540
rect 149834 128500 149874 128540
rect 149916 128500 149956 128540
rect 149998 128500 150038 128540
rect 150080 128500 150120 128540
rect 75392 127744 75432 127784
rect 75474 127744 75514 127784
rect 75556 127744 75596 127784
rect 75638 127744 75678 127784
rect 75720 127744 75760 127784
rect 90512 127744 90552 127784
rect 90594 127744 90634 127784
rect 90676 127744 90716 127784
rect 90758 127744 90798 127784
rect 90840 127744 90880 127784
rect 105632 127744 105672 127784
rect 105714 127744 105754 127784
rect 105796 127744 105836 127784
rect 105878 127744 105918 127784
rect 105960 127744 106000 127784
rect 120752 127744 120792 127784
rect 120834 127744 120874 127784
rect 120916 127744 120956 127784
rect 120998 127744 121038 127784
rect 121080 127744 121120 127784
rect 135872 127744 135912 127784
rect 135954 127744 135994 127784
rect 136036 127744 136076 127784
rect 136118 127744 136158 127784
rect 136200 127744 136240 127784
rect 150992 127744 151032 127784
rect 151074 127744 151114 127784
rect 151156 127744 151196 127784
rect 151238 127744 151278 127784
rect 151320 127744 151360 127784
rect 74152 126988 74192 127028
rect 74234 126988 74274 127028
rect 74316 126988 74356 127028
rect 74398 126988 74438 127028
rect 74480 126988 74520 127028
rect 89272 126988 89312 127028
rect 89354 126988 89394 127028
rect 89436 126988 89476 127028
rect 89518 126988 89558 127028
rect 89600 126988 89640 127028
rect 104392 126988 104432 127028
rect 104474 126988 104514 127028
rect 104556 126988 104596 127028
rect 104638 126988 104678 127028
rect 104720 126988 104760 127028
rect 119512 126988 119552 127028
rect 119594 126988 119634 127028
rect 119676 126988 119716 127028
rect 119758 126988 119798 127028
rect 119840 126988 119880 127028
rect 134632 126988 134672 127028
rect 134714 126988 134754 127028
rect 134796 126988 134836 127028
rect 134878 126988 134918 127028
rect 134960 126988 135000 127028
rect 149752 126988 149792 127028
rect 149834 126988 149874 127028
rect 149916 126988 149956 127028
rect 149998 126988 150038 127028
rect 150080 126988 150120 127028
rect 75392 126232 75432 126272
rect 75474 126232 75514 126272
rect 75556 126232 75596 126272
rect 75638 126232 75678 126272
rect 75720 126232 75760 126272
rect 90512 126232 90552 126272
rect 90594 126232 90634 126272
rect 90676 126232 90716 126272
rect 90758 126232 90798 126272
rect 90840 126232 90880 126272
rect 105632 126232 105672 126272
rect 105714 126232 105754 126272
rect 105796 126232 105836 126272
rect 105878 126232 105918 126272
rect 105960 126232 106000 126272
rect 120752 126232 120792 126272
rect 120834 126232 120874 126272
rect 120916 126232 120956 126272
rect 120998 126232 121038 126272
rect 121080 126232 121120 126272
rect 135872 126232 135912 126272
rect 135954 126232 135994 126272
rect 136036 126232 136076 126272
rect 136118 126232 136158 126272
rect 136200 126232 136240 126272
rect 150992 126232 151032 126272
rect 151074 126232 151114 126272
rect 151156 126232 151196 126272
rect 151238 126232 151278 126272
rect 151320 126232 151360 126272
rect 74152 125476 74192 125516
rect 74234 125476 74274 125516
rect 74316 125476 74356 125516
rect 74398 125476 74438 125516
rect 74480 125476 74520 125516
rect 89272 125476 89312 125516
rect 89354 125476 89394 125516
rect 89436 125476 89476 125516
rect 89518 125476 89558 125516
rect 89600 125476 89640 125516
rect 104392 125476 104432 125516
rect 104474 125476 104514 125516
rect 104556 125476 104596 125516
rect 104638 125476 104678 125516
rect 104720 125476 104760 125516
rect 119512 125476 119552 125516
rect 119594 125476 119634 125516
rect 119676 125476 119716 125516
rect 119758 125476 119798 125516
rect 119840 125476 119880 125516
rect 134632 125476 134672 125516
rect 134714 125476 134754 125516
rect 134796 125476 134836 125516
rect 134878 125476 134918 125516
rect 134960 125476 135000 125516
rect 149752 125476 149792 125516
rect 149834 125476 149874 125516
rect 149916 125476 149956 125516
rect 149998 125476 150038 125516
rect 150080 125476 150120 125516
rect 75392 124720 75432 124760
rect 75474 124720 75514 124760
rect 75556 124720 75596 124760
rect 75638 124720 75678 124760
rect 75720 124720 75760 124760
rect 90512 124720 90552 124760
rect 90594 124720 90634 124760
rect 90676 124720 90716 124760
rect 90758 124720 90798 124760
rect 90840 124720 90880 124760
rect 105632 124720 105672 124760
rect 105714 124720 105754 124760
rect 105796 124720 105836 124760
rect 105878 124720 105918 124760
rect 105960 124720 106000 124760
rect 120752 124720 120792 124760
rect 120834 124720 120874 124760
rect 120916 124720 120956 124760
rect 120998 124720 121038 124760
rect 121080 124720 121120 124760
rect 135872 124720 135912 124760
rect 135954 124720 135994 124760
rect 136036 124720 136076 124760
rect 136118 124720 136158 124760
rect 136200 124720 136240 124760
rect 150992 124720 151032 124760
rect 151074 124720 151114 124760
rect 151156 124720 151196 124760
rect 151238 124720 151278 124760
rect 151320 124720 151360 124760
rect 74152 123964 74192 124004
rect 74234 123964 74274 124004
rect 74316 123964 74356 124004
rect 74398 123964 74438 124004
rect 74480 123964 74520 124004
rect 89272 123964 89312 124004
rect 89354 123964 89394 124004
rect 89436 123964 89476 124004
rect 89518 123964 89558 124004
rect 89600 123964 89640 124004
rect 104392 123964 104432 124004
rect 104474 123964 104514 124004
rect 104556 123964 104596 124004
rect 104638 123964 104678 124004
rect 104720 123964 104760 124004
rect 119512 123964 119552 124004
rect 119594 123964 119634 124004
rect 119676 123964 119716 124004
rect 119758 123964 119798 124004
rect 119840 123964 119880 124004
rect 134632 123964 134672 124004
rect 134714 123964 134754 124004
rect 134796 123964 134836 124004
rect 134878 123964 134918 124004
rect 134960 123964 135000 124004
rect 149752 123964 149792 124004
rect 149834 123964 149874 124004
rect 149916 123964 149956 124004
rect 149998 123964 150038 124004
rect 150080 123964 150120 124004
rect 75392 123208 75432 123248
rect 75474 123208 75514 123248
rect 75556 123208 75596 123248
rect 75638 123208 75678 123248
rect 75720 123208 75760 123248
rect 90512 123208 90552 123248
rect 90594 123208 90634 123248
rect 90676 123208 90716 123248
rect 90758 123208 90798 123248
rect 90840 123208 90880 123248
rect 105632 123208 105672 123248
rect 105714 123208 105754 123248
rect 105796 123208 105836 123248
rect 105878 123208 105918 123248
rect 105960 123208 106000 123248
rect 120752 123208 120792 123248
rect 120834 123208 120874 123248
rect 120916 123208 120956 123248
rect 120998 123208 121038 123248
rect 121080 123208 121120 123248
rect 135872 123208 135912 123248
rect 135954 123208 135994 123248
rect 136036 123208 136076 123248
rect 136118 123208 136158 123248
rect 136200 123208 136240 123248
rect 150992 123208 151032 123248
rect 151074 123208 151114 123248
rect 151156 123208 151196 123248
rect 151238 123208 151278 123248
rect 151320 123208 151360 123248
rect 74152 122452 74192 122492
rect 74234 122452 74274 122492
rect 74316 122452 74356 122492
rect 74398 122452 74438 122492
rect 74480 122452 74520 122492
rect 89272 122452 89312 122492
rect 89354 122452 89394 122492
rect 89436 122452 89476 122492
rect 89518 122452 89558 122492
rect 89600 122452 89640 122492
rect 104392 122452 104432 122492
rect 104474 122452 104514 122492
rect 104556 122452 104596 122492
rect 104638 122452 104678 122492
rect 104720 122452 104760 122492
rect 119512 122452 119552 122492
rect 119594 122452 119634 122492
rect 119676 122452 119716 122492
rect 119758 122452 119798 122492
rect 119840 122452 119880 122492
rect 134632 122452 134672 122492
rect 134714 122452 134754 122492
rect 134796 122452 134836 122492
rect 134878 122452 134918 122492
rect 134960 122452 135000 122492
rect 149752 122452 149792 122492
rect 149834 122452 149874 122492
rect 149916 122452 149956 122492
rect 149998 122452 150038 122492
rect 150080 122452 150120 122492
rect 75392 121696 75432 121736
rect 75474 121696 75514 121736
rect 75556 121696 75596 121736
rect 75638 121696 75678 121736
rect 75720 121696 75760 121736
rect 90512 121696 90552 121736
rect 90594 121696 90634 121736
rect 90676 121696 90716 121736
rect 90758 121696 90798 121736
rect 90840 121696 90880 121736
rect 105632 121696 105672 121736
rect 105714 121696 105754 121736
rect 105796 121696 105836 121736
rect 105878 121696 105918 121736
rect 105960 121696 106000 121736
rect 120752 121696 120792 121736
rect 120834 121696 120874 121736
rect 120916 121696 120956 121736
rect 120998 121696 121038 121736
rect 121080 121696 121120 121736
rect 135872 121696 135912 121736
rect 135954 121696 135994 121736
rect 136036 121696 136076 121736
rect 136118 121696 136158 121736
rect 136200 121696 136240 121736
rect 150992 121696 151032 121736
rect 151074 121696 151114 121736
rect 151156 121696 151196 121736
rect 151238 121696 151278 121736
rect 151320 121696 151360 121736
rect 74152 120940 74192 120980
rect 74234 120940 74274 120980
rect 74316 120940 74356 120980
rect 74398 120940 74438 120980
rect 74480 120940 74520 120980
rect 89272 120940 89312 120980
rect 89354 120940 89394 120980
rect 89436 120940 89476 120980
rect 89518 120940 89558 120980
rect 89600 120940 89640 120980
rect 104392 120940 104432 120980
rect 104474 120940 104514 120980
rect 104556 120940 104596 120980
rect 104638 120940 104678 120980
rect 104720 120940 104760 120980
rect 119512 120940 119552 120980
rect 119594 120940 119634 120980
rect 119676 120940 119716 120980
rect 119758 120940 119798 120980
rect 119840 120940 119880 120980
rect 134632 120940 134672 120980
rect 134714 120940 134754 120980
rect 134796 120940 134836 120980
rect 134878 120940 134918 120980
rect 134960 120940 135000 120980
rect 149752 120940 149792 120980
rect 149834 120940 149874 120980
rect 149916 120940 149956 120980
rect 149998 120940 150038 120980
rect 150080 120940 150120 120980
rect 75392 120184 75432 120224
rect 75474 120184 75514 120224
rect 75556 120184 75596 120224
rect 75638 120184 75678 120224
rect 75720 120184 75760 120224
rect 90512 120184 90552 120224
rect 90594 120184 90634 120224
rect 90676 120184 90716 120224
rect 90758 120184 90798 120224
rect 90840 120184 90880 120224
rect 105632 120184 105672 120224
rect 105714 120184 105754 120224
rect 105796 120184 105836 120224
rect 105878 120184 105918 120224
rect 105960 120184 106000 120224
rect 120752 120184 120792 120224
rect 120834 120184 120874 120224
rect 120916 120184 120956 120224
rect 120998 120184 121038 120224
rect 121080 120184 121120 120224
rect 135872 120184 135912 120224
rect 135954 120184 135994 120224
rect 136036 120184 136076 120224
rect 136118 120184 136158 120224
rect 136200 120184 136240 120224
rect 150992 120184 151032 120224
rect 151074 120184 151114 120224
rect 151156 120184 151196 120224
rect 151238 120184 151278 120224
rect 151320 120184 151360 120224
rect 74152 119428 74192 119468
rect 74234 119428 74274 119468
rect 74316 119428 74356 119468
rect 74398 119428 74438 119468
rect 74480 119428 74520 119468
rect 89272 119428 89312 119468
rect 89354 119428 89394 119468
rect 89436 119428 89476 119468
rect 89518 119428 89558 119468
rect 89600 119428 89640 119468
rect 104392 119428 104432 119468
rect 104474 119428 104514 119468
rect 104556 119428 104596 119468
rect 104638 119428 104678 119468
rect 104720 119428 104760 119468
rect 119512 119428 119552 119468
rect 119594 119428 119634 119468
rect 119676 119428 119716 119468
rect 119758 119428 119798 119468
rect 119840 119428 119880 119468
rect 134632 119428 134672 119468
rect 134714 119428 134754 119468
rect 134796 119428 134836 119468
rect 134878 119428 134918 119468
rect 134960 119428 135000 119468
rect 149752 119428 149792 119468
rect 149834 119428 149874 119468
rect 149916 119428 149956 119468
rect 149998 119428 150038 119468
rect 150080 119428 150120 119468
rect 75392 118672 75432 118712
rect 75474 118672 75514 118712
rect 75556 118672 75596 118712
rect 75638 118672 75678 118712
rect 75720 118672 75760 118712
rect 90512 118672 90552 118712
rect 90594 118672 90634 118712
rect 90676 118672 90716 118712
rect 90758 118672 90798 118712
rect 90840 118672 90880 118712
rect 105632 118672 105672 118712
rect 105714 118672 105754 118712
rect 105796 118672 105836 118712
rect 105878 118672 105918 118712
rect 105960 118672 106000 118712
rect 120752 118672 120792 118712
rect 120834 118672 120874 118712
rect 120916 118672 120956 118712
rect 120998 118672 121038 118712
rect 121080 118672 121120 118712
rect 135872 118672 135912 118712
rect 135954 118672 135994 118712
rect 136036 118672 136076 118712
rect 136118 118672 136158 118712
rect 136200 118672 136240 118712
rect 150992 118672 151032 118712
rect 151074 118672 151114 118712
rect 151156 118672 151196 118712
rect 151238 118672 151278 118712
rect 151320 118672 151360 118712
rect 74152 117916 74192 117956
rect 74234 117916 74274 117956
rect 74316 117916 74356 117956
rect 74398 117916 74438 117956
rect 74480 117916 74520 117956
rect 89272 117916 89312 117956
rect 89354 117916 89394 117956
rect 89436 117916 89476 117956
rect 89518 117916 89558 117956
rect 89600 117916 89640 117956
rect 104392 117916 104432 117956
rect 104474 117916 104514 117956
rect 104556 117916 104596 117956
rect 104638 117916 104678 117956
rect 104720 117916 104760 117956
rect 119512 117916 119552 117956
rect 119594 117916 119634 117956
rect 119676 117916 119716 117956
rect 119758 117916 119798 117956
rect 119840 117916 119880 117956
rect 134632 117916 134672 117956
rect 134714 117916 134754 117956
rect 134796 117916 134836 117956
rect 134878 117916 134918 117956
rect 134960 117916 135000 117956
rect 149752 117916 149792 117956
rect 149834 117916 149874 117956
rect 149916 117916 149956 117956
rect 149998 117916 150038 117956
rect 150080 117916 150120 117956
rect 75392 117160 75432 117200
rect 75474 117160 75514 117200
rect 75556 117160 75596 117200
rect 75638 117160 75678 117200
rect 75720 117160 75760 117200
rect 90512 117160 90552 117200
rect 90594 117160 90634 117200
rect 90676 117160 90716 117200
rect 90758 117160 90798 117200
rect 90840 117160 90880 117200
rect 105632 117160 105672 117200
rect 105714 117160 105754 117200
rect 105796 117160 105836 117200
rect 105878 117160 105918 117200
rect 105960 117160 106000 117200
rect 120752 117160 120792 117200
rect 120834 117160 120874 117200
rect 120916 117160 120956 117200
rect 120998 117160 121038 117200
rect 121080 117160 121120 117200
rect 135872 117160 135912 117200
rect 135954 117160 135994 117200
rect 136036 117160 136076 117200
rect 136118 117160 136158 117200
rect 136200 117160 136240 117200
rect 150992 117160 151032 117200
rect 151074 117160 151114 117200
rect 151156 117160 151196 117200
rect 151238 117160 151278 117200
rect 151320 117160 151360 117200
rect 74152 116404 74192 116444
rect 74234 116404 74274 116444
rect 74316 116404 74356 116444
rect 74398 116404 74438 116444
rect 74480 116404 74520 116444
rect 89272 116404 89312 116444
rect 89354 116404 89394 116444
rect 89436 116404 89476 116444
rect 89518 116404 89558 116444
rect 89600 116404 89640 116444
rect 104392 116404 104432 116444
rect 104474 116404 104514 116444
rect 104556 116404 104596 116444
rect 104638 116404 104678 116444
rect 104720 116404 104760 116444
rect 119512 116404 119552 116444
rect 119594 116404 119634 116444
rect 119676 116404 119716 116444
rect 119758 116404 119798 116444
rect 119840 116404 119880 116444
rect 134632 116404 134672 116444
rect 134714 116404 134754 116444
rect 134796 116404 134836 116444
rect 134878 116404 134918 116444
rect 134960 116404 135000 116444
rect 149752 116404 149792 116444
rect 149834 116404 149874 116444
rect 149916 116404 149956 116444
rect 149998 116404 150038 116444
rect 150080 116404 150120 116444
rect 75392 115648 75432 115688
rect 75474 115648 75514 115688
rect 75556 115648 75596 115688
rect 75638 115648 75678 115688
rect 75720 115648 75760 115688
rect 90512 115648 90552 115688
rect 90594 115648 90634 115688
rect 90676 115648 90716 115688
rect 90758 115648 90798 115688
rect 90840 115648 90880 115688
rect 105632 115648 105672 115688
rect 105714 115648 105754 115688
rect 105796 115648 105836 115688
rect 105878 115648 105918 115688
rect 105960 115648 106000 115688
rect 120752 115648 120792 115688
rect 120834 115648 120874 115688
rect 120916 115648 120956 115688
rect 120998 115648 121038 115688
rect 121080 115648 121120 115688
rect 135872 115648 135912 115688
rect 135954 115648 135994 115688
rect 136036 115648 136076 115688
rect 136118 115648 136158 115688
rect 136200 115648 136240 115688
rect 150992 115648 151032 115688
rect 151074 115648 151114 115688
rect 151156 115648 151196 115688
rect 151238 115648 151278 115688
rect 151320 115648 151360 115688
rect 74152 114892 74192 114932
rect 74234 114892 74274 114932
rect 74316 114892 74356 114932
rect 74398 114892 74438 114932
rect 74480 114892 74520 114932
rect 89272 114892 89312 114932
rect 89354 114892 89394 114932
rect 89436 114892 89476 114932
rect 89518 114892 89558 114932
rect 89600 114892 89640 114932
rect 104392 114892 104432 114932
rect 104474 114892 104514 114932
rect 104556 114892 104596 114932
rect 104638 114892 104678 114932
rect 104720 114892 104760 114932
rect 119512 114892 119552 114932
rect 119594 114892 119634 114932
rect 119676 114892 119716 114932
rect 119758 114892 119798 114932
rect 119840 114892 119880 114932
rect 134632 114892 134672 114932
rect 134714 114892 134754 114932
rect 134796 114892 134836 114932
rect 134878 114892 134918 114932
rect 134960 114892 135000 114932
rect 149752 114892 149792 114932
rect 149834 114892 149874 114932
rect 149916 114892 149956 114932
rect 149998 114892 150038 114932
rect 150080 114892 150120 114932
rect 75392 114136 75432 114176
rect 75474 114136 75514 114176
rect 75556 114136 75596 114176
rect 75638 114136 75678 114176
rect 75720 114136 75760 114176
rect 90512 114136 90552 114176
rect 90594 114136 90634 114176
rect 90676 114136 90716 114176
rect 90758 114136 90798 114176
rect 90840 114136 90880 114176
rect 105632 114136 105672 114176
rect 105714 114136 105754 114176
rect 105796 114136 105836 114176
rect 105878 114136 105918 114176
rect 105960 114136 106000 114176
rect 120752 114136 120792 114176
rect 120834 114136 120874 114176
rect 120916 114136 120956 114176
rect 120998 114136 121038 114176
rect 121080 114136 121120 114176
rect 135872 114136 135912 114176
rect 135954 114136 135994 114176
rect 136036 114136 136076 114176
rect 136118 114136 136158 114176
rect 136200 114136 136240 114176
rect 150992 114136 151032 114176
rect 151074 114136 151114 114176
rect 151156 114136 151196 114176
rect 151238 114136 151278 114176
rect 151320 114136 151360 114176
rect 74152 113380 74192 113420
rect 74234 113380 74274 113420
rect 74316 113380 74356 113420
rect 74398 113380 74438 113420
rect 74480 113380 74520 113420
rect 89272 113380 89312 113420
rect 89354 113380 89394 113420
rect 89436 113380 89476 113420
rect 89518 113380 89558 113420
rect 89600 113380 89640 113420
rect 104392 113380 104432 113420
rect 104474 113380 104514 113420
rect 104556 113380 104596 113420
rect 104638 113380 104678 113420
rect 104720 113380 104760 113420
rect 119512 113380 119552 113420
rect 119594 113380 119634 113420
rect 119676 113380 119716 113420
rect 119758 113380 119798 113420
rect 119840 113380 119880 113420
rect 134632 113380 134672 113420
rect 134714 113380 134754 113420
rect 134796 113380 134836 113420
rect 134878 113380 134918 113420
rect 134960 113380 135000 113420
rect 149752 113380 149792 113420
rect 149834 113380 149874 113420
rect 149916 113380 149956 113420
rect 149998 113380 150038 113420
rect 150080 113380 150120 113420
rect 75392 112624 75432 112664
rect 75474 112624 75514 112664
rect 75556 112624 75596 112664
rect 75638 112624 75678 112664
rect 75720 112624 75760 112664
rect 90512 112624 90552 112664
rect 90594 112624 90634 112664
rect 90676 112624 90716 112664
rect 90758 112624 90798 112664
rect 90840 112624 90880 112664
rect 105632 112624 105672 112664
rect 105714 112624 105754 112664
rect 105796 112624 105836 112664
rect 105878 112624 105918 112664
rect 105960 112624 106000 112664
rect 120752 112624 120792 112664
rect 120834 112624 120874 112664
rect 120916 112624 120956 112664
rect 120998 112624 121038 112664
rect 121080 112624 121120 112664
rect 135872 112624 135912 112664
rect 135954 112624 135994 112664
rect 136036 112624 136076 112664
rect 136118 112624 136158 112664
rect 136200 112624 136240 112664
rect 150992 112624 151032 112664
rect 151074 112624 151114 112664
rect 151156 112624 151196 112664
rect 151238 112624 151278 112664
rect 151320 112624 151360 112664
rect 74152 111868 74192 111908
rect 74234 111868 74274 111908
rect 74316 111868 74356 111908
rect 74398 111868 74438 111908
rect 74480 111868 74520 111908
rect 89272 111868 89312 111908
rect 89354 111868 89394 111908
rect 89436 111868 89476 111908
rect 89518 111868 89558 111908
rect 89600 111868 89640 111908
rect 104392 111868 104432 111908
rect 104474 111868 104514 111908
rect 104556 111868 104596 111908
rect 104638 111868 104678 111908
rect 104720 111868 104760 111908
rect 119512 111868 119552 111908
rect 119594 111868 119634 111908
rect 119676 111868 119716 111908
rect 119758 111868 119798 111908
rect 119840 111868 119880 111908
rect 134632 111868 134672 111908
rect 134714 111868 134754 111908
rect 134796 111868 134836 111908
rect 134878 111868 134918 111908
rect 134960 111868 135000 111908
rect 149752 111868 149792 111908
rect 149834 111868 149874 111908
rect 149916 111868 149956 111908
rect 149998 111868 150038 111908
rect 150080 111868 150120 111908
rect 75392 111112 75432 111152
rect 75474 111112 75514 111152
rect 75556 111112 75596 111152
rect 75638 111112 75678 111152
rect 75720 111112 75760 111152
rect 90512 111112 90552 111152
rect 90594 111112 90634 111152
rect 90676 111112 90716 111152
rect 90758 111112 90798 111152
rect 90840 111112 90880 111152
rect 105632 111112 105672 111152
rect 105714 111112 105754 111152
rect 105796 111112 105836 111152
rect 105878 111112 105918 111152
rect 105960 111112 106000 111152
rect 120752 111112 120792 111152
rect 120834 111112 120874 111152
rect 120916 111112 120956 111152
rect 120998 111112 121038 111152
rect 121080 111112 121120 111152
rect 135872 111112 135912 111152
rect 135954 111112 135994 111152
rect 136036 111112 136076 111152
rect 136118 111112 136158 111152
rect 136200 111112 136240 111152
rect 150992 111112 151032 111152
rect 151074 111112 151114 111152
rect 151156 111112 151196 111152
rect 151238 111112 151278 111152
rect 151320 111112 151360 111152
rect 74152 110356 74192 110396
rect 74234 110356 74274 110396
rect 74316 110356 74356 110396
rect 74398 110356 74438 110396
rect 74480 110356 74520 110396
rect 89272 110356 89312 110396
rect 89354 110356 89394 110396
rect 89436 110356 89476 110396
rect 89518 110356 89558 110396
rect 89600 110356 89640 110396
rect 104392 110356 104432 110396
rect 104474 110356 104514 110396
rect 104556 110356 104596 110396
rect 104638 110356 104678 110396
rect 104720 110356 104760 110396
rect 119512 110356 119552 110396
rect 119594 110356 119634 110396
rect 119676 110356 119716 110396
rect 119758 110356 119798 110396
rect 119840 110356 119880 110396
rect 134632 110356 134672 110396
rect 134714 110356 134754 110396
rect 134796 110356 134836 110396
rect 134878 110356 134918 110396
rect 134960 110356 135000 110396
rect 149752 110356 149792 110396
rect 149834 110356 149874 110396
rect 149916 110356 149956 110396
rect 149998 110356 150038 110396
rect 150080 110356 150120 110396
rect 75392 109600 75432 109640
rect 75474 109600 75514 109640
rect 75556 109600 75596 109640
rect 75638 109600 75678 109640
rect 75720 109600 75760 109640
rect 90512 109600 90552 109640
rect 90594 109600 90634 109640
rect 90676 109600 90716 109640
rect 90758 109600 90798 109640
rect 90840 109600 90880 109640
rect 105632 109600 105672 109640
rect 105714 109600 105754 109640
rect 105796 109600 105836 109640
rect 105878 109600 105918 109640
rect 105960 109600 106000 109640
rect 120752 109600 120792 109640
rect 120834 109600 120874 109640
rect 120916 109600 120956 109640
rect 120998 109600 121038 109640
rect 121080 109600 121120 109640
rect 135872 109600 135912 109640
rect 135954 109600 135994 109640
rect 136036 109600 136076 109640
rect 136118 109600 136158 109640
rect 136200 109600 136240 109640
rect 150992 109600 151032 109640
rect 151074 109600 151114 109640
rect 151156 109600 151196 109640
rect 151238 109600 151278 109640
rect 151320 109600 151360 109640
rect 74152 108844 74192 108884
rect 74234 108844 74274 108884
rect 74316 108844 74356 108884
rect 74398 108844 74438 108884
rect 74480 108844 74520 108884
rect 89272 108844 89312 108884
rect 89354 108844 89394 108884
rect 89436 108844 89476 108884
rect 89518 108844 89558 108884
rect 89600 108844 89640 108884
rect 104392 108844 104432 108884
rect 104474 108844 104514 108884
rect 104556 108844 104596 108884
rect 104638 108844 104678 108884
rect 104720 108844 104760 108884
rect 119512 108844 119552 108884
rect 119594 108844 119634 108884
rect 119676 108844 119716 108884
rect 119758 108844 119798 108884
rect 119840 108844 119880 108884
rect 134632 108844 134672 108884
rect 134714 108844 134754 108884
rect 134796 108844 134836 108884
rect 134878 108844 134918 108884
rect 134960 108844 135000 108884
rect 149752 108844 149792 108884
rect 149834 108844 149874 108884
rect 149916 108844 149956 108884
rect 149998 108844 150038 108884
rect 150080 108844 150120 108884
rect 75392 108088 75432 108128
rect 75474 108088 75514 108128
rect 75556 108088 75596 108128
rect 75638 108088 75678 108128
rect 75720 108088 75760 108128
rect 90512 108088 90552 108128
rect 90594 108088 90634 108128
rect 90676 108088 90716 108128
rect 90758 108088 90798 108128
rect 90840 108088 90880 108128
rect 105632 108088 105672 108128
rect 105714 108088 105754 108128
rect 105796 108088 105836 108128
rect 105878 108088 105918 108128
rect 105960 108088 106000 108128
rect 120752 108088 120792 108128
rect 120834 108088 120874 108128
rect 120916 108088 120956 108128
rect 120998 108088 121038 108128
rect 121080 108088 121120 108128
rect 135872 108088 135912 108128
rect 135954 108088 135994 108128
rect 136036 108088 136076 108128
rect 136118 108088 136158 108128
rect 136200 108088 136240 108128
rect 150992 108088 151032 108128
rect 151074 108088 151114 108128
rect 151156 108088 151196 108128
rect 151238 108088 151278 108128
rect 151320 108088 151360 108128
rect 74152 107332 74192 107372
rect 74234 107332 74274 107372
rect 74316 107332 74356 107372
rect 74398 107332 74438 107372
rect 74480 107332 74520 107372
rect 89272 107332 89312 107372
rect 89354 107332 89394 107372
rect 89436 107332 89476 107372
rect 89518 107332 89558 107372
rect 89600 107332 89640 107372
rect 104392 107332 104432 107372
rect 104474 107332 104514 107372
rect 104556 107332 104596 107372
rect 104638 107332 104678 107372
rect 104720 107332 104760 107372
rect 119512 107332 119552 107372
rect 119594 107332 119634 107372
rect 119676 107332 119716 107372
rect 119758 107332 119798 107372
rect 119840 107332 119880 107372
rect 134632 107332 134672 107372
rect 134714 107332 134754 107372
rect 134796 107332 134836 107372
rect 134878 107332 134918 107372
rect 134960 107332 135000 107372
rect 149752 107332 149792 107372
rect 149834 107332 149874 107372
rect 149916 107332 149956 107372
rect 149998 107332 150038 107372
rect 150080 107332 150120 107372
rect 75392 106576 75432 106616
rect 75474 106576 75514 106616
rect 75556 106576 75596 106616
rect 75638 106576 75678 106616
rect 75720 106576 75760 106616
rect 90512 106576 90552 106616
rect 90594 106576 90634 106616
rect 90676 106576 90716 106616
rect 90758 106576 90798 106616
rect 90840 106576 90880 106616
rect 105632 106576 105672 106616
rect 105714 106576 105754 106616
rect 105796 106576 105836 106616
rect 105878 106576 105918 106616
rect 105960 106576 106000 106616
rect 120752 106576 120792 106616
rect 120834 106576 120874 106616
rect 120916 106576 120956 106616
rect 120998 106576 121038 106616
rect 121080 106576 121120 106616
rect 135872 106576 135912 106616
rect 135954 106576 135994 106616
rect 136036 106576 136076 106616
rect 136118 106576 136158 106616
rect 136200 106576 136240 106616
rect 150992 106576 151032 106616
rect 151074 106576 151114 106616
rect 151156 106576 151196 106616
rect 151238 106576 151278 106616
rect 151320 106576 151360 106616
rect 74152 105820 74192 105860
rect 74234 105820 74274 105860
rect 74316 105820 74356 105860
rect 74398 105820 74438 105860
rect 74480 105820 74520 105860
rect 89272 105820 89312 105860
rect 89354 105820 89394 105860
rect 89436 105820 89476 105860
rect 89518 105820 89558 105860
rect 89600 105820 89640 105860
rect 104392 105820 104432 105860
rect 104474 105820 104514 105860
rect 104556 105820 104596 105860
rect 104638 105820 104678 105860
rect 104720 105820 104760 105860
rect 119512 105820 119552 105860
rect 119594 105820 119634 105860
rect 119676 105820 119716 105860
rect 119758 105820 119798 105860
rect 119840 105820 119880 105860
rect 134632 105820 134672 105860
rect 134714 105820 134754 105860
rect 134796 105820 134836 105860
rect 134878 105820 134918 105860
rect 134960 105820 135000 105860
rect 149752 105820 149792 105860
rect 149834 105820 149874 105860
rect 149916 105820 149956 105860
rect 149998 105820 150038 105860
rect 150080 105820 150120 105860
rect 75392 105064 75432 105104
rect 75474 105064 75514 105104
rect 75556 105064 75596 105104
rect 75638 105064 75678 105104
rect 75720 105064 75760 105104
rect 90512 105064 90552 105104
rect 90594 105064 90634 105104
rect 90676 105064 90716 105104
rect 90758 105064 90798 105104
rect 90840 105064 90880 105104
rect 105632 105064 105672 105104
rect 105714 105064 105754 105104
rect 105796 105064 105836 105104
rect 105878 105064 105918 105104
rect 105960 105064 106000 105104
rect 120752 105064 120792 105104
rect 120834 105064 120874 105104
rect 120916 105064 120956 105104
rect 120998 105064 121038 105104
rect 121080 105064 121120 105104
rect 135872 105064 135912 105104
rect 135954 105064 135994 105104
rect 136036 105064 136076 105104
rect 136118 105064 136158 105104
rect 136200 105064 136240 105104
rect 150992 105064 151032 105104
rect 151074 105064 151114 105104
rect 151156 105064 151196 105104
rect 151238 105064 151278 105104
rect 151320 105064 151360 105104
rect 74152 104308 74192 104348
rect 74234 104308 74274 104348
rect 74316 104308 74356 104348
rect 74398 104308 74438 104348
rect 74480 104308 74520 104348
rect 89272 104308 89312 104348
rect 89354 104308 89394 104348
rect 89436 104308 89476 104348
rect 89518 104308 89558 104348
rect 89600 104308 89640 104348
rect 104392 104308 104432 104348
rect 104474 104308 104514 104348
rect 104556 104308 104596 104348
rect 104638 104308 104678 104348
rect 104720 104308 104760 104348
rect 119512 104308 119552 104348
rect 119594 104308 119634 104348
rect 119676 104308 119716 104348
rect 119758 104308 119798 104348
rect 119840 104308 119880 104348
rect 134632 104308 134672 104348
rect 134714 104308 134754 104348
rect 134796 104308 134836 104348
rect 134878 104308 134918 104348
rect 134960 104308 135000 104348
rect 149752 104308 149792 104348
rect 149834 104308 149874 104348
rect 149916 104308 149956 104348
rect 149998 104308 150038 104348
rect 150080 104308 150120 104348
rect 75392 103552 75432 103592
rect 75474 103552 75514 103592
rect 75556 103552 75596 103592
rect 75638 103552 75678 103592
rect 75720 103552 75760 103592
rect 90512 103552 90552 103592
rect 90594 103552 90634 103592
rect 90676 103552 90716 103592
rect 90758 103552 90798 103592
rect 90840 103552 90880 103592
rect 105632 103552 105672 103592
rect 105714 103552 105754 103592
rect 105796 103552 105836 103592
rect 105878 103552 105918 103592
rect 105960 103552 106000 103592
rect 120752 103552 120792 103592
rect 120834 103552 120874 103592
rect 120916 103552 120956 103592
rect 120998 103552 121038 103592
rect 121080 103552 121120 103592
rect 135872 103552 135912 103592
rect 135954 103552 135994 103592
rect 136036 103552 136076 103592
rect 136118 103552 136158 103592
rect 136200 103552 136240 103592
rect 150992 103552 151032 103592
rect 151074 103552 151114 103592
rect 151156 103552 151196 103592
rect 151238 103552 151278 103592
rect 151320 103552 151360 103592
rect 74152 102796 74192 102836
rect 74234 102796 74274 102836
rect 74316 102796 74356 102836
rect 74398 102796 74438 102836
rect 74480 102796 74520 102836
rect 89272 102796 89312 102836
rect 89354 102796 89394 102836
rect 89436 102796 89476 102836
rect 89518 102796 89558 102836
rect 89600 102796 89640 102836
rect 104392 102796 104432 102836
rect 104474 102796 104514 102836
rect 104556 102796 104596 102836
rect 104638 102796 104678 102836
rect 104720 102796 104760 102836
rect 119512 102796 119552 102836
rect 119594 102796 119634 102836
rect 119676 102796 119716 102836
rect 119758 102796 119798 102836
rect 119840 102796 119880 102836
rect 134632 102796 134672 102836
rect 134714 102796 134754 102836
rect 134796 102796 134836 102836
rect 134878 102796 134918 102836
rect 134960 102796 135000 102836
rect 149752 102796 149792 102836
rect 149834 102796 149874 102836
rect 149916 102796 149956 102836
rect 149998 102796 150038 102836
rect 150080 102796 150120 102836
rect 75392 102040 75432 102080
rect 75474 102040 75514 102080
rect 75556 102040 75596 102080
rect 75638 102040 75678 102080
rect 75720 102040 75760 102080
rect 90512 102040 90552 102080
rect 90594 102040 90634 102080
rect 90676 102040 90716 102080
rect 90758 102040 90798 102080
rect 90840 102040 90880 102080
rect 105632 102040 105672 102080
rect 105714 102040 105754 102080
rect 105796 102040 105836 102080
rect 105878 102040 105918 102080
rect 105960 102040 106000 102080
rect 120752 102040 120792 102080
rect 120834 102040 120874 102080
rect 120916 102040 120956 102080
rect 120998 102040 121038 102080
rect 121080 102040 121120 102080
rect 135872 102040 135912 102080
rect 135954 102040 135994 102080
rect 136036 102040 136076 102080
rect 136118 102040 136158 102080
rect 136200 102040 136240 102080
rect 150992 102040 151032 102080
rect 151074 102040 151114 102080
rect 151156 102040 151196 102080
rect 151238 102040 151278 102080
rect 151320 102040 151360 102080
rect 74152 101284 74192 101324
rect 74234 101284 74274 101324
rect 74316 101284 74356 101324
rect 74398 101284 74438 101324
rect 74480 101284 74520 101324
rect 89272 101284 89312 101324
rect 89354 101284 89394 101324
rect 89436 101284 89476 101324
rect 89518 101284 89558 101324
rect 89600 101284 89640 101324
rect 104392 101284 104432 101324
rect 104474 101284 104514 101324
rect 104556 101284 104596 101324
rect 104638 101284 104678 101324
rect 104720 101284 104760 101324
rect 119512 101284 119552 101324
rect 119594 101284 119634 101324
rect 119676 101284 119716 101324
rect 119758 101284 119798 101324
rect 119840 101284 119880 101324
rect 134632 101284 134672 101324
rect 134714 101284 134754 101324
rect 134796 101284 134836 101324
rect 134878 101284 134918 101324
rect 134960 101284 135000 101324
rect 149752 101284 149792 101324
rect 149834 101284 149874 101324
rect 149916 101284 149956 101324
rect 149998 101284 150038 101324
rect 150080 101284 150120 101324
rect 75392 100528 75432 100568
rect 75474 100528 75514 100568
rect 75556 100528 75596 100568
rect 75638 100528 75678 100568
rect 75720 100528 75760 100568
rect 90512 100528 90552 100568
rect 90594 100528 90634 100568
rect 90676 100528 90716 100568
rect 90758 100528 90798 100568
rect 90840 100528 90880 100568
rect 105632 100528 105672 100568
rect 105714 100528 105754 100568
rect 105796 100528 105836 100568
rect 105878 100528 105918 100568
rect 105960 100528 106000 100568
rect 120752 100528 120792 100568
rect 120834 100528 120874 100568
rect 120916 100528 120956 100568
rect 120998 100528 121038 100568
rect 121080 100528 121120 100568
rect 135872 100528 135912 100568
rect 135954 100528 135994 100568
rect 136036 100528 136076 100568
rect 136118 100528 136158 100568
rect 136200 100528 136240 100568
rect 150992 100528 151032 100568
rect 151074 100528 151114 100568
rect 151156 100528 151196 100568
rect 151238 100528 151278 100568
rect 151320 100528 151360 100568
rect 74152 99772 74192 99812
rect 74234 99772 74274 99812
rect 74316 99772 74356 99812
rect 74398 99772 74438 99812
rect 74480 99772 74520 99812
rect 89272 99772 89312 99812
rect 89354 99772 89394 99812
rect 89436 99772 89476 99812
rect 89518 99772 89558 99812
rect 89600 99772 89640 99812
rect 104392 99772 104432 99812
rect 104474 99772 104514 99812
rect 104556 99772 104596 99812
rect 104638 99772 104678 99812
rect 104720 99772 104760 99812
rect 119512 99772 119552 99812
rect 119594 99772 119634 99812
rect 119676 99772 119716 99812
rect 119758 99772 119798 99812
rect 119840 99772 119880 99812
rect 134632 99772 134672 99812
rect 134714 99772 134754 99812
rect 134796 99772 134836 99812
rect 134878 99772 134918 99812
rect 134960 99772 135000 99812
rect 149752 99772 149792 99812
rect 149834 99772 149874 99812
rect 149916 99772 149956 99812
rect 149998 99772 150038 99812
rect 150080 99772 150120 99812
rect 75392 99016 75432 99056
rect 75474 99016 75514 99056
rect 75556 99016 75596 99056
rect 75638 99016 75678 99056
rect 75720 99016 75760 99056
rect 90512 99016 90552 99056
rect 90594 99016 90634 99056
rect 90676 99016 90716 99056
rect 90758 99016 90798 99056
rect 90840 99016 90880 99056
rect 105632 99016 105672 99056
rect 105714 99016 105754 99056
rect 105796 99016 105836 99056
rect 105878 99016 105918 99056
rect 105960 99016 106000 99056
rect 120752 99016 120792 99056
rect 120834 99016 120874 99056
rect 120916 99016 120956 99056
rect 120998 99016 121038 99056
rect 121080 99016 121120 99056
rect 135872 99016 135912 99056
rect 135954 99016 135994 99056
rect 136036 99016 136076 99056
rect 136118 99016 136158 99056
rect 136200 99016 136240 99056
rect 150992 99016 151032 99056
rect 151074 99016 151114 99056
rect 151156 99016 151196 99056
rect 151238 99016 151278 99056
rect 151320 99016 151360 99056
rect 74152 98260 74192 98300
rect 74234 98260 74274 98300
rect 74316 98260 74356 98300
rect 74398 98260 74438 98300
rect 74480 98260 74520 98300
rect 89272 98260 89312 98300
rect 89354 98260 89394 98300
rect 89436 98260 89476 98300
rect 89518 98260 89558 98300
rect 89600 98260 89640 98300
rect 104392 98260 104432 98300
rect 104474 98260 104514 98300
rect 104556 98260 104596 98300
rect 104638 98260 104678 98300
rect 104720 98260 104760 98300
rect 119512 98260 119552 98300
rect 119594 98260 119634 98300
rect 119676 98260 119716 98300
rect 119758 98260 119798 98300
rect 119840 98260 119880 98300
rect 134632 98260 134672 98300
rect 134714 98260 134754 98300
rect 134796 98260 134836 98300
rect 134878 98260 134918 98300
rect 134960 98260 135000 98300
rect 149752 98260 149792 98300
rect 149834 98260 149874 98300
rect 149916 98260 149956 98300
rect 149998 98260 150038 98300
rect 150080 98260 150120 98300
rect 75392 97504 75432 97544
rect 75474 97504 75514 97544
rect 75556 97504 75596 97544
rect 75638 97504 75678 97544
rect 75720 97504 75760 97544
rect 90512 97504 90552 97544
rect 90594 97504 90634 97544
rect 90676 97504 90716 97544
rect 90758 97504 90798 97544
rect 90840 97504 90880 97544
rect 105632 97504 105672 97544
rect 105714 97504 105754 97544
rect 105796 97504 105836 97544
rect 105878 97504 105918 97544
rect 105960 97504 106000 97544
rect 120752 97504 120792 97544
rect 120834 97504 120874 97544
rect 120916 97504 120956 97544
rect 120998 97504 121038 97544
rect 121080 97504 121120 97544
rect 135872 97504 135912 97544
rect 135954 97504 135994 97544
rect 136036 97504 136076 97544
rect 136118 97504 136158 97544
rect 136200 97504 136240 97544
rect 150992 97504 151032 97544
rect 151074 97504 151114 97544
rect 151156 97504 151196 97544
rect 151238 97504 151278 97544
rect 151320 97504 151360 97544
rect 74152 96748 74192 96788
rect 74234 96748 74274 96788
rect 74316 96748 74356 96788
rect 74398 96748 74438 96788
rect 74480 96748 74520 96788
rect 89272 96748 89312 96788
rect 89354 96748 89394 96788
rect 89436 96748 89476 96788
rect 89518 96748 89558 96788
rect 89600 96748 89640 96788
rect 104392 96748 104432 96788
rect 104474 96748 104514 96788
rect 104556 96748 104596 96788
rect 104638 96748 104678 96788
rect 104720 96748 104760 96788
rect 119512 96748 119552 96788
rect 119594 96748 119634 96788
rect 119676 96748 119716 96788
rect 119758 96748 119798 96788
rect 119840 96748 119880 96788
rect 134632 96748 134672 96788
rect 134714 96748 134754 96788
rect 134796 96748 134836 96788
rect 134878 96748 134918 96788
rect 134960 96748 135000 96788
rect 149752 96748 149792 96788
rect 149834 96748 149874 96788
rect 149916 96748 149956 96788
rect 149998 96748 150038 96788
rect 150080 96748 150120 96788
rect 75392 95992 75432 96032
rect 75474 95992 75514 96032
rect 75556 95992 75596 96032
rect 75638 95992 75678 96032
rect 75720 95992 75760 96032
rect 90512 95992 90552 96032
rect 90594 95992 90634 96032
rect 90676 95992 90716 96032
rect 90758 95992 90798 96032
rect 90840 95992 90880 96032
rect 105632 95992 105672 96032
rect 105714 95992 105754 96032
rect 105796 95992 105836 96032
rect 105878 95992 105918 96032
rect 105960 95992 106000 96032
rect 120752 95992 120792 96032
rect 120834 95992 120874 96032
rect 120916 95992 120956 96032
rect 120998 95992 121038 96032
rect 121080 95992 121120 96032
rect 135872 95992 135912 96032
rect 135954 95992 135994 96032
rect 136036 95992 136076 96032
rect 136118 95992 136158 96032
rect 136200 95992 136240 96032
rect 150992 95992 151032 96032
rect 151074 95992 151114 96032
rect 151156 95992 151196 96032
rect 151238 95992 151278 96032
rect 151320 95992 151360 96032
rect 74152 95236 74192 95276
rect 74234 95236 74274 95276
rect 74316 95236 74356 95276
rect 74398 95236 74438 95276
rect 74480 95236 74520 95276
rect 89272 95236 89312 95276
rect 89354 95236 89394 95276
rect 89436 95236 89476 95276
rect 89518 95236 89558 95276
rect 89600 95236 89640 95276
rect 104392 95236 104432 95276
rect 104474 95236 104514 95276
rect 104556 95236 104596 95276
rect 104638 95236 104678 95276
rect 104720 95236 104760 95276
rect 119512 95236 119552 95276
rect 119594 95236 119634 95276
rect 119676 95236 119716 95276
rect 119758 95236 119798 95276
rect 119840 95236 119880 95276
rect 134632 95236 134672 95276
rect 134714 95236 134754 95276
rect 134796 95236 134836 95276
rect 134878 95236 134918 95276
rect 134960 95236 135000 95276
rect 149752 95236 149792 95276
rect 149834 95236 149874 95276
rect 149916 95236 149956 95276
rect 149998 95236 150038 95276
rect 150080 95236 150120 95276
rect 75392 94480 75432 94520
rect 75474 94480 75514 94520
rect 75556 94480 75596 94520
rect 75638 94480 75678 94520
rect 75720 94480 75760 94520
rect 90512 94480 90552 94520
rect 90594 94480 90634 94520
rect 90676 94480 90716 94520
rect 90758 94480 90798 94520
rect 90840 94480 90880 94520
rect 105632 94480 105672 94520
rect 105714 94480 105754 94520
rect 105796 94480 105836 94520
rect 105878 94480 105918 94520
rect 105960 94480 106000 94520
rect 120752 94480 120792 94520
rect 120834 94480 120874 94520
rect 120916 94480 120956 94520
rect 120998 94480 121038 94520
rect 121080 94480 121120 94520
rect 135872 94480 135912 94520
rect 135954 94480 135994 94520
rect 136036 94480 136076 94520
rect 136118 94480 136158 94520
rect 136200 94480 136240 94520
rect 150992 94480 151032 94520
rect 151074 94480 151114 94520
rect 151156 94480 151196 94520
rect 151238 94480 151278 94520
rect 151320 94480 151360 94520
rect 74152 93724 74192 93764
rect 74234 93724 74274 93764
rect 74316 93724 74356 93764
rect 74398 93724 74438 93764
rect 74480 93724 74520 93764
rect 89272 93724 89312 93764
rect 89354 93724 89394 93764
rect 89436 93724 89476 93764
rect 89518 93724 89558 93764
rect 89600 93724 89640 93764
rect 104392 93724 104432 93764
rect 104474 93724 104514 93764
rect 104556 93724 104596 93764
rect 104638 93724 104678 93764
rect 104720 93724 104760 93764
rect 119512 93724 119552 93764
rect 119594 93724 119634 93764
rect 119676 93724 119716 93764
rect 119758 93724 119798 93764
rect 119840 93724 119880 93764
rect 134632 93724 134672 93764
rect 134714 93724 134754 93764
rect 134796 93724 134836 93764
rect 134878 93724 134918 93764
rect 134960 93724 135000 93764
rect 149752 93724 149792 93764
rect 149834 93724 149874 93764
rect 149916 93724 149956 93764
rect 149998 93724 150038 93764
rect 150080 93724 150120 93764
rect 75392 92968 75432 93008
rect 75474 92968 75514 93008
rect 75556 92968 75596 93008
rect 75638 92968 75678 93008
rect 75720 92968 75760 93008
rect 90512 92968 90552 93008
rect 90594 92968 90634 93008
rect 90676 92968 90716 93008
rect 90758 92968 90798 93008
rect 90840 92968 90880 93008
rect 105632 92968 105672 93008
rect 105714 92968 105754 93008
rect 105796 92968 105836 93008
rect 105878 92968 105918 93008
rect 105960 92968 106000 93008
rect 120752 92968 120792 93008
rect 120834 92968 120874 93008
rect 120916 92968 120956 93008
rect 120998 92968 121038 93008
rect 121080 92968 121120 93008
rect 135872 92968 135912 93008
rect 135954 92968 135994 93008
rect 136036 92968 136076 93008
rect 136118 92968 136158 93008
rect 136200 92968 136240 93008
rect 150992 92968 151032 93008
rect 151074 92968 151114 93008
rect 151156 92968 151196 93008
rect 151238 92968 151278 93008
rect 151320 92968 151360 93008
rect 74152 92212 74192 92252
rect 74234 92212 74274 92252
rect 74316 92212 74356 92252
rect 74398 92212 74438 92252
rect 74480 92212 74520 92252
rect 89272 92212 89312 92252
rect 89354 92212 89394 92252
rect 89436 92212 89476 92252
rect 89518 92212 89558 92252
rect 89600 92212 89640 92252
rect 104392 92212 104432 92252
rect 104474 92212 104514 92252
rect 104556 92212 104596 92252
rect 104638 92212 104678 92252
rect 104720 92212 104760 92252
rect 119512 92212 119552 92252
rect 119594 92212 119634 92252
rect 119676 92212 119716 92252
rect 119758 92212 119798 92252
rect 119840 92212 119880 92252
rect 134632 92212 134672 92252
rect 134714 92212 134754 92252
rect 134796 92212 134836 92252
rect 134878 92212 134918 92252
rect 134960 92212 135000 92252
rect 149752 92212 149792 92252
rect 149834 92212 149874 92252
rect 149916 92212 149956 92252
rect 149998 92212 150038 92252
rect 150080 92212 150120 92252
rect 75392 91456 75432 91496
rect 75474 91456 75514 91496
rect 75556 91456 75596 91496
rect 75638 91456 75678 91496
rect 75720 91456 75760 91496
rect 90512 91456 90552 91496
rect 90594 91456 90634 91496
rect 90676 91456 90716 91496
rect 90758 91456 90798 91496
rect 90840 91456 90880 91496
rect 105632 91456 105672 91496
rect 105714 91456 105754 91496
rect 105796 91456 105836 91496
rect 105878 91456 105918 91496
rect 105960 91456 106000 91496
rect 120752 91456 120792 91496
rect 120834 91456 120874 91496
rect 120916 91456 120956 91496
rect 120998 91456 121038 91496
rect 121080 91456 121120 91496
rect 135872 91456 135912 91496
rect 135954 91456 135994 91496
rect 136036 91456 136076 91496
rect 136118 91456 136158 91496
rect 136200 91456 136240 91496
rect 150992 91456 151032 91496
rect 151074 91456 151114 91496
rect 151156 91456 151196 91496
rect 151238 91456 151278 91496
rect 151320 91456 151360 91496
rect 74152 90700 74192 90740
rect 74234 90700 74274 90740
rect 74316 90700 74356 90740
rect 74398 90700 74438 90740
rect 74480 90700 74520 90740
rect 89272 90700 89312 90740
rect 89354 90700 89394 90740
rect 89436 90700 89476 90740
rect 89518 90700 89558 90740
rect 89600 90700 89640 90740
rect 104392 90700 104432 90740
rect 104474 90700 104514 90740
rect 104556 90700 104596 90740
rect 104638 90700 104678 90740
rect 104720 90700 104760 90740
rect 119512 90700 119552 90740
rect 119594 90700 119634 90740
rect 119676 90700 119716 90740
rect 119758 90700 119798 90740
rect 119840 90700 119880 90740
rect 134632 90700 134672 90740
rect 134714 90700 134754 90740
rect 134796 90700 134836 90740
rect 134878 90700 134918 90740
rect 134960 90700 135000 90740
rect 149752 90700 149792 90740
rect 149834 90700 149874 90740
rect 149916 90700 149956 90740
rect 149998 90700 150038 90740
rect 150080 90700 150120 90740
rect 75392 89944 75432 89984
rect 75474 89944 75514 89984
rect 75556 89944 75596 89984
rect 75638 89944 75678 89984
rect 75720 89944 75760 89984
rect 90512 89944 90552 89984
rect 90594 89944 90634 89984
rect 90676 89944 90716 89984
rect 90758 89944 90798 89984
rect 90840 89944 90880 89984
rect 105632 89944 105672 89984
rect 105714 89944 105754 89984
rect 105796 89944 105836 89984
rect 105878 89944 105918 89984
rect 105960 89944 106000 89984
rect 120752 89944 120792 89984
rect 120834 89944 120874 89984
rect 120916 89944 120956 89984
rect 120998 89944 121038 89984
rect 121080 89944 121120 89984
rect 135872 89944 135912 89984
rect 135954 89944 135994 89984
rect 136036 89944 136076 89984
rect 136118 89944 136158 89984
rect 136200 89944 136240 89984
rect 150992 89944 151032 89984
rect 151074 89944 151114 89984
rect 151156 89944 151196 89984
rect 151238 89944 151278 89984
rect 151320 89944 151360 89984
rect 74152 89188 74192 89228
rect 74234 89188 74274 89228
rect 74316 89188 74356 89228
rect 74398 89188 74438 89228
rect 74480 89188 74520 89228
rect 89272 89188 89312 89228
rect 89354 89188 89394 89228
rect 89436 89188 89476 89228
rect 89518 89188 89558 89228
rect 89600 89188 89640 89228
rect 104392 89188 104432 89228
rect 104474 89188 104514 89228
rect 104556 89188 104596 89228
rect 104638 89188 104678 89228
rect 104720 89188 104760 89228
rect 119512 89188 119552 89228
rect 119594 89188 119634 89228
rect 119676 89188 119716 89228
rect 119758 89188 119798 89228
rect 119840 89188 119880 89228
rect 134632 89188 134672 89228
rect 134714 89188 134754 89228
rect 134796 89188 134836 89228
rect 134878 89188 134918 89228
rect 134960 89188 135000 89228
rect 149752 89188 149792 89228
rect 149834 89188 149874 89228
rect 149916 89188 149956 89228
rect 149998 89188 150038 89228
rect 150080 89188 150120 89228
rect 75392 88432 75432 88472
rect 75474 88432 75514 88472
rect 75556 88432 75596 88472
rect 75638 88432 75678 88472
rect 75720 88432 75760 88472
rect 90512 88432 90552 88472
rect 90594 88432 90634 88472
rect 90676 88432 90716 88472
rect 90758 88432 90798 88472
rect 90840 88432 90880 88472
rect 105632 88432 105672 88472
rect 105714 88432 105754 88472
rect 105796 88432 105836 88472
rect 105878 88432 105918 88472
rect 105960 88432 106000 88472
rect 120752 88432 120792 88472
rect 120834 88432 120874 88472
rect 120916 88432 120956 88472
rect 120998 88432 121038 88472
rect 121080 88432 121120 88472
rect 135872 88432 135912 88472
rect 135954 88432 135994 88472
rect 136036 88432 136076 88472
rect 136118 88432 136158 88472
rect 136200 88432 136240 88472
rect 150992 88432 151032 88472
rect 151074 88432 151114 88472
rect 151156 88432 151196 88472
rect 151238 88432 151278 88472
rect 151320 88432 151360 88472
rect 74152 87676 74192 87716
rect 74234 87676 74274 87716
rect 74316 87676 74356 87716
rect 74398 87676 74438 87716
rect 74480 87676 74520 87716
rect 89272 87676 89312 87716
rect 89354 87676 89394 87716
rect 89436 87676 89476 87716
rect 89518 87676 89558 87716
rect 89600 87676 89640 87716
rect 104392 87676 104432 87716
rect 104474 87676 104514 87716
rect 104556 87676 104596 87716
rect 104638 87676 104678 87716
rect 104720 87676 104760 87716
rect 119512 87676 119552 87716
rect 119594 87676 119634 87716
rect 119676 87676 119716 87716
rect 119758 87676 119798 87716
rect 119840 87676 119880 87716
rect 134632 87676 134672 87716
rect 134714 87676 134754 87716
rect 134796 87676 134836 87716
rect 134878 87676 134918 87716
rect 134960 87676 135000 87716
rect 149752 87676 149792 87716
rect 149834 87676 149874 87716
rect 149916 87676 149956 87716
rect 149998 87676 150038 87716
rect 150080 87676 150120 87716
rect 75392 86920 75432 86960
rect 75474 86920 75514 86960
rect 75556 86920 75596 86960
rect 75638 86920 75678 86960
rect 75720 86920 75760 86960
rect 90512 86920 90552 86960
rect 90594 86920 90634 86960
rect 90676 86920 90716 86960
rect 90758 86920 90798 86960
rect 90840 86920 90880 86960
rect 105632 86920 105672 86960
rect 105714 86920 105754 86960
rect 105796 86920 105836 86960
rect 105878 86920 105918 86960
rect 105960 86920 106000 86960
rect 120752 86920 120792 86960
rect 120834 86920 120874 86960
rect 120916 86920 120956 86960
rect 120998 86920 121038 86960
rect 121080 86920 121120 86960
rect 135872 86920 135912 86960
rect 135954 86920 135994 86960
rect 136036 86920 136076 86960
rect 136118 86920 136158 86960
rect 136200 86920 136240 86960
rect 150992 86920 151032 86960
rect 151074 86920 151114 86960
rect 151156 86920 151196 86960
rect 151238 86920 151278 86960
rect 151320 86920 151360 86960
rect 74152 86164 74192 86204
rect 74234 86164 74274 86204
rect 74316 86164 74356 86204
rect 74398 86164 74438 86204
rect 74480 86164 74520 86204
rect 89272 86164 89312 86204
rect 89354 86164 89394 86204
rect 89436 86164 89476 86204
rect 89518 86164 89558 86204
rect 89600 86164 89640 86204
rect 104392 86164 104432 86204
rect 104474 86164 104514 86204
rect 104556 86164 104596 86204
rect 104638 86164 104678 86204
rect 104720 86164 104760 86204
rect 119512 86164 119552 86204
rect 119594 86164 119634 86204
rect 119676 86164 119716 86204
rect 119758 86164 119798 86204
rect 119840 86164 119880 86204
rect 134632 86164 134672 86204
rect 134714 86164 134754 86204
rect 134796 86164 134836 86204
rect 134878 86164 134918 86204
rect 134960 86164 135000 86204
rect 149752 86164 149792 86204
rect 149834 86164 149874 86204
rect 149916 86164 149956 86204
rect 149998 86164 150038 86204
rect 150080 86164 150120 86204
rect 75392 85408 75432 85448
rect 75474 85408 75514 85448
rect 75556 85408 75596 85448
rect 75638 85408 75678 85448
rect 75720 85408 75760 85448
rect 90512 85408 90552 85448
rect 90594 85408 90634 85448
rect 90676 85408 90716 85448
rect 90758 85408 90798 85448
rect 90840 85408 90880 85448
rect 105632 85408 105672 85448
rect 105714 85408 105754 85448
rect 105796 85408 105836 85448
rect 105878 85408 105918 85448
rect 105960 85408 106000 85448
rect 120752 85408 120792 85448
rect 120834 85408 120874 85448
rect 120916 85408 120956 85448
rect 120998 85408 121038 85448
rect 121080 85408 121120 85448
rect 135872 85408 135912 85448
rect 135954 85408 135994 85448
rect 136036 85408 136076 85448
rect 136118 85408 136158 85448
rect 136200 85408 136240 85448
rect 150992 85408 151032 85448
rect 151074 85408 151114 85448
rect 151156 85408 151196 85448
rect 151238 85408 151278 85448
rect 151320 85408 151360 85448
rect 74152 84652 74192 84692
rect 74234 84652 74274 84692
rect 74316 84652 74356 84692
rect 74398 84652 74438 84692
rect 74480 84652 74520 84692
rect 89272 84652 89312 84692
rect 89354 84652 89394 84692
rect 89436 84652 89476 84692
rect 89518 84652 89558 84692
rect 89600 84652 89640 84692
rect 104392 84652 104432 84692
rect 104474 84652 104514 84692
rect 104556 84652 104596 84692
rect 104638 84652 104678 84692
rect 104720 84652 104760 84692
rect 119512 84652 119552 84692
rect 119594 84652 119634 84692
rect 119676 84652 119716 84692
rect 119758 84652 119798 84692
rect 119840 84652 119880 84692
rect 134632 84652 134672 84692
rect 134714 84652 134754 84692
rect 134796 84652 134836 84692
rect 134878 84652 134918 84692
rect 134960 84652 135000 84692
rect 149752 84652 149792 84692
rect 149834 84652 149874 84692
rect 149916 84652 149956 84692
rect 149998 84652 150038 84692
rect 150080 84652 150120 84692
rect 75392 83896 75432 83936
rect 75474 83896 75514 83936
rect 75556 83896 75596 83936
rect 75638 83896 75678 83936
rect 75720 83896 75760 83936
rect 90512 83896 90552 83936
rect 90594 83896 90634 83936
rect 90676 83896 90716 83936
rect 90758 83896 90798 83936
rect 90840 83896 90880 83936
rect 105632 83896 105672 83936
rect 105714 83896 105754 83936
rect 105796 83896 105836 83936
rect 105878 83896 105918 83936
rect 105960 83896 106000 83936
rect 120752 83896 120792 83936
rect 120834 83896 120874 83936
rect 120916 83896 120956 83936
rect 120998 83896 121038 83936
rect 121080 83896 121120 83936
rect 135872 83896 135912 83936
rect 135954 83896 135994 83936
rect 136036 83896 136076 83936
rect 136118 83896 136158 83936
rect 136200 83896 136240 83936
rect 150992 83896 151032 83936
rect 151074 83896 151114 83936
rect 151156 83896 151196 83936
rect 151238 83896 151278 83936
rect 151320 83896 151360 83936
rect 74152 83140 74192 83180
rect 74234 83140 74274 83180
rect 74316 83140 74356 83180
rect 74398 83140 74438 83180
rect 74480 83140 74520 83180
rect 89272 83140 89312 83180
rect 89354 83140 89394 83180
rect 89436 83140 89476 83180
rect 89518 83140 89558 83180
rect 89600 83140 89640 83180
rect 104392 83140 104432 83180
rect 104474 83140 104514 83180
rect 104556 83140 104596 83180
rect 104638 83140 104678 83180
rect 104720 83140 104760 83180
rect 119512 83140 119552 83180
rect 119594 83140 119634 83180
rect 119676 83140 119716 83180
rect 119758 83140 119798 83180
rect 119840 83140 119880 83180
rect 134632 83140 134672 83180
rect 134714 83140 134754 83180
rect 134796 83140 134836 83180
rect 134878 83140 134918 83180
rect 134960 83140 135000 83180
rect 149752 83140 149792 83180
rect 149834 83140 149874 83180
rect 149916 83140 149956 83180
rect 149998 83140 150038 83180
rect 150080 83140 150120 83180
rect 75392 82384 75432 82424
rect 75474 82384 75514 82424
rect 75556 82384 75596 82424
rect 75638 82384 75678 82424
rect 75720 82384 75760 82424
rect 90512 82384 90552 82424
rect 90594 82384 90634 82424
rect 90676 82384 90716 82424
rect 90758 82384 90798 82424
rect 90840 82384 90880 82424
rect 105632 82384 105672 82424
rect 105714 82384 105754 82424
rect 105796 82384 105836 82424
rect 105878 82384 105918 82424
rect 105960 82384 106000 82424
rect 120752 82384 120792 82424
rect 120834 82384 120874 82424
rect 120916 82384 120956 82424
rect 120998 82384 121038 82424
rect 121080 82384 121120 82424
rect 135872 82384 135912 82424
rect 135954 82384 135994 82424
rect 136036 82384 136076 82424
rect 136118 82384 136158 82424
rect 136200 82384 136240 82424
rect 150992 82384 151032 82424
rect 151074 82384 151114 82424
rect 151156 82384 151196 82424
rect 151238 82384 151278 82424
rect 151320 82384 151360 82424
rect 74152 81628 74192 81668
rect 74234 81628 74274 81668
rect 74316 81628 74356 81668
rect 74398 81628 74438 81668
rect 74480 81628 74520 81668
rect 89272 81628 89312 81668
rect 89354 81628 89394 81668
rect 89436 81628 89476 81668
rect 89518 81628 89558 81668
rect 89600 81628 89640 81668
rect 104392 81628 104432 81668
rect 104474 81628 104514 81668
rect 104556 81628 104596 81668
rect 104638 81628 104678 81668
rect 104720 81628 104760 81668
rect 119512 81628 119552 81668
rect 119594 81628 119634 81668
rect 119676 81628 119716 81668
rect 119758 81628 119798 81668
rect 119840 81628 119880 81668
rect 134632 81628 134672 81668
rect 134714 81628 134754 81668
rect 134796 81628 134836 81668
rect 134878 81628 134918 81668
rect 134960 81628 135000 81668
rect 149752 81628 149792 81668
rect 149834 81628 149874 81668
rect 149916 81628 149956 81668
rect 149998 81628 150038 81668
rect 150080 81628 150120 81668
rect 75392 80872 75432 80912
rect 75474 80872 75514 80912
rect 75556 80872 75596 80912
rect 75638 80872 75678 80912
rect 75720 80872 75760 80912
rect 90512 80872 90552 80912
rect 90594 80872 90634 80912
rect 90676 80872 90716 80912
rect 90758 80872 90798 80912
rect 90840 80872 90880 80912
rect 105632 80872 105672 80912
rect 105714 80872 105754 80912
rect 105796 80872 105836 80912
rect 105878 80872 105918 80912
rect 105960 80872 106000 80912
rect 120752 80872 120792 80912
rect 120834 80872 120874 80912
rect 120916 80872 120956 80912
rect 120998 80872 121038 80912
rect 121080 80872 121120 80912
rect 135872 80872 135912 80912
rect 135954 80872 135994 80912
rect 136036 80872 136076 80912
rect 136118 80872 136158 80912
rect 136200 80872 136240 80912
rect 150992 80872 151032 80912
rect 151074 80872 151114 80912
rect 151156 80872 151196 80912
rect 151238 80872 151278 80912
rect 151320 80872 151360 80912
rect 74152 80116 74192 80156
rect 74234 80116 74274 80156
rect 74316 80116 74356 80156
rect 74398 80116 74438 80156
rect 74480 80116 74520 80156
rect 89272 80116 89312 80156
rect 89354 80116 89394 80156
rect 89436 80116 89476 80156
rect 89518 80116 89558 80156
rect 89600 80116 89640 80156
rect 104392 80116 104432 80156
rect 104474 80116 104514 80156
rect 104556 80116 104596 80156
rect 104638 80116 104678 80156
rect 104720 80116 104760 80156
rect 119512 80116 119552 80156
rect 119594 80116 119634 80156
rect 119676 80116 119716 80156
rect 119758 80116 119798 80156
rect 119840 80116 119880 80156
rect 134632 80116 134672 80156
rect 134714 80116 134754 80156
rect 134796 80116 134836 80156
rect 134878 80116 134918 80156
rect 134960 80116 135000 80156
rect 149752 80116 149792 80156
rect 149834 80116 149874 80156
rect 149916 80116 149956 80156
rect 149998 80116 150038 80156
rect 150080 80116 150120 80156
rect 75392 79360 75432 79400
rect 75474 79360 75514 79400
rect 75556 79360 75596 79400
rect 75638 79360 75678 79400
rect 75720 79360 75760 79400
rect 90512 79360 90552 79400
rect 90594 79360 90634 79400
rect 90676 79360 90716 79400
rect 90758 79360 90798 79400
rect 90840 79360 90880 79400
rect 105632 79360 105672 79400
rect 105714 79360 105754 79400
rect 105796 79360 105836 79400
rect 105878 79360 105918 79400
rect 105960 79360 106000 79400
rect 120752 79360 120792 79400
rect 120834 79360 120874 79400
rect 120916 79360 120956 79400
rect 120998 79360 121038 79400
rect 121080 79360 121120 79400
rect 135872 79360 135912 79400
rect 135954 79360 135994 79400
rect 136036 79360 136076 79400
rect 136118 79360 136158 79400
rect 136200 79360 136240 79400
rect 150992 79360 151032 79400
rect 151074 79360 151114 79400
rect 151156 79360 151196 79400
rect 151238 79360 151278 79400
rect 151320 79360 151360 79400
rect 74152 78604 74192 78644
rect 74234 78604 74274 78644
rect 74316 78604 74356 78644
rect 74398 78604 74438 78644
rect 74480 78604 74520 78644
rect 89272 78604 89312 78644
rect 89354 78604 89394 78644
rect 89436 78604 89476 78644
rect 89518 78604 89558 78644
rect 89600 78604 89640 78644
rect 104392 78604 104432 78644
rect 104474 78604 104514 78644
rect 104556 78604 104596 78644
rect 104638 78604 104678 78644
rect 104720 78604 104760 78644
rect 119512 78604 119552 78644
rect 119594 78604 119634 78644
rect 119676 78604 119716 78644
rect 119758 78604 119798 78644
rect 119840 78604 119880 78644
rect 134632 78604 134672 78644
rect 134714 78604 134754 78644
rect 134796 78604 134836 78644
rect 134878 78604 134918 78644
rect 134960 78604 135000 78644
rect 149752 78604 149792 78644
rect 149834 78604 149874 78644
rect 149916 78604 149956 78644
rect 149998 78604 150038 78644
rect 150080 78604 150120 78644
rect 75392 77848 75432 77888
rect 75474 77848 75514 77888
rect 75556 77848 75596 77888
rect 75638 77848 75678 77888
rect 75720 77848 75760 77888
rect 90512 77848 90552 77888
rect 90594 77848 90634 77888
rect 90676 77848 90716 77888
rect 90758 77848 90798 77888
rect 90840 77848 90880 77888
rect 105632 77848 105672 77888
rect 105714 77848 105754 77888
rect 105796 77848 105836 77888
rect 105878 77848 105918 77888
rect 105960 77848 106000 77888
rect 120752 77848 120792 77888
rect 120834 77848 120874 77888
rect 120916 77848 120956 77888
rect 120998 77848 121038 77888
rect 121080 77848 121120 77888
rect 135872 77848 135912 77888
rect 135954 77848 135994 77888
rect 136036 77848 136076 77888
rect 136118 77848 136158 77888
rect 136200 77848 136240 77888
rect 150992 77848 151032 77888
rect 151074 77848 151114 77888
rect 151156 77848 151196 77888
rect 151238 77848 151278 77888
rect 151320 77848 151360 77888
rect 74152 77092 74192 77132
rect 74234 77092 74274 77132
rect 74316 77092 74356 77132
rect 74398 77092 74438 77132
rect 74480 77092 74520 77132
rect 89272 77092 89312 77132
rect 89354 77092 89394 77132
rect 89436 77092 89476 77132
rect 89518 77092 89558 77132
rect 89600 77092 89640 77132
rect 104392 77092 104432 77132
rect 104474 77092 104514 77132
rect 104556 77092 104596 77132
rect 104638 77092 104678 77132
rect 104720 77092 104760 77132
rect 119512 77092 119552 77132
rect 119594 77092 119634 77132
rect 119676 77092 119716 77132
rect 119758 77092 119798 77132
rect 119840 77092 119880 77132
rect 134632 77092 134672 77132
rect 134714 77092 134754 77132
rect 134796 77092 134836 77132
rect 134878 77092 134918 77132
rect 134960 77092 135000 77132
rect 149752 77092 149792 77132
rect 149834 77092 149874 77132
rect 149916 77092 149956 77132
rect 149998 77092 150038 77132
rect 150080 77092 150120 77132
rect 75392 76336 75432 76376
rect 75474 76336 75514 76376
rect 75556 76336 75596 76376
rect 75638 76336 75678 76376
rect 75720 76336 75760 76376
rect 90512 76336 90552 76376
rect 90594 76336 90634 76376
rect 90676 76336 90716 76376
rect 90758 76336 90798 76376
rect 90840 76336 90880 76376
rect 105632 76336 105672 76376
rect 105714 76336 105754 76376
rect 105796 76336 105836 76376
rect 105878 76336 105918 76376
rect 105960 76336 106000 76376
rect 120752 76336 120792 76376
rect 120834 76336 120874 76376
rect 120916 76336 120956 76376
rect 120998 76336 121038 76376
rect 121080 76336 121120 76376
rect 135872 76336 135912 76376
rect 135954 76336 135994 76376
rect 136036 76336 136076 76376
rect 136118 76336 136158 76376
rect 136200 76336 136240 76376
rect 150992 76336 151032 76376
rect 151074 76336 151114 76376
rect 151156 76336 151196 76376
rect 151238 76336 151278 76376
rect 151320 76336 151360 76376
rect 74152 75580 74192 75620
rect 74234 75580 74274 75620
rect 74316 75580 74356 75620
rect 74398 75580 74438 75620
rect 74480 75580 74520 75620
rect 89272 75580 89312 75620
rect 89354 75580 89394 75620
rect 89436 75580 89476 75620
rect 89518 75580 89558 75620
rect 89600 75580 89640 75620
rect 104392 75580 104432 75620
rect 104474 75580 104514 75620
rect 104556 75580 104596 75620
rect 104638 75580 104678 75620
rect 104720 75580 104760 75620
rect 119512 75580 119552 75620
rect 119594 75580 119634 75620
rect 119676 75580 119716 75620
rect 119758 75580 119798 75620
rect 119840 75580 119880 75620
rect 134632 75580 134672 75620
rect 134714 75580 134754 75620
rect 134796 75580 134836 75620
rect 134878 75580 134918 75620
rect 134960 75580 135000 75620
rect 149752 75580 149792 75620
rect 149834 75580 149874 75620
rect 149916 75580 149956 75620
rect 149998 75580 150038 75620
rect 150080 75580 150120 75620
rect 75392 74824 75432 74864
rect 75474 74824 75514 74864
rect 75556 74824 75596 74864
rect 75638 74824 75678 74864
rect 75720 74824 75760 74864
rect 90512 74824 90552 74864
rect 90594 74824 90634 74864
rect 90676 74824 90716 74864
rect 90758 74824 90798 74864
rect 90840 74824 90880 74864
rect 105632 74824 105672 74864
rect 105714 74824 105754 74864
rect 105796 74824 105836 74864
rect 105878 74824 105918 74864
rect 105960 74824 106000 74864
rect 120752 74824 120792 74864
rect 120834 74824 120874 74864
rect 120916 74824 120956 74864
rect 120998 74824 121038 74864
rect 121080 74824 121120 74864
rect 135872 74824 135912 74864
rect 135954 74824 135994 74864
rect 136036 74824 136076 74864
rect 136118 74824 136158 74864
rect 136200 74824 136240 74864
rect 150992 74824 151032 74864
rect 151074 74824 151114 74864
rect 151156 74824 151196 74864
rect 151238 74824 151278 74864
rect 151320 74824 151360 74864
rect 74152 74068 74192 74108
rect 74234 74068 74274 74108
rect 74316 74068 74356 74108
rect 74398 74068 74438 74108
rect 74480 74068 74520 74108
rect 89272 74068 89312 74108
rect 89354 74068 89394 74108
rect 89436 74068 89476 74108
rect 89518 74068 89558 74108
rect 89600 74068 89640 74108
rect 104392 74068 104432 74108
rect 104474 74068 104514 74108
rect 104556 74068 104596 74108
rect 104638 74068 104678 74108
rect 104720 74068 104760 74108
rect 119512 74068 119552 74108
rect 119594 74068 119634 74108
rect 119676 74068 119716 74108
rect 119758 74068 119798 74108
rect 119840 74068 119880 74108
rect 134632 74068 134672 74108
rect 134714 74068 134754 74108
rect 134796 74068 134836 74108
rect 134878 74068 134918 74108
rect 134960 74068 135000 74108
rect 149752 74068 149792 74108
rect 149834 74068 149874 74108
rect 149916 74068 149956 74108
rect 149998 74068 150038 74108
rect 150080 74068 150120 74108
rect 75392 73312 75432 73352
rect 75474 73312 75514 73352
rect 75556 73312 75596 73352
rect 75638 73312 75678 73352
rect 75720 73312 75760 73352
rect 90512 73312 90552 73352
rect 90594 73312 90634 73352
rect 90676 73312 90716 73352
rect 90758 73312 90798 73352
rect 90840 73312 90880 73352
rect 105632 73312 105672 73352
rect 105714 73312 105754 73352
rect 105796 73312 105836 73352
rect 105878 73312 105918 73352
rect 105960 73312 106000 73352
rect 120752 73312 120792 73352
rect 120834 73312 120874 73352
rect 120916 73312 120956 73352
rect 120998 73312 121038 73352
rect 121080 73312 121120 73352
rect 135872 73312 135912 73352
rect 135954 73312 135994 73352
rect 136036 73312 136076 73352
rect 136118 73312 136158 73352
rect 136200 73312 136240 73352
rect 150992 73312 151032 73352
rect 151074 73312 151114 73352
rect 151156 73312 151196 73352
rect 151238 73312 151278 73352
rect 151320 73312 151360 73352
rect 74152 72556 74192 72596
rect 74234 72556 74274 72596
rect 74316 72556 74356 72596
rect 74398 72556 74438 72596
rect 74480 72556 74520 72596
rect 89272 72556 89312 72596
rect 89354 72556 89394 72596
rect 89436 72556 89476 72596
rect 89518 72556 89558 72596
rect 89600 72556 89640 72596
rect 104392 72556 104432 72596
rect 104474 72556 104514 72596
rect 104556 72556 104596 72596
rect 104638 72556 104678 72596
rect 104720 72556 104760 72596
rect 119512 72556 119552 72596
rect 119594 72556 119634 72596
rect 119676 72556 119716 72596
rect 119758 72556 119798 72596
rect 119840 72556 119880 72596
rect 134632 72556 134672 72596
rect 134714 72556 134754 72596
rect 134796 72556 134836 72596
rect 134878 72556 134918 72596
rect 134960 72556 135000 72596
rect 149752 72556 149792 72596
rect 149834 72556 149874 72596
rect 149916 72556 149956 72596
rect 149998 72556 150038 72596
rect 150080 72556 150120 72596
rect 75392 71800 75432 71840
rect 75474 71800 75514 71840
rect 75556 71800 75596 71840
rect 75638 71800 75678 71840
rect 75720 71800 75760 71840
rect 90512 71800 90552 71840
rect 90594 71800 90634 71840
rect 90676 71800 90716 71840
rect 90758 71800 90798 71840
rect 90840 71800 90880 71840
rect 105632 71800 105672 71840
rect 105714 71800 105754 71840
rect 105796 71800 105836 71840
rect 105878 71800 105918 71840
rect 105960 71800 106000 71840
rect 120752 71800 120792 71840
rect 120834 71800 120874 71840
rect 120916 71800 120956 71840
rect 120998 71800 121038 71840
rect 121080 71800 121120 71840
rect 135872 71800 135912 71840
rect 135954 71800 135994 71840
rect 136036 71800 136076 71840
rect 136118 71800 136158 71840
rect 136200 71800 136240 71840
rect 150992 71800 151032 71840
rect 151074 71800 151114 71840
rect 151156 71800 151196 71840
rect 151238 71800 151278 71840
rect 151320 71800 151360 71840
<< metal5 >>
rect 75383 151999 75769 152018
rect 75383 151976 75449 151999
rect 75535 151976 75617 151999
rect 75703 151976 75769 151999
rect 75383 151936 75392 151976
rect 75432 151936 75449 151976
rect 75535 151936 75556 151976
rect 75596 151936 75617 151976
rect 75703 151936 75720 151976
rect 75760 151936 75769 151976
rect 75383 151913 75449 151936
rect 75535 151913 75617 151936
rect 75703 151913 75769 151936
rect 75383 151894 75769 151913
rect 90503 151999 90889 152018
rect 90503 151976 90569 151999
rect 90655 151976 90737 151999
rect 90823 151976 90889 151999
rect 90503 151936 90512 151976
rect 90552 151936 90569 151976
rect 90655 151936 90676 151976
rect 90716 151936 90737 151976
rect 90823 151936 90840 151976
rect 90880 151936 90889 151976
rect 90503 151913 90569 151936
rect 90655 151913 90737 151936
rect 90823 151913 90889 151936
rect 90503 151894 90889 151913
rect 105623 151999 106009 152018
rect 105623 151976 105689 151999
rect 105775 151976 105857 151999
rect 105943 151976 106009 151999
rect 105623 151936 105632 151976
rect 105672 151936 105689 151976
rect 105775 151936 105796 151976
rect 105836 151936 105857 151976
rect 105943 151936 105960 151976
rect 106000 151936 106009 151976
rect 105623 151913 105689 151936
rect 105775 151913 105857 151936
rect 105943 151913 106009 151936
rect 105623 151894 106009 151913
rect 120743 151999 121129 152018
rect 120743 151976 120809 151999
rect 120895 151976 120977 151999
rect 121063 151976 121129 151999
rect 120743 151936 120752 151976
rect 120792 151936 120809 151976
rect 120895 151936 120916 151976
rect 120956 151936 120977 151976
rect 121063 151936 121080 151976
rect 121120 151936 121129 151976
rect 120743 151913 120809 151936
rect 120895 151913 120977 151936
rect 121063 151913 121129 151936
rect 120743 151894 121129 151913
rect 135863 151999 136249 152018
rect 135863 151976 135929 151999
rect 136015 151976 136097 151999
rect 136183 151976 136249 151999
rect 135863 151936 135872 151976
rect 135912 151936 135929 151976
rect 136015 151936 136036 151976
rect 136076 151936 136097 151976
rect 136183 151936 136200 151976
rect 136240 151936 136249 151976
rect 135863 151913 135929 151936
rect 136015 151913 136097 151936
rect 136183 151913 136249 151936
rect 135863 151894 136249 151913
rect 150983 151999 151369 152018
rect 150983 151976 151049 151999
rect 151135 151976 151217 151999
rect 151303 151976 151369 151999
rect 150983 151936 150992 151976
rect 151032 151936 151049 151976
rect 151135 151936 151156 151976
rect 151196 151936 151217 151976
rect 151303 151936 151320 151976
rect 151360 151936 151369 151976
rect 150983 151913 151049 151936
rect 151135 151913 151217 151936
rect 151303 151913 151369 151936
rect 150983 151894 151369 151913
rect 74143 151243 74529 151262
rect 74143 151220 74209 151243
rect 74295 151220 74377 151243
rect 74463 151220 74529 151243
rect 74143 151180 74152 151220
rect 74192 151180 74209 151220
rect 74295 151180 74316 151220
rect 74356 151180 74377 151220
rect 74463 151180 74480 151220
rect 74520 151180 74529 151220
rect 74143 151157 74209 151180
rect 74295 151157 74377 151180
rect 74463 151157 74529 151180
rect 74143 151138 74529 151157
rect 89263 151243 89649 151262
rect 89263 151220 89329 151243
rect 89415 151220 89497 151243
rect 89583 151220 89649 151243
rect 89263 151180 89272 151220
rect 89312 151180 89329 151220
rect 89415 151180 89436 151220
rect 89476 151180 89497 151220
rect 89583 151180 89600 151220
rect 89640 151180 89649 151220
rect 89263 151157 89329 151180
rect 89415 151157 89497 151180
rect 89583 151157 89649 151180
rect 89263 151138 89649 151157
rect 104383 151243 104769 151262
rect 104383 151220 104449 151243
rect 104535 151220 104617 151243
rect 104703 151220 104769 151243
rect 104383 151180 104392 151220
rect 104432 151180 104449 151220
rect 104535 151180 104556 151220
rect 104596 151180 104617 151220
rect 104703 151180 104720 151220
rect 104760 151180 104769 151220
rect 104383 151157 104449 151180
rect 104535 151157 104617 151180
rect 104703 151157 104769 151180
rect 104383 151138 104769 151157
rect 119503 151243 119889 151262
rect 119503 151220 119569 151243
rect 119655 151220 119737 151243
rect 119823 151220 119889 151243
rect 119503 151180 119512 151220
rect 119552 151180 119569 151220
rect 119655 151180 119676 151220
rect 119716 151180 119737 151220
rect 119823 151180 119840 151220
rect 119880 151180 119889 151220
rect 119503 151157 119569 151180
rect 119655 151157 119737 151180
rect 119823 151157 119889 151180
rect 119503 151138 119889 151157
rect 134623 151243 135009 151262
rect 134623 151220 134689 151243
rect 134775 151220 134857 151243
rect 134943 151220 135009 151243
rect 134623 151180 134632 151220
rect 134672 151180 134689 151220
rect 134775 151180 134796 151220
rect 134836 151180 134857 151220
rect 134943 151180 134960 151220
rect 135000 151180 135009 151220
rect 134623 151157 134689 151180
rect 134775 151157 134857 151180
rect 134943 151157 135009 151180
rect 134623 151138 135009 151157
rect 149743 151243 150129 151262
rect 149743 151220 149809 151243
rect 149895 151220 149977 151243
rect 150063 151220 150129 151243
rect 149743 151180 149752 151220
rect 149792 151180 149809 151220
rect 149895 151180 149916 151220
rect 149956 151180 149977 151220
rect 150063 151180 150080 151220
rect 150120 151180 150129 151220
rect 149743 151157 149809 151180
rect 149895 151157 149977 151180
rect 150063 151157 150129 151180
rect 149743 151138 150129 151157
rect 75383 150487 75769 150506
rect 75383 150464 75449 150487
rect 75535 150464 75617 150487
rect 75703 150464 75769 150487
rect 75383 150424 75392 150464
rect 75432 150424 75449 150464
rect 75535 150424 75556 150464
rect 75596 150424 75617 150464
rect 75703 150424 75720 150464
rect 75760 150424 75769 150464
rect 75383 150401 75449 150424
rect 75535 150401 75617 150424
rect 75703 150401 75769 150424
rect 75383 150382 75769 150401
rect 90503 150487 90889 150506
rect 90503 150464 90569 150487
rect 90655 150464 90737 150487
rect 90823 150464 90889 150487
rect 90503 150424 90512 150464
rect 90552 150424 90569 150464
rect 90655 150424 90676 150464
rect 90716 150424 90737 150464
rect 90823 150424 90840 150464
rect 90880 150424 90889 150464
rect 90503 150401 90569 150424
rect 90655 150401 90737 150424
rect 90823 150401 90889 150424
rect 90503 150382 90889 150401
rect 105623 150487 106009 150506
rect 105623 150464 105689 150487
rect 105775 150464 105857 150487
rect 105943 150464 106009 150487
rect 105623 150424 105632 150464
rect 105672 150424 105689 150464
rect 105775 150424 105796 150464
rect 105836 150424 105857 150464
rect 105943 150424 105960 150464
rect 106000 150424 106009 150464
rect 105623 150401 105689 150424
rect 105775 150401 105857 150424
rect 105943 150401 106009 150424
rect 105623 150382 106009 150401
rect 120743 150487 121129 150506
rect 120743 150464 120809 150487
rect 120895 150464 120977 150487
rect 121063 150464 121129 150487
rect 120743 150424 120752 150464
rect 120792 150424 120809 150464
rect 120895 150424 120916 150464
rect 120956 150424 120977 150464
rect 121063 150424 121080 150464
rect 121120 150424 121129 150464
rect 120743 150401 120809 150424
rect 120895 150401 120977 150424
rect 121063 150401 121129 150424
rect 120743 150382 121129 150401
rect 135863 150487 136249 150506
rect 135863 150464 135929 150487
rect 136015 150464 136097 150487
rect 136183 150464 136249 150487
rect 135863 150424 135872 150464
rect 135912 150424 135929 150464
rect 136015 150424 136036 150464
rect 136076 150424 136097 150464
rect 136183 150424 136200 150464
rect 136240 150424 136249 150464
rect 135863 150401 135929 150424
rect 136015 150401 136097 150424
rect 136183 150401 136249 150424
rect 135863 150382 136249 150401
rect 150983 150487 151369 150506
rect 150983 150464 151049 150487
rect 151135 150464 151217 150487
rect 151303 150464 151369 150487
rect 150983 150424 150992 150464
rect 151032 150424 151049 150464
rect 151135 150424 151156 150464
rect 151196 150424 151217 150464
rect 151303 150424 151320 150464
rect 151360 150424 151369 150464
rect 150983 150401 151049 150424
rect 151135 150401 151217 150424
rect 151303 150401 151369 150424
rect 150983 150382 151369 150401
rect 74143 149731 74529 149750
rect 74143 149708 74209 149731
rect 74295 149708 74377 149731
rect 74463 149708 74529 149731
rect 74143 149668 74152 149708
rect 74192 149668 74209 149708
rect 74295 149668 74316 149708
rect 74356 149668 74377 149708
rect 74463 149668 74480 149708
rect 74520 149668 74529 149708
rect 74143 149645 74209 149668
rect 74295 149645 74377 149668
rect 74463 149645 74529 149668
rect 74143 149626 74529 149645
rect 89263 149731 89649 149750
rect 89263 149708 89329 149731
rect 89415 149708 89497 149731
rect 89583 149708 89649 149731
rect 89263 149668 89272 149708
rect 89312 149668 89329 149708
rect 89415 149668 89436 149708
rect 89476 149668 89497 149708
rect 89583 149668 89600 149708
rect 89640 149668 89649 149708
rect 89263 149645 89329 149668
rect 89415 149645 89497 149668
rect 89583 149645 89649 149668
rect 89263 149626 89649 149645
rect 104383 149731 104769 149750
rect 104383 149708 104449 149731
rect 104535 149708 104617 149731
rect 104703 149708 104769 149731
rect 104383 149668 104392 149708
rect 104432 149668 104449 149708
rect 104535 149668 104556 149708
rect 104596 149668 104617 149708
rect 104703 149668 104720 149708
rect 104760 149668 104769 149708
rect 104383 149645 104449 149668
rect 104535 149645 104617 149668
rect 104703 149645 104769 149668
rect 104383 149626 104769 149645
rect 119503 149731 119889 149750
rect 119503 149708 119569 149731
rect 119655 149708 119737 149731
rect 119823 149708 119889 149731
rect 119503 149668 119512 149708
rect 119552 149668 119569 149708
rect 119655 149668 119676 149708
rect 119716 149668 119737 149708
rect 119823 149668 119840 149708
rect 119880 149668 119889 149708
rect 119503 149645 119569 149668
rect 119655 149645 119737 149668
rect 119823 149645 119889 149668
rect 119503 149626 119889 149645
rect 134623 149731 135009 149750
rect 134623 149708 134689 149731
rect 134775 149708 134857 149731
rect 134943 149708 135009 149731
rect 134623 149668 134632 149708
rect 134672 149668 134689 149708
rect 134775 149668 134796 149708
rect 134836 149668 134857 149708
rect 134943 149668 134960 149708
rect 135000 149668 135009 149708
rect 134623 149645 134689 149668
rect 134775 149645 134857 149668
rect 134943 149645 135009 149668
rect 134623 149626 135009 149645
rect 149743 149731 150129 149750
rect 149743 149708 149809 149731
rect 149895 149708 149977 149731
rect 150063 149708 150129 149731
rect 149743 149668 149752 149708
rect 149792 149668 149809 149708
rect 149895 149668 149916 149708
rect 149956 149668 149977 149708
rect 150063 149668 150080 149708
rect 150120 149668 150129 149708
rect 149743 149645 149809 149668
rect 149895 149645 149977 149668
rect 150063 149645 150129 149668
rect 149743 149626 150129 149645
rect 75383 148975 75769 148994
rect 75383 148952 75449 148975
rect 75535 148952 75617 148975
rect 75703 148952 75769 148975
rect 75383 148912 75392 148952
rect 75432 148912 75449 148952
rect 75535 148912 75556 148952
rect 75596 148912 75617 148952
rect 75703 148912 75720 148952
rect 75760 148912 75769 148952
rect 75383 148889 75449 148912
rect 75535 148889 75617 148912
rect 75703 148889 75769 148912
rect 75383 148870 75769 148889
rect 90503 148975 90889 148994
rect 90503 148952 90569 148975
rect 90655 148952 90737 148975
rect 90823 148952 90889 148975
rect 90503 148912 90512 148952
rect 90552 148912 90569 148952
rect 90655 148912 90676 148952
rect 90716 148912 90737 148952
rect 90823 148912 90840 148952
rect 90880 148912 90889 148952
rect 90503 148889 90569 148912
rect 90655 148889 90737 148912
rect 90823 148889 90889 148912
rect 90503 148870 90889 148889
rect 105623 148975 106009 148994
rect 105623 148952 105689 148975
rect 105775 148952 105857 148975
rect 105943 148952 106009 148975
rect 105623 148912 105632 148952
rect 105672 148912 105689 148952
rect 105775 148912 105796 148952
rect 105836 148912 105857 148952
rect 105943 148912 105960 148952
rect 106000 148912 106009 148952
rect 105623 148889 105689 148912
rect 105775 148889 105857 148912
rect 105943 148889 106009 148912
rect 105623 148870 106009 148889
rect 120743 148975 121129 148994
rect 120743 148952 120809 148975
rect 120895 148952 120977 148975
rect 121063 148952 121129 148975
rect 120743 148912 120752 148952
rect 120792 148912 120809 148952
rect 120895 148912 120916 148952
rect 120956 148912 120977 148952
rect 121063 148912 121080 148952
rect 121120 148912 121129 148952
rect 120743 148889 120809 148912
rect 120895 148889 120977 148912
rect 121063 148889 121129 148912
rect 120743 148870 121129 148889
rect 135863 148975 136249 148994
rect 135863 148952 135929 148975
rect 136015 148952 136097 148975
rect 136183 148952 136249 148975
rect 135863 148912 135872 148952
rect 135912 148912 135929 148952
rect 136015 148912 136036 148952
rect 136076 148912 136097 148952
rect 136183 148912 136200 148952
rect 136240 148912 136249 148952
rect 135863 148889 135929 148912
rect 136015 148889 136097 148912
rect 136183 148889 136249 148912
rect 135863 148870 136249 148889
rect 150983 148975 151369 148994
rect 150983 148952 151049 148975
rect 151135 148952 151217 148975
rect 151303 148952 151369 148975
rect 150983 148912 150992 148952
rect 151032 148912 151049 148952
rect 151135 148912 151156 148952
rect 151196 148912 151217 148952
rect 151303 148912 151320 148952
rect 151360 148912 151369 148952
rect 150983 148889 151049 148912
rect 151135 148889 151217 148912
rect 151303 148889 151369 148912
rect 150983 148870 151369 148889
rect 74143 148219 74529 148238
rect 74143 148196 74209 148219
rect 74295 148196 74377 148219
rect 74463 148196 74529 148219
rect 74143 148156 74152 148196
rect 74192 148156 74209 148196
rect 74295 148156 74316 148196
rect 74356 148156 74377 148196
rect 74463 148156 74480 148196
rect 74520 148156 74529 148196
rect 74143 148133 74209 148156
rect 74295 148133 74377 148156
rect 74463 148133 74529 148156
rect 74143 148114 74529 148133
rect 89263 148219 89649 148238
rect 89263 148196 89329 148219
rect 89415 148196 89497 148219
rect 89583 148196 89649 148219
rect 89263 148156 89272 148196
rect 89312 148156 89329 148196
rect 89415 148156 89436 148196
rect 89476 148156 89497 148196
rect 89583 148156 89600 148196
rect 89640 148156 89649 148196
rect 89263 148133 89329 148156
rect 89415 148133 89497 148156
rect 89583 148133 89649 148156
rect 89263 148114 89649 148133
rect 104383 148219 104769 148238
rect 104383 148196 104449 148219
rect 104535 148196 104617 148219
rect 104703 148196 104769 148219
rect 104383 148156 104392 148196
rect 104432 148156 104449 148196
rect 104535 148156 104556 148196
rect 104596 148156 104617 148196
rect 104703 148156 104720 148196
rect 104760 148156 104769 148196
rect 104383 148133 104449 148156
rect 104535 148133 104617 148156
rect 104703 148133 104769 148156
rect 104383 148114 104769 148133
rect 119503 148219 119889 148238
rect 119503 148196 119569 148219
rect 119655 148196 119737 148219
rect 119823 148196 119889 148219
rect 119503 148156 119512 148196
rect 119552 148156 119569 148196
rect 119655 148156 119676 148196
rect 119716 148156 119737 148196
rect 119823 148156 119840 148196
rect 119880 148156 119889 148196
rect 119503 148133 119569 148156
rect 119655 148133 119737 148156
rect 119823 148133 119889 148156
rect 119503 148114 119889 148133
rect 134623 148219 135009 148238
rect 134623 148196 134689 148219
rect 134775 148196 134857 148219
rect 134943 148196 135009 148219
rect 134623 148156 134632 148196
rect 134672 148156 134689 148196
rect 134775 148156 134796 148196
rect 134836 148156 134857 148196
rect 134943 148156 134960 148196
rect 135000 148156 135009 148196
rect 134623 148133 134689 148156
rect 134775 148133 134857 148156
rect 134943 148133 135009 148156
rect 134623 148114 135009 148133
rect 149743 148219 150129 148238
rect 149743 148196 149809 148219
rect 149895 148196 149977 148219
rect 150063 148196 150129 148219
rect 149743 148156 149752 148196
rect 149792 148156 149809 148196
rect 149895 148156 149916 148196
rect 149956 148156 149977 148196
rect 150063 148156 150080 148196
rect 150120 148156 150129 148196
rect 149743 148133 149809 148156
rect 149895 148133 149977 148156
rect 150063 148133 150129 148156
rect 149743 148114 150129 148133
rect 75383 147463 75769 147482
rect 75383 147440 75449 147463
rect 75535 147440 75617 147463
rect 75703 147440 75769 147463
rect 75383 147400 75392 147440
rect 75432 147400 75449 147440
rect 75535 147400 75556 147440
rect 75596 147400 75617 147440
rect 75703 147400 75720 147440
rect 75760 147400 75769 147440
rect 75383 147377 75449 147400
rect 75535 147377 75617 147400
rect 75703 147377 75769 147400
rect 75383 147358 75769 147377
rect 90503 147463 90889 147482
rect 90503 147440 90569 147463
rect 90655 147440 90737 147463
rect 90823 147440 90889 147463
rect 90503 147400 90512 147440
rect 90552 147400 90569 147440
rect 90655 147400 90676 147440
rect 90716 147400 90737 147440
rect 90823 147400 90840 147440
rect 90880 147400 90889 147440
rect 90503 147377 90569 147400
rect 90655 147377 90737 147400
rect 90823 147377 90889 147400
rect 90503 147358 90889 147377
rect 105623 147463 106009 147482
rect 105623 147440 105689 147463
rect 105775 147440 105857 147463
rect 105943 147440 106009 147463
rect 105623 147400 105632 147440
rect 105672 147400 105689 147440
rect 105775 147400 105796 147440
rect 105836 147400 105857 147440
rect 105943 147400 105960 147440
rect 106000 147400 106009 147440
rect 105623 147377 105689 147400
rect 105775 147377 105857 147400
rect 105943 147377 106009 147400
rect 105623 147358 106009 147377
rect 120743 147463 121129 147482
rect 120743 147440 120809 147463
rect 120895 147440 120977 147463
rect 121063 147440 121129 147463
rect 120743 147400 120752 147440
rect 120792 147400 120809 147440
rect 120895 147400 120916 147440
rect 120956 147400 120977 147440
rect 121063 147400 121080 147440
rect 121120 147400 121129 147440
rect 120743 147377 120809 147400
rect 120895 147377 120977 147400
rect 121063 147377 121129 147400
rect 120743 147358 121129 147377
rect 135863 147463 136249 147482
rect 135863 147440 135929 147463
rect 136015 147440 136097 147463
rect 136183 147440 136249 147463
rect 135863 147400 135872 147440
rect 135912 147400 135929 147440
rect 136015 147400 136036 147440
rect 136076 147400 136097 147440
rect 136183 147400 136200 147440
rect 136240 147400 136249 147440
rect 135863 147377 135929 147400
rect 136015 147377 136097 147400
rect 136183 147377 136249 147400
rect 135863 147358 136249 147377
rect 150983 147463 151369 147482
rect 150983 147440 151049 147463
rect 151135 147440 151217 147463
rect 151303 147440 151369 147463
rect 150983 147400 150992 147440
rect 151032 147400 151049 147440
rect 151135 147400 151156 147440
rect 151196 147400 151217 147440
rect 151303 147400 151320 147440
rect 151360 147400 151369 147440
rect 150983 147377 151049 147400
rect 151135 147377 151217 147400
rect 151303 147377 151369 147400
rect 150983 147358 151369 147377
rect 74143 146707 74529 146726
rect 74143 146684 74209 146707
rect 74295 146684 74377 146707
rect 74463 146684 74529 146707
rect 74143 146644 74152 146684
rect 74192 146644 74209 146684
rect 74295 146644 74316 146684
rect 74356 146644 74377 146684
rect 74463 146644 74480 146684
rect 74520 146644 74529 146684
rect 74143 146621 74209 146644
rect 74295 146621 74377 146644
rect 74463 146621 74529 146644
rect 74143 146602 74529 146621
rect 89263 146707 89649 146726
rect 89263 146684 89329 146707
rect 89415 146684 89497 146707
rect 89583 146684 89649 146707
rect 89263 146644 89272 146684
rect 89312 146644 89329 146684
rect 89415 146644 89436 146684
rect 89476 146644 89497 146684
rect 89583 146644 89600 146684
rect 89640 146644 89649 146684
rect 89263 146621 89329 146644
rect 89415 146621 89497 146644
rect 89583 146621 89649 146644
rect 89263 146602 89649 146621
rect 104383 146707 104769 146726
rect 104383 146684 104449 146707
rect 104535 146684 104617 146707
rect 104703 146684 104769 146707
rect 104383 146644 104392 146684
rect 104432 146644 104449 146684
rect 104535 146644 104556 146684
rect 104596 146644 104617 146684
rect 104703 146644 104720 146684
rect 104760 146644 104769 146684
rect 104383 146621 104449 146644
rect 104535 146621 104617 146644
rect 104703 146621 104769 146644
rect 104383 146602 104769 146621
rect 119503 146707 119889 146726
rect 119503 146684 119569 146707
rect 119655 146684 119737 146707
rect 119823 146684 119889 146707
rect 119503 146644 119512 146684
rect 119552 146644 119569 146684
rect 119655 146644 119676 146684
rect 119716 146644 119737 146684
rect 119823 146644 119840 146684
rect 119880 146644 119889 146684
rect 119503 146621 119569 146644
rect 119655 146621 119737 146644
rect 119823 146621 119889 146644
rect 119503 146602 119889 146621
rect 134623 146707 135009 146726
rect 134623 146684 134689 146707
rect 134775 146684 134857 146707
rect 134943 146684 135009 146707
rect 134623 146644 134632 146684
rect 134672 146644 134689 146684
rect 134775 146644 134796 146684
rect 134836 146644 134857 146684
rect 134943 146644 134960 146684
rect 135000 146644 135009 146684
rect 134623 146621 134689 146644
rect 134775 146621 134857 146644
rect 134943 146621 135009 146644
rect 134623 146602 135009 146621
rect 149743 146707 150129 146726
rect 149743 146684 149809 146707
rect 149895 146684 149977 146707
rect 150063 146684 150129 146707
rect 149743 146644 149752 146684
rect 149792 146644 149809 146684
rect 149895 146644 149916 146684
rect 149956 146644 149977 146684
rect 150063 146644 150080 146684
rect 150120 146644 150129 146684
rect 149743 146621 149809 146644
rect 149895 146621 149977 146644
rect 150063 146621 150129 146644
rect 149743 146602 150129 146621
rect 75383 145951 75769 145970
rect 75383 145928 75449 145951
rect 75535 145928 75617 145951
rect 75703 145928 75769 145951
rect 75383 145888 75392 145928
rect 75432 145888 75449 145928
rect 75535 145888 75556 145928
rect 75596 145888 75617 145928
rect 75703 145888 75720 145928
rect 75760 145888 75769 145928
rect 75383 145865 75449 145888
rect 75535 145865 75617 145888
rect 75703 145865 75769 145888
rect 75383 145846 75769 145865
rect 90503 145951 90889 145970
rect 90503 145928 90569 145951
rect 90655 145928 90737 145951
rect 90823 145928 90889 145951
rect 90503 145888 90512 145928
rect 90552 145888 90569 145928
rect 90655 145888 90676 145928
rect 90716 145888 90737 145928
rect 90823 145888 90840 145928
rect 90880 145888 90889 145928
rect 90503 145865 90569 145888
rect 90655 145865 90737 145888
rect 90823 145865 90889 145888
rect 90503 145846 90889 145865
rect 105623 145951 106009 145970
rect 105623 145928 105689 145951
rect 105775 145928 105857 145951
rect 105943 145928 106009 145951
rect 105623 145888 105632 145928
rect 105672 145888 105689 145928
rect 105775 145888 105796 145928
rect 105836 145888 105857 145928
rect 105943 145888 105960 145928
rect 106000 145888 106009 145928
rect 105623 145865 105689 145888
rect 105775 145865 105857 145888
rect 105943 145865 106009 145888
rect 105623 145846 106009 145865
rect 120743 145951 121129 145970
rect 120743 145928 120809 145951
rect 120895 145928 120977 145951
rect 121063 145928 121129 145951
rect 120743 145888 120752 145928
rect 120792 145888 120809 145928
rect 120895 145888 120916 145928
rect 120956 145888 120977 145928
rect 121063 145888 121080 145928
rect 121120 145888 121129 145928
rect 120743 145865 120809 145888
rect 120895 145865 120977 145888
rect 121063 145865 121129 145888
rect 120743 145846 121129 145865
rect 135863 145951 136249 145970
rect 135863 145928 135929 145951
rect 136015 145928 136097 145951
rect 136183 145928 136249 145951
rect 135863 145888 135872 145928
rect 135912 145888 135929 145928
rect 136015 145888 136036 145928
rect 136076 145888 136097 145928
rect 136183 145888 136200 145928
rect 136240 145888 136249 145928
rect 135863 145865 135929 145888
rect 136015 145865 136097 145888
rect 136183 145865 136249 145888
rect 135863 145846 136249 145865
rect 150983 145951 151369 145970
rect 150983 145928 151049 145951
rect 151135 145928 151217 145951
rect 151303 145928 151369 145951
rect 150983 145888 150992 145928
rect 151032 145888 151049 145928
rect 151135 145888 151156 145928
rect 151196 145888 151217 145928
rect 151303 145888 151320 145928
rect 151360 145888 151369 145928
rect 150983 145865 151049 145888
rect 151135 145865 151217 145888
rect 151303 145865 151369 145888
rect 150983 145846 151369 145865
rect 74143 145195 74529 145214
rect 74143 145172 74209 145195
rect 74295 145172 74377 145195
rect 74463 145172 74529 145195
rect 74143 145132 74152 145172
rect 74192 145132 74209 145172
rect 74295 145132 74316 145172
rect 74356 145132 74377 145172
rect 74463 145132 74480 145172
rect 74520 145132 74529 145172
rect 74143 145109 74209 145132
rect 74295 145109 74377 145132
rect 74463 145109 74529 145132
rect 74143 145090 74529 145109
rect 89263 145195 89649 145214
rect 89263 145172 89329 145195
rect 89415 145172 89497 145195
rect 89583 145172 89649 145195
rect 89263 145132 89272 145172
rect 89312 145132 89329 145172
rect 89415 145132 89436 145172
rect 89476 145132 89497 145172
rect 89583 145132 89600 145172
rect 89640 145132 89649 145172
rect 89263 145109 89329 145132
rect 89415 145109 89497 145132
rect 89583 145109 89649 145132
rect 89263 145090 89649 145109
rect 104383 145195 104769 145214
rect 104383 145172 104449 145195
rect 104535 145172 104617 145195
rect 104703 145172 104769 145195
rect 104383 145132 104392 145172
rect 104432 145132 104449 145172
rect 104535 145132 104556 145172
rect 104596 145132 104617 145172
rect 104703 145132 104720 145172
rect 104760 145132 104769 145172
rect 104383 145109 104449 145132
rect 104535 145109 104617 145132
rect 104703 145109 104769 145132
rect 104383 145090 104769 145109
rect 119503 145195 119889 145214
rect 119503 145172 119569 145195
rect 119655 145172 119737 145195
rect 119823 145172 119889 145195
rect 119503 145132 119512 145172
rect 119552 145132 119569 145172
rect 119655 145132 119676 145172
rect 119716 145132 119737 145172
rect 119823 145132 119840 145172
rect 119880 145132 119889 145172
rect 119503 145109 119569 145132
rect 119655 145109 119737 145132
rect 119823 145109 119889 145132
rect 119503 145090 119889 145109
rect 134623 145195 135009 145214
rect 134623 145172 134689 145195
rect 134775 145172 134857 145195
rect 134943 145172 135009 145195
rect 134623 145132 134632 145172
rect 134672 145132 134689 145172
rect 134775 145132 134796 145172
rect 134836 145132 134857 145172
rect 134943 145132 134960 145172
rect 135000 145132 135009 145172
rect 134623 145109 134689 145132
rect 134775 145109 134857 145132
rect 134943 145109 135009 145132
rect 134623 145090 135009 145109
rect 149743 145195 150129 145214
rect 149743 145172 149809 145195
rect 149895 145172 149977 145195
rect 150063 145172 150129 145195
rect 149743 145132 149752 145172
rect 149792 145132 149809 145172
rect 149895 145132 149916 145172
rect 149956 145132 149977 145172
rect 150063 145132 150080 145172
rect 150120 145132 150129 145172
rect 149743 145109 149809 145132
rect 149895 145109 149977 145132
rect 150063 145109 150129 145132
rect 149743 145090 150129 145109
rect 75383 144439 75769 144458
rect 75383 144416 75449 144439
rect 75535 144416 75617 144439
rect 75703 144416 75769 144439
rect 75383 144376 75392 144416
rect 75432 144376 75449 144416
rect 75535 144376 75556 144416
rect 75596 144376 75617 144416
rect 75703 144376 75720 144416
rect 75760 144376 75769 144416
rect 75383 144353 75449 144376
rect 75535 144353 75617 144376
rect 75703 144353 75769 144376
rect 75383 144334 75769 144353
rect 90503 144439 90889 144458
rect 90503 144416 90569 144439
rect 90655 144416 90737 144439
rect 90823 144416 90889 144439
rect 90503 144376 90512 144416
rect 90552 144376 90569 144416
rect 90655 144376 90676 144416
rect 90716 144376 90737 144416
rect 90823 144376 90840 144416
rect 90880 144376 90889 144416
rect 90503 144353 90569 144376
rect 90655 144353 90737 144376
rect 90823 144353 90889 144376
rect 90503 144334 90889 144353
rect 105623 144439 106009 144458
rect 105623 144416 105689 144439
rect 105775 144416 105857 144439
rect 105943 144416 106009 144439
rect 105623 144376 105632 144416
rect 105672 144376 105689 144416
rect 105775 144376 105796 144416
rect 105836 144376 105857 144416
rect 105943 144376 105960 144416
rect 106000 144376 106009 144416
rect 105623 144353 105689 144376
rect 105775 144353 105857 144376
rect 105943 144353 106009 144376
rect 105623 144334 106009 144353
rect 120743 144439 121129 144458
rect 120743 144416 120809 144439
rect 120895 144416 120977 144439
rect 121063 144416 121129 144439
rect 120743 144376 120752 144416
rect 120792 144376 120809 144416
rect 120895 144376 120916 144416
rect 120956 144376 120977 144416
rect 121063 144376 121080 144416
rect 121120 144376 121129 144416
rect 120743 144353 120809 144376
rect 120895 144353 120977 144376
rect 121063 144353 121129 144376
rect 120743 144334 121129 144353
rect 135863 144439 136249 144458
rect 135863 144416 135929 144439
rect 136015 144416 136097 144439
rect 136183 144416 136249 144439
rect 135863 144376 135872 144416
rect 135912 144376 135929 144416
rect 136015 144376 136036 144416
rect 136076 144376 136097 144416
rect 136183 144376 136200 144416
rect 136240 144376 136249 144416
rect 135863 144353 135929 144376
rect 136015 144353 136097 144376
rect 136183 144353 136249 144376
rect 135863 144334 136249 144353
rect 150983 144439 151369 144458
rect 150983 144416 151049 144439
rect 151135 144416 151217 144439
rect 151303 144416 151369 144439
rect 150983 144376 150992 144416
rect 151032 144376 151049 144416
rect 151135 144376 151156 144416
rect 151196 144376 151217 144416
rect 151303 144376 151320 144416
rect 151360 144376 151369 144416
rect 150983 144353 151049 144376
rect 151135 144353 151217 144376
rect 151303 144353 151369 144376
rect 150983 144334 151369 144353
rect 74143 143683 74529 143702
rect 74143 143660 74209 143683
rect 74295 143660 74377 143683
rect 74463 143660 74529 143683
rect 74143 143620 74152 143660
rect 74192 143620 74209 143660
rect 74295 143620 74316 143660
rect 74356 143620 74377 143660
rect 74463 143620 74480 143660
rect 74520 143620 74529 143660
rect 74143 143597 74209 143620
rect 74295 143597 74377 143620
rect 74463 143597 74529 143620
rect 74143 143578 74529 143597
rect 89263 143683 89649 143702
rect 89263 143660 89329 143683
rect 89415 143660 89497 143683
rect 89583 143660 89649 143683
rect 89263 143620 89272 143660
rect 89312 143620 89329 143660
rect 89415 143620 89436 143660
rect 89476 143620 89497 143660
rect 89583 143620 89600 143660
rect 89640 143620 89649 143660
rect 89263 143597 89329 143620
rect 89415 143597 89497 143620
rect 89583 143597 89649 143620
rect 89263 143578 89649 143597
rect 104383 143683 104769 143702
rect 104383 143660 104449 143683
rect 104535 143660 104617 143683
rect 104703 143660 104769 143683
rect 104383 143620 104392 143660
rect 104432 143620 104449 143660
rect 104535 143620 104556 143660
rect 104596 143620 104617 143660
rect 104703 143620 104720 143660
rect 104760 143620 104769 143660
rect 104383 143597 104449 143620
rect 104535 143597 104617 143620
rect 104703 143597 104769 143620
rect 104383 143578 104769 143597
rect 119503 143683 119889 143702
rect 119503 143660 119569 143683
rect 119655 143660 119737 143683
rect 119823 143660 119889 143683
rect 119503 143620 119512 143660
rect 119552 143620 119569 143660
rect 119655 143620 119676 143660
rect 119716 143620 119737 143660
rect 119823 143620 119840 143660
rect 119880 143620 119889 143660
rect 119503 143597 119569 143620
rect 119655 143597 119737 143620
rect 119823 143597 119889 143620
rect 119503 143578 119889 143597
rect 134623 143683 135009 143702
rect 134623 143660 134689 143683
rect 134775 143660 134857 143683
rect 134943 143660 135009 143683
rect 134623 143620 134632 143660
rect 134672 143620 134689 143660
rect 134775 143620 134796 143660
rect 134836 143620 134857 143660
rect 134943 143620 134960 143660
rect 135000 143620 135009 143660
rect 134623 143597 134689 143620
rect 134775 143597 134857 143620
rect 134943 143597 135009 143620
rect 134623 143578 135009 143597
rect 149743 143683 150129 143702
rect 149743 143660 149809 143683
rect 149895 143660 149977 143683
rect 150063 143660 150129 143683
rect 149743 143620 149752 143660
rect 149792 143620 149809 143660
rect 149895 143620 149916 143660
rect 149956 143620 149977 143660
rect 150063 143620 150080 143660
rect 150120 143620 150129 143660
rect 149743 143597 149809 143620
rect 149895 143597 149977 143620
rect 150063 143597 150129 143620
rect 149743 143578 150129 143597
rect 75383 142927 75769 142946
rect 75383 142904 75449 142927
rect 75535 142904 75617 142927
rect 75703 142904 75769 142927
rect 75383 142864 75392 142904
rect 75432 142864 75449 142904
rect 75535 142864 75556 142904
rect 75596 142864 75617 142904
rect 75703 142864 75720 142904
rect 75760 142864 75769 142904
rect 75383 142841 75449 142864
rect 75535 142841 75617 142864
rect 75703 142841 75769 142864
rect 75383 142822 75769 142841
rect 90503 142927 90889 142946
rect 90503 142904 90569 142927
rect 90655 142904 90737 142927
rect 90823 142904 90889 142927
rect 90503 142864 90512 142904
rect 90552 142864 90569 142904
rect 90655 142864 90676 142904
rect 90716 142864 90737 142904
rect 90823 142864 90840 142904
rect 90880 142864 90889 142904
rect 90503 142841 90569 142864
rect 90655 142841 90737 142864
rect 90823 142841 90889 142864
rect 90503 142822 90889 142841
rect 105623 142927 106009 142946
rect 105623 142904 105689 142927
rect 105775 142904 105857 142927
rect 105943 142904 106009 142927
rect 105623 142864 105632 142904
rect 105672 142864 105689 142904
rect 105775 142864 105796 142904
rect 105836 142864 105857 142904
rect 105943 142864 105960 142904
rect 106000 142864 106009 142904
rect 105623 142841 105689 142864
rect 105775 142841 105857 142864
rect 105943 142841 106009 142864
rect 105623 142822 106009 142841
rect 120743 142927 121129 142946
rect 120743 142904 120809 142927
rect 120895 142904 120977 142927
rect 121063 142904 121129 142927
rect 120743 142864 120752 142904
rect 120792 142864 120809 142904
rect 120895 142864 120916 142904
rect 120956 142864 120977 142904
rect 121063 142864 121080 142904
rect 121120 142864 121129 142904
rect 120743 142841 120809 142864
rect 120895 142841 120977 142864
rect 121063 142841 121129 142864
rect 120743 142822 121129 142841
rect 135863 142927 136249 142946
rect 135863 142904 135929 142927
rect 136015 142904 136097 142927
rect 136183 142904 136249 142927
rect 135863 142864 135872 142904
rect 135912 142864 135929 142904
rect 136015 142864 136036 142904
rect 136076 142864 136097 142904
rect 136183 142864 136200 142904
rect 136240 142864 136249 142904
rect 135863 142841 135929 142864
rect 136015 142841 136097 142864
rect 136183 142841 136249 142864
rect 135863 142822 136249 142841
rect 150983 142927 151369 142946
rect 150983 142904 151049 142927
rect 151135 142904 151217 142927
rect 151303 142904 151369 142927
rect 150983 142864 150992 142904
rect 151032 142864 151049 142904
rect 151135 142864 151156 142904
rect 151196 142864 151217 142904
rect 151303 142864 151320 142904
rect 151360 142864 151369 142904
rect 150983 142841 151049 142864
rect 151135 142841 151217 142864
rect 151303 142841 151369 142864
rect 150983 142822 151369 142841
rect 74143 142171 74529 142190
rect 74143 142148 74209 142171
rect 74295 142148 74377 142171
rect 74463 142148 74529 142171
rect 74143 142108 74152 142148
rect 74192 142108 74209 142148
rect 74295 142108 74316 142148
rect 74356 142108 74377 142148
rect 74463 142108 74480 142148
rect 74520 142108 74529 142148
rect 74143 142085 74209 142108
rect 74295 142085 74377 142108
rect 74463 142085 74529 142108
rect 74143 142066 74529 142085
rect 89263 142171 89649 142190
rect 89263 142148 89329 142171
rect 89415 142148 89497 142171
rect 89583 142148 89649 142171
rect 89263 142108 89272 142148
rect 89312 142108 89329 142148
rect 89415 142108 89436 142148
rect 89476 142108 89497 142148
rect 89583 142108 89600 142148
rect 89640 142108 89649 142148
rect 89263 142085 89329 142108
rect 89415 142085 89497 142108
rect 89583 142085 89649 142108
rect 89263 142066 89649 142085
rect 104383 142171 104769 142190
rect 104383 142148 104449 142171
rect 104535 142148 104617 142171
rect 104703 142148 104769 142171
rect 104383 142108 104392 142148
rect 104432 142108 104449 142148
rect 104535 142108 104556 142148
rect 104596 142108 104617 142148
rect 104703 142108 104720 142148
rect 104760 142108 104769 142148
rect 104383 142085 104449 142108
rect 104535 142085 104617 142108
rect 104703 142085 104769 142108
rect 104383 142066 104769 142085
rect 119503 142171 119889 142190
rect 119503 142148 119569 142171
rect 119655 142148 119737 142171
rect 119823 142148 119889 142171
rect 119503 142108 119512 142148
rect 119552 142108 119569 142148
rect 119655 142108 119676 142148
rect 119716 142108 119737 142148
rect 119823 142108 119840 142148
rect 119880 142108 119889 142148
rect 119503 142085 119569 142108
rect 119655 142085 119737 142108
rect 119823 142085 119889 142108
rect 119503 142066 119889 142085
rect 134623 142171 135009 142190
rect 134623 142148 134689 142171
rect 134775 142148 134857 142171
rect 134943 142148 135009 142171
rect 134623 142108 134632 142148
rect 134672 142108 134689 142148
rect 134775 142108 134796 142148
rect 134836 142108 134857 142148
rect 134943 142108 134960 142148
rect 135000 142108 135009 142148
rect 134623 142085 134689 142108
rect 134775 142085 134857 142108
rect 134943 142085 135009 142108
rect 134623 142066 135009 142085
rect 149743 142171 150129 142190
rect 149743 142148 149809 142171
rect 149895 142148 149977 142171
rect 150063 142148 150129 142171
rect 149743 142108 149752 142148
rect 149792 142108 149809 142148
rect 149895 142108 149916 142148
rect 149956 142108 149977 142148
rect 150063 142108 150080 142148
rect 150120 142108 150129 142148
rect 149743 142085 149809 142108
rect 149895 142085 149977 142108
rect 150063 142085 150129 142108
rect 149743 142066 150129 142085
rect 75383 141415 75769 141434
rect 75383 141392 75449 141415
rect 75535 141392 75617 141415
rect 75703 141392 75769 141415
rect 75383 141352 75392 141392
rect 75432 141352 75449 141392
rect 75535 141352 75556 141392
rect 75596 141352 75617 141392
rect 75703 141352 75720 141392
rect 75760 141352 75769 141392
rect 75383 141329 75449 141352
rect 75535 141329 75617 141352
rect 75703 141329 75769 141352
rect 75383 141310 75769 141329
rect 90503 141415 90889 141434
rect 90503 141392 90569 141415
rect 90655 141392 90737 141415
rect 90823 141392 90889 141415
rect 90503 141352 90512 141392
rect 90552 141352 90569 141392
rect 90655 141352 90676 141392
rect 90716 141352 90737 141392
rect 90823 141352 90840 141392
rect 90880 141352 90889 141392
rect 90503 141329 90569 141352
rect 90655 141329 90737 141352
rect 90823 141329 90889 141352
rect 90503 141310 90889 141329
rect 105623 141415 106009 141434
rect 105623 141392 105689 141415
rect 105775 141392 105857 141415
rect 105943 141392 106009 141415
rect 105623 141352 105632 141392
rect 105672 141352 105689 141392
rect 105775 141352 105796 141392
rect 105836 141352 105857 141392
rect 105943 141352 105960 141392
rect 106000 141352 106009 141392
rect 105623 141329 105689 141352
rect 105775 141329 105857 141352
rect 105943 141329 106009 141352
rect 105623 141310 106009 141329
rect 120743 141415 121129 141434
rect 120743 141392 120809 141415
rect 120895 141392 120977 141415
rect 121063 141392 121129 141415
rect 120743 141352 120752 141392
rect 120792 141352 120809 141392
rect 120895 141352 120916 141392
rect 120956 141352 120977 141392
rect 121063 141352 121080 141392
rect 121120 141352 121129 141392
rect 120743 141329 120809 141352
rect 120895 141329 120977 141352
rect 121063 141329 121129 141352
rect 120743 141310 121129 141329
rect 135863 141415 136249 141434
rect 135863 141392 135929 141415
rect 136015 141392 136097 141415
rect 136183 141392 136249 141415
rect 135863 141352 135872 141392
rect 135912 141352 135929 141392
rect 136015 141352 136036 141392
rect 136076 141352 136097 141392
rect 136183 141352 136200 141392
rect 136240 141352 136249 141392
rect 135863 141329 135929 141352
rect 136015 141329 136097 141352
rect 136183 141329 136249 141352
rect 135863 141310 136249 141329
rect 150983 141415 151369 141434
rect 150983 141392 151049 141415
rect 151135 141392 151217 141415
rect 151303 141392 151369 141415
rect 150983 141352 150992 141392
rect 151032 141352 151049 141392
rect 151135 141352 151156 141392
rect 151196 141352 151217 141392
rect 151303 141352 151320 141392
rect 151360 141352 151369 141392
rect 150983 141329 151049 141352
rect 151135 141329 151217 141352
rect 151303 141329 151369 141352
rect 150983 141310 151369 141329
rect 74143 140659 74529 140678
rect 74143 140636 74209 140659
rect 74295 140636 74377 140659
rect 74463 140636 74529 140659
rect 74143 140596 74152 140636
rect 74192 140596 74209 140636
rect 74295 140596 74316 140636
rect 74356 140596 74377 140636
rect 74463 140596 74480 140636
rect 74520 140596 74529 140636
rect 74143 140573 74209 140596
rect 74295 140573 74377 140596
rect 74463 140573 74529 140596
rect 74143 140554 74529 140573
rect 89263 140659 89649 140678
rect 89263 140636 89329 140659
rect 89415 140636 89497 140659
rect 89583 140636 89649 140659
rect 89263 140596 89272 140636
rect 89312 140596 89329 140636
rect 89415 140596 89436 140636
rect 89476 140596 89497 140636
rect 89583 140596 89600 140636
rect 89640 140596 89649 140636
rect 89263 140573 89329 140596
rect 89415 140573 89497 140596
rect 89583 140573 89649 140596
rect 89263 140554 89649 140573
rect 104383 140659 104769 140678
rect 104383 140636 104449 140659
rect 104535 140636 104617 140659
rect 104703 140636 104769 140659
rect 104383 140596 104392 140636
rect 104432 140596 104449 140636
rect 104535 140596 104556 140636
rect 104596 140596 104617 140636
rect 104703 140596 104720 140636
rect 104760 140596 104769 140636
rect 104383 140573 104449 140596
rect 104535 140573 104617 140596
rect 104703 140573 104769 140596
rect 104383 140554 104769 140573
rect 119503 140659 119889 140678
rect 119503 140636 119569 140659
rect 119655 140636 119737 140659
rect 119823 140636 119889 140659
rect 119503 140596 119512 140636
rect 119552 140596 119569 140636
rect 119655 140596 119676 140636
rect 119716 140596 119737 140636
rect 119823 140596 119840 140636
rect 119880 140596 119889 140636
rect 119503 140573 119569 140596
rect 119655 140573 119737 140596
rect 119823 140573 119889 140596
rect 119503 140554 119889 140573
rect 134623 140659 135009 140678
rect 134623 140636 134689 140659
rect 134775 140636 134857 140659
rect 134943 140636 135009 140659
rect 134623 140596 134632 140636
rect 134672 140596 134689 140636
rect 134775 140596 134796 140636
rect 134836 140596 134857 140636
rect 134943 140596 134960 140636
rect 135000 140596 135009 140636
rect 134623 140573 134689 140596
rect 134775 140573 134857 140596
rect 134943 140573 135009 140596
rect 134623 140554 135009 140573
rect 149743 140659 150129 140678
rect 149743 140636 149809 140659
rect 149895 140636 149977 140659
rect 150063 140636 150129 140659
rect 149743 140596 149752 140636
rect 149792 140596 149809 140636
rect 149895 140596 149916 140636
rect 149956 140596 149977 140636
rect 150063 140596 150080 140636
rect 150120 140596 150129 140636
rect 149743 140573 149809 140596
rect 149895 140573 149977 140596
rect 150063 140573 150129 140596
rect 149743 140554 150129 140573
rect 75383 139903 75769 139922
rect 75383 139880 75449 139903
rect 75535 139880 75617 139903
rect 75703 139880 75769 139903
rect 75383 139840 75392 139880
rect 75432 139840 75449 139880
rect 75535 139840 75556 139880
rect 75596 139840 75617 139880
rect 75703 139840 75720 139880
rect 75760 139840 75769 139880
rect 75383 139817 75449 139840
rect 75535 139817 75617 139840
rect 75703 139817 75769 139840
rect 75383 139798 75769 139817
rect 90503 139903 90889 139922
rect 90503 139880 90569 139903
rect 90655 139880 90737 139903
rect 90823 139880 90889 139903
rect 90503 139840 90512 139880
rect 90552 139840 90569 139880
rect 90655 139840 90676 139880
rect 90716 139840 90737 139880
rect 90823 139840 90840 139880
rect 90880 139840 90889 139880
rect 90503 139817 90569 139840
rect 90655 139817 90737 139840
rect 90823 139817 90889 139840
rect 90503 139798 90889 139817
rect 105623 139903 106009 139922
rect 105623 139880 105689 139903
rect 105775 139880 105857 139903
rect 105943 139880 106009 139903
rect 105623 139840 105632 139880
rect 105672 139840 105689 139880
rect 105775 139840 105796 139880
rect 105836 139840 105857 139880
rect 105943 139840 105960 139880
rect 106000 139840 106009 139880
rect 105623 139817 105689 139840
rect 105775 139817 105857 139840
rect 105943 139817 106009 139840
rect 105623 139798 106009 139817
rect 120743 139903 121129 139922
rect 120743 139880 120809 139903
rect 120895 139880 120977 139903
rect 121063 139880 121129 139903
rect 120743 139840 120752 139880
rect 120792 139840 120809 139880
rect 120895 139840 120916 139880
rect 120956 139840 120977 139880
rect 121063 139840 121080 139880
rect 121120 139840 121129 139880
rect 120743 139817 120809 139840
rect 120895 139817 120977 139840
rect 121063 139817 121129 139840
rect 120743 139798 121129 139817
rect 135863 139903 136249 139922
rect 135863 139880 135929 139903
rect 136015 139880 136097 139903
rect 136183 139880 136249 139903
rect 135863 139840 135872 139880
rect 135912 139840 135929 139880
rect 136015 139840 136036 139880
rect 136076 139840 136097 139880
rect 136183 139840 136200 139880
rect 136240 139840 136249 139880
rect 135863 139817 135929 139840
rect 136015 139817 136097 139840
rect 136183 139817 136249 139840
rect 135863 139798 136249 139817
rect 150983 139903 151369 139922
rect 150983 139880 151049 139903
rect 151135 139880 151217 139903
rect 151303 139880 151369 139903
rect 150983 139840 150992 139880
rect 151032 139840 151049 139880
rect 151135 139840 151156 139880
rect 151196 139840 151217 139880
rect 151303 139840 151320 139880
rect 151360 139840 151369 139880
rect 150983 139817 151049 139840
rect 151135 139817 151217 139840
rect 151303 139817 151369 139840
rect 150983 139798 151369 139817
rect 74143 139147 74529 139166
rect 74143 139124 74209 139147
rect 74295 139124 74377 139147
rect 74463 139124 74529 139147
rect 74143 139084 74152 139124
rect 74192 139084 74209 139124
rect 74295 139084 74316 139124
rect 74356 139084 74377 139124
rect 74463 139084 74480 139124
rect 74520 139084 74529 139124
rect 74143 139061 74209 139084
rect 74295 139061 74377 139084
rect 74463 139061 74529 139084
rect 74143 139042 74529 139061
rect 89263 139147 89649 139166
rect 89263 139124 89329 139147
rect 89415 139124 89497 139147
rect 89583 139124 89649 139147
rect 89263 139084 89272 139124
rect 89312 139084 89329 139124
rect 89415 139084 89436 139124
rect 89476 139084 89497 139124
rect 89583 139084 89600 139124
rect 89640 139084 89649 139124
rect 89263 139061 89329 139084
rect 89415 139061 89497 139084
rect 89583 139061 89649 139084
rect 89263 139042 89649 139061
rect 104383 139147 104769 139166
rect 104383 139124 104449 139147
rect 104535 139124 104617 139147
rect 104703 139124 104769 139147
rect 104383 139084 104392 139124
rect 104432 139084 104449 139124
rect 104535 139084 104556 139124
rect 104596 139084 104617 139124
rect 104703 139084 104720 139124
rect 104760 139084 104769 139124
rect 104383 139061 104449 139084
rect 104535 139061 104617 139084
rect 104703 139061 104769 139084
rect 104383 139042 104769 139061
rect 119503 139147 119889 139166
rect 119503 139124 119569 139147
rect 119655 139124 119737 139147
rect 119823 139124 119889 139147
rect 119503 139084 119512 139124
rect 119552 139084 119569 139124
rect 119655 139084 119676 139124
rect 119716 139084 119737 139124
rect 119823 139084 119840 139124
rect 119880 139084 119889 139124
rect 119503 139061 119569 139084
rect 119655 139061 119737 139084
rect 119823 139061 119889 139084
rect 119503 139042 119889 139061
rect 134623 139147 135009 139166
rect 134623 139124 134689 139147
rect 134775 139124 134857 139147
rect 134943 139124 135009 139147
rect 134623 139084 134632 139124
rect 134672 139084 134689 139124
rect 134775 139084 134796 139124
rect 134836 139084 134857 139124
rect 134943 139084 134960 139124
rect 135000 139084 135009 139124
rect 134623 139061 134689 139084
rect 134775 139061 134857 139084
rect 134943 139061 135009 139084
rect 134623 139042 135009 139061
rect 149743 139147 150129 139166
rect 149743 139124 149809 139147
rect 149895 139124 149977 139147
rect 150063 139124 150129 139147
rect 149743 139084 149752 139124
rect 149792 139084 149809 139124
rect 149895 139084 149916 139124
rect 149956 139084 149977 139124
rect 150063 139084 150080 139124
rect 150120 139084 150129 139124
rect 149743 139061 149809 139084
rect 149895 139061 149977 139084
rect 150063 139061 150129 139084
rect 149743 139042 150129 139061
rect 75383 138391 75769 138410
rect 75383 138368 75449 138391
rect 75535 138368 75617 138391
rect 75703 138368 75769 138391
rect 75383 138328 75392 138368
rect 75432 138328 75449 138368
rect 75535 138328 75556 138368
rect 75596 138328 75617 138368
rect 75703 138328 75720 138368
rect 75760 138328 75769 138368
rect 75383 138305 75449 138328
rect 75535 138305 75617 138328
rect 75703 138305 75769 138328
rect 75383 138286 75769 138305
rect 90503 138391 90889 138410
rect 90503 138368 90569 138391
rect 90655 138368 90737 138391
rect 90823 138368 90889 138391
rect 90503 138328 90512 138368
rect 90552 138328 90569 138368
rect 90655 138328 90676 138368
rect 90716 138328 90737 138368
rect 90823 138328 90840 138368
rect 90880 138328 90889 138368
rect 90503 138305 90569 138328
rect 90655 138305 90737 138328
rect 90823 138305 90889 138328
rect 90503 138286 90889 138305
rect 105623 138391 106009 138410
rect 105623 138368 105689 138391
rect 105775 138368 105857 138391
rect 105943 138368 106009 138391
rect 105623 138328 105632 138368
rect 105672 138328 105689 138368
rect 105775 138328 105796 138368
rect 105836 138328 105857 138368
rect 105943 138328 105960 138368
rect 106000 138328 106009 138368
rect 105623 138305 105689 138328
rect 105775 138305 105857 138328
rect 105943 138305 106009 138328
rect 105623 138286 106009 138305
rect 120743 138391 121129 138410
rect 120743 138368 120809 138391
rect 120895 138368 120977 138391
rect 121063 138368 121129 138391
rect 120743 138328 120752 138368
rect 120792 138328 120809 138368
rect 120895 138328 120916 138368
rect 120956 138328 120977 138368
rect 121063 138328 121080 138368
rect 121120 138328 121129 138368
rect 120743 138305 120809 138328
rect 120895 138305 120977 138328
rect 121063 138305 121129 138328
rect 120743 138286 121129 138305
rect 135863 138391 136249 138410
rect 135863 138368 135929 138391
rect 136015 138368 136097 138391
rect 136183 138368 136249 138391
rect 135863 138328 135872 138368
rect 135912 138328 135929 138368
rect 136015 138328 136036 138368
rect 136076 138328 136097 138368
rect 136183 138328 136200 138368
rect 136240 138328 136249 138368
rect 135863 138305 135929 138328
rect 136015 138305 136097 138328
rect 136183 138305 136249 138328
rect 135863 138286 136249 138305
rect 150983 138391 151369 138410
rect 150983 138368 151049 138391
rect 151135 138368 151217 138391
rect 151303 138368 151369 138391
rect 150983 138328 150992 138368
rect 151032 138328 151049 138368
rect 151135 138328 151156 138368
rect 151196 138328 151217 138368
rect 151303 138328 151320 138368
rect 151360 138328 151369 138368
rect 150983 138305 151049 138328
rect 151135 138305 151217 138328
rect 151303 138305 151369 138328
rect 150983 138286 151369 138305
rect 74143 137635 74529 137654
rect 74143 137612 74209 137635
rect 74295 137612 74377 137635
rect 74463 137612 74529 137635
rect 74143 137572 74152 137612
rect 74192 137572 74209 137612
rect 74295 137572 74316 137612
rect 74356 137572 74377 137612
rect 74463 137572 74480 137612
rect 74520 137572 74529 137612
rect 74143 137549 74209 137572
rect 74295 137549 74377 137572
rect 74463 137549 74529 137572
rect 74143 137530 74529 137549
rect 89263 137635 89649 137654
rect 89263 137612 89329 137635
rect 89415 137612 89497 137635
rect 89583 137612 89649 137635
rect 89263 137572 89272 137612
rect 89312 137572 89329 137612
rect 89415 137572 89436 137612
rect 89476 137572 89497 137612
rect 89583 137572 89600 137612
rect 89640 137572 89649 137612
rect 89263 137549 89329 137572
rect 89415 137549 89497 137572
rect 89583 137549 89649 137572
rect 89263 137530 89649 137549
rect 104383 137635 104769 137654
rect 104383 137612 104449 137635
rect 104535 137612 104617 137635
rect 104703 137612 104769 137635
rect 104383 137572 104392 137612
rect 104432 137572 104449 137612
rect 104535 137572 104556 137612
rect 104596 137572 104617 137612
rect 104703 137572 104720 137612
rect 104760 137572 104769 137612
rect 104383 137549 104449 137572
rect 104535 137549 104617 137572
rect 104703 137549 104769 137572
rect 104383 137530 104769 137549
rect 119503 137635 119889 137654
rect 119503 137612 119569 137635
rect 119655 137612 119737 137635
rect 119823 137612 119889 137635
rect 119503 137572 119512 137612
rect 119552 137572 119569 137612
rect 119655 137572 119676 137612
rect 119716 137572 119737 137612
rect 119823 137572 119840 137612
rect 119880 137572 119889 137612
rect 119503 137549 119569 137572
rect 119655 137549 119737 137572
rect 119823 137549 119889 137572
rect 119503 137530 119889 137549
rect 134623 137635 135009 137654
rect 134623 137612 134689 137635
rect 134775 137612 134857 137635
rect 134943 137612 135009 137635
rect 134623 137572 134632 137612
rect 134672 137572 134689 137612
rect 134775 137572 134796 137612
rect 134836 137572 134857 137612
rect 134943 137572 134960 137612
rect 135000 137572 135009 137612
rect 134623 137549 134689 137572
rect 134775 137549 134857 137572
rect 134943 137549 135009 137572
rect 134623 137530 135009 137549
rect 149743 137635 150129 137654
rect 149743 137612 149809 137635
rect 149895 137612 149977 137635
rect 150063 137612 150129 137635
rect 149743 137572 149752 137612
rect 149792 137572 149809 137612
rect 149895 137572 149916 137612
rect 149956 137572 149977 137612
rect 150063 137572 150080 137612
rect 150120 137572 150129 137612
rect 149743 137549 149809 137572
rect 149895 137549 149977 137572
rect 150063 137549 150129 137572
rect 149743 137530 150129 137549
rect 75383 136879 75769 136898
rect 75383 136856 75449 136879
rect 75535 136856 75617 136879
rect 75703 136856 75769 136879
rect 75383 136816 75392 136856
rect 75432 136816 75449 136856
rect 75535 136816 75556 136856
rect 75596 136816 75617 136856
rect 75703 136816 75720 136856
rect 75760 136816 75769 136856
rect 75383 136793 75449 136816
rect 75535 136793 75617 136816
rect 75703 136793 75769 136816
rect 75383 136774 75769 136793
rect 90503 136879 90889 136898
rect 90503 136856 90569 136879
rect 90655 136856 90737 136879
rect 90823 136856 90889 136879
rect 90503 136816 90512 136856
rect 90552 136816 90569 136856
rect 90655 136816 90676 136856
rect 90716 136816 90737 136856
rect 90823 136816 90840 136856
rect 90880 136816 90889 136856
rect 90503 136793 90569 136816
rect 90655 136793 90737 136816
rect 90823 136793 90889 136816
rect 90503 136774 90889 136793
rect 105623 136879 106009 136898
rect 105623 136856 105689 136879
rect 105775 136856 105857 136879
rect 105943 136856 106009 136879
rect 105623 136816 105632 136856
rect 105672 136816 105689 136856
rect 105775 136816 105796 136856
rect 105836 136816 105857 136856
rect 105943 136816 105960 136856
rect 106000 136816 106009 136856
rect 105623 136793 105689 136816
rect 105775 136793 105857 136816
rect 105943 136793 106009 136816
rect 105623 136774 106009 136793
rect 120743 136879 121129 136898
rect 120743 136856 120809 136879
rect 120895 136856 120977 136879
rect 121063 136856 121129 136879
rect 120743 136816 120752 136856
rect 120792 136816 120809 136856
rect 120895 136816 120916 136856
rect 120956 136816 120977 136856
rect 121063 136816 121080 136856
rect 121120 136816 121129 136856
rect 120743 136793 120809 136816
rect 120895 136793 120977 136816
rect 121063 136793 121129 136816
rect 120743 136774 121129 136793
rect 135863 136879 136249 136898
rect 135863 136856 135929 136879
rect 136015 136856 136097 136879
rect 136183 136856 136249 136879
rect 135863 136816 135872 136856
rect 135912 136816 135929 136856
rect 136015 136816 136036 136856
rect 136076 136816 136097 136856
rect 136183 136816 136200 136856
rect 136240 136816 136249 136856
rect 135863 136793 135929 136816
rect 136015 136793 136097 136816
rect 136183 136793 136249 136816
rect 135863 136774 136249 136793
rect 150983 136879 151369 136898
rect 150983 136856 151049 136879
rect 151135 136856 151217 136879
rect 151303 136856 151369 136879
rect 150983 136816 150992 136856
rect 151032 136816 151049 136856
rect 151135 136816 151156 136856
rect 151196 136816 151217 136856
rect 151303 136816 151320 136856
rect 151360 136816 151369 136856
rect 150983 136793 151049 136816
rect 151135 136793 151217 136816
rect 151303 136793 151369 136816
rect 150983 136774 151369 136793
rect 74143 136123 74529 136142
rect 74143 136100 74209 136123
rect 74295 136100 74377 136123
rect 74463 136100 74529 136123
rect 74143 136060 74152 136100
rect 74192 136060 74209 136100
rect 74295 136060 74316 136100
rect 74356 136060 74377 136100
rect 74463 136060 74480 136100
rect 74520 136060 74529 136100
rect 74143 136037 74209 136060
rect 74295 136037 74377 136060
rect 74463 136037 74529 136060
rect 74143 136018 74529 136037
rect 89263 136123 89649 136142
rect 89263 136100 89329 136123
rect 89415 136100 89497 136123
rect 89583 136100 89649 136123
rect 89263 136060 89272 136100
rect 89312 136060 89329 136100
rect 89415 136060 89436 136100
rect 89476 136060 89497 136100
rect 89583 136060 89600 136100
rect 89640 136060 89649 136100
rect 89263 136037 89329 136060
rect 89415 136037 89497 136060
rect 89583 136037 89649 136060
rect 89263 136018 89649 136037
rect 104383 136123 104769 136142
rect 104383 136100 104449 136123
rect 104535 136100 104617 136123
rect 104703 136100 104769 136123
rect 104383 136060 104392 136100
rect 104432 136060 104449 136100
rect 104535 136060 104556 136100
rect 104596 136060 104617 136100
rect 104703 136060 104720 136100
rect 104760 136060 104769 136100
rect 104383 136037 104449 136060
rect 104535 136037 104617 136060
rect 104703 136037 104769 136060
rect 104383 136018 104769 136037
rect 119503 136123 119889 136142
rect 119503 136100 119569 136123
rect 119655 136100 119737 136123
rect 119823 136100 119889 136123
rect 119503 136060 119512 136100
rect 119552 136060 119569 136100
rect 119655 136060 119676 136100
rect 119716 136060 119737 136100
rect 119823 136060 119840 136100
rect 119880 136060 119889 136100
rect 119503 136037 119569 136060
rect 119655 136037 119737 136060
rect 119823 136037 119889 136060
rect 119503 136018 119889 136037
rect 134623 136123 135009 136142
rect 134623 136100 134689 136123
rect 134775 136100 134857 136123
rect 134943 136100 135009 136123
rect 134623 136060 134632 136100
rect 134672 136060 134689 136100
rect 134775 136060 134796 136100
rect 134836 136060 134857 136100
rect 134943 136060 134960 136100
rect 135000 136060 135009 136100
rect 134623 136037 134689 136060
rect 134775 136037 134857 136060
rect 134943 136037 135009 136060
rect 134623 136018 135009 136037
rect 149743 136123 150129 136142
rect 149743 136100 149809 136123
rect 149895 136100 149977 136123
rect 150063 136100 150129 136123
rect 149743 136060 149752 136100
rect 149792 136060 149809 136100
rect 149895 136060 149916 136100
rect 149956 136060 149977 136100
rect 150063 136060 150080 136100
rect 150120 136060 150129 136100
rect 149743 136037 149809 136060
rect 149895 136037 149977 136060
rect 150063 136037 150129 136060
rect 149743 136018 150129 136037
rect 75383 135367 75769 135386
rect 75383 135344 75449 135367
rect 75535 135344 75617 135367
rect 75703 135344 75769 135367
rect 75383 135304 75392 135344
rect 75432 135304 75449 135344
rect 75535 135304 75556 135344
rect 75596 135304 75617 135344
rect 75703 135304 75720 135344
rect 75760 135304 75769 135344
rect 75383 135281 75449 135304
rect 75535 135281 75617 135304
rect 75703 135281 75769 135304
rect 75383 135262 75769 135281
rect 90503 135367 90889 135386
rect 90503 135344 90569 135367
rect 90655 135344 90737 135367
rect 90823 135344 90889 135367
rect 90503 135304 90512 135344
rect 90552 135304 90569 135344
rect 90655 135304 90676 135344
rect 90716 135304 90737 135344
rect 90823 135304 90840 135344
rect 90880 135304 90889 135344
rect 90503 135281 90569 135304
rect 90655 135281 90737 135304
rect 90823 135281 90889 135304
rect 90503 135262 90889 135281
rect 105623 135367 106009 135386
rect 105623 135344 105689 135367
rect 105775 135344 105857 135367
rect 105943 135344 106009 135367
rect 105623 135304 105632 135344
rect 105672 135304 105689 135344
rect 105775 135304 105796 135344
rect 105836 135304 105857 135344
rect 105943 135304 105960 135344
rect 106000 135304 106009 135344
rect 105623 135281 105689 135304
rect 105775 135281 105857 135304
rect 105943 135281 106009 135304
rect 105623 135262 106009 135281
rect 120743 135367 121129 135386
rect 120743 135344 120809 135367
rect 120895 135344 120977 135367
rect 121063 135344 121129 135367
rect 120743 135304 120752 135344
rect 120792 135304 120809 135344
rect 120895 135304 120916 135344
rect 120956 135304 120977 135344
rect 121063 135304 121080 135344
rect 121120 135304 121129 135344
rect 120743 135281 120809 135304
rect 120895 135281 120977 135304
rect 121063 135281 121129 135304
rect 120743 135262 121129 135281
rect 135863 135367 136249 135386
rect 135863 135344 135929 135367
rect 136015 135344 136097 135367
rect 136183 135344 136249 135367
rect 135863 135304 135872 135344
rect 135912 135304 135929 135344
rect 136015 135304 136036 135344
rect 136076 135304 136097 135344
rect 136183 135304 136200 135344
rect 136240 135304 136249 135344
rect 135863 135281 135929 135304
rect 136015 135281 136097 135304
rect 136183 135281 136249 135304
rect 135863 135262 136249 135281
rect 150983 135367 151369 135386
rect 150983 135344 151049 135367
rect 151135 135344 151217 135367
rect 151303 135344 151369 135367
rect 150983 135304 150992 135344
rect 151032 135304 151049 135344
rect 151135 135304 151156 135344
rect 151196 135304 151217 135344
rect 151303 135304 151320 135344
rect 151360 135304 151369 135344
rect 150983 135281 151049 135304
rect 151135 135281 151217 135304
rect 151303 135281 151369 135304
rect 150983 135262 151369 135281
rect 74143 134611 74529 134630
rect 74143 134588 74209 134611
rect 74295 134588 74377 134611
rect 74463 134588 74529 134611
rect 74143 134548 74152 134588
rect 74192 134548 74209 134588
rect 74295 134548 74316 134588
rect 74356 134548 74377 134588
rect 74463 134548 74480 134588
rect 74520 134548 74529 134588
rect 74143 134525 74209 134548
rect 74295 134525 74377 134548
rect 74463 134525 74529 134548
rect 74143 134506 74529 134525
rect 89263 134611 89649 134630
rect 89263 134588 89329 134611
rect 89415 134588 89497 134611
rect 89583 134588 89649 134611
rect 89263 134548 89272 134588
rect 89312 134548 89329 134588
rect 89415 134548 89436 134588
rect 89476 134548 89497 134588
rect 89583 134548 89600 134588
rect 89640 134548 89649 134588
rect 89263 134525 89329 134548
rect 89415 134525 89497 134548
rect 89583 134525 89649 134548
rect 89263 134506 89649 134525
rect 104383 134611 104769 134630
rect 104383 134588 104449 134611
rect 104535 134588 104617 134611
rect 104703 134588 104769 134611
rect 104383 134548 104392 134588
rect 104432 134548 104449 134588
rect 104535 134548 104556 134588
rect 104596 134548 104617 134588
rect 104703 134548 104720 134588
rect 104760 134548 104769 134588
rect 104383 134525 104449 134548
rect 104535 134525 104617 134548
rect 104703 134525 104769 134548
rect 104383 134506 104769 134525
rect 119503 134611 119889 134630
rect 119503 134588 119569 134611
rect 119655 134588 119737 134611
rect 119823 134588 119889 134611
rect 119503 134548 119512 134588
rect 119552 134548 119569 134588
rect 119655 134548 119676 134588
rect 119716 134548 119737 134588
rect 119823 134548 119840 134588
rect 119880 134548 119889 134588
rect 119503 134525 119569 134548
rect 119655 134525 119737 134548
rect 119823 134525 119889 134548
rect 119503 134506 119889 134525
rect 134623 134611 135009 134630
rect 134623 134588 134689 134611
rect 134775 134588 134857 134611
rect 134943 134588 135009 134611
rect 134623 134548 134632 134588
rect 134672 134548 134689 134588
rect 134775 134548 134796 134588
rect 134836 134548 134857 134588
rect 134943 134548 134960 134588
rect 135000 134548 135009 134588
rect 134623 134525 134689 134548
rect 134775 134525 134857 134548
rect 134943 134525 135009 134548
rect 134623 134506 135009 134525
rect 149743 134611 150129 134630
rect 149743 134588 149809 134611
rect 149895 134588 149977 134611
rect 150063 134588 150129 134611
rect 149743 134548 149752 134588
rect 149792 134548 149809 134588
rect 149895 134548 149916 134588
rect 149956 134548 149977 134588
rect 150063 134548 150080 134588
rect 150120 134548 150129 134588
rect 149743 134525 149809 134548
rect 149895 134525 149977 134548
rect 150063 134525 150129 134548
rect 149743 134506 150129 134525
rect 75383 133855 75769 133874
rect 75383 133832 75449 133855
rect 75535 133832 75617 133855
rect 75703 133832 75769 133855
rect 75383 133792 75392 133832
rect 75432 133792 75449 133832
rect 75535 133792 75556 133832
rect 75596 133792 75617 133832
rect 75703 133792 75720 133832
rect 75760 133792 75769 133832
rect 75383 133769 75449 133792
rect 75535 133769 75617 133792
rect 75703 133769 75769 133792
rect 75383 133750 75769 133769
rect 90503 133855 90889 133874
rect 90503 133832 90569 133855
rect 90655 133832 90737 133855
rect 90823 133832 90889 133855
rect 90503 133792 90512 133832
rect 90552 133792 90569 133832
rect 90655 133792 90676 133832
rect 90716 133792 90737 133832
rect 90823 133792 90840 133832
rect 90880 133792 90889 133832
rect 90503 133769 90569 133792
rect 90655 133769 90737 133792
rect 90823 133769 90889 133792
rect 90503 133750 90889 133769
rect 105623 133855 106009 133874
rect 105623 133832 105689 133855
rect 105775 133832 105857 133855
rect 105943 133832 106009 133855
rect 105623 133792 105632 133832
rect 105672 133792 105689 133832
rect 105775 133792 105796 133832
rect 105836 133792 105857 133832
rect 105943 133792 105960 133832
rect 106000 133792 106009 133832
rect 105623 133769 105689 133792
rect 105775 133769 105857 133792
rect 105943 133769 106009 133792
rect 105623 133750 106009 133769
rect 120743 133855 121129 133874
rect 120743 133832 120809 133855
rect 120895 133832 120977 133855
rect 121063 133832 121129 133855
rect 120743 133792 120752 133832
rect 120792 133792 120809 133832
rect 120895 133792 120916 133832
rect 120956 133792 120977 133832
rect 121063 133792 121080 133832
rect 121120 133792 121129 133832
rect 120743 133769 120809 133792
rect 120895 133769 120977 133792
rect 121063 133769 121129 133792
rect 120743 133750 121129 133769
rect 135863 133855 136249 133874
rect 135863 133832 135929 133855
rect 136015 133832 136097 133855
rect 136183 133832 136249 133855
rect 135863 133792 135872 133832
rect 135912 133792 135929 133832
rect 136015 133792 136036 133832
rect 136076 133792 136097 133832
rect 136183 133792 136200 133832
rect 136240 133792 136249 133832
rect 135863 133769 135929 133792
rect 136015 133769 136097 133792
rect 136183 133769 136249 133792
rect 135863 133750 136249 133769
rect 150983 133855 151369 133874
rect 150983 133832 151049 133855
rect 151135 133832 151217 133855
rect 151303 133832 151369 133855
rect 150983 133792 150992 133832
rect 151032 133792 151049 133832
rect 151135 133792 151156 133832
rect 151196 133792 151217 133832
rect 151303 133792 151320 133832
rect 151360 133792 151369 133832
rect 150983 133769 151049 133792
rect 151135 133769 151217 133792
rect 151303 133769 151369 133792
rect 150983 133750 151369 133769
rect 74143 133099 74529 133118
rect 74143 133076 74209 133099
rect 74295 133076 74377 133099
rect 74463 133076 74529 133099
rect 74143 133036 74152 133076
rect 74192 133036 74209 133076
rect 74295 133036 74316 133076
rect 74356 133036 74377 133076
rect 74463 133036 74480 133076
rect 74520 133036 74529 133076
rect 74143 133013 74209 133036
rect 74295 133013 74377 133036
rect 74463 133013 74529 133036
rect 74143 132994 74529 133013
rect 89263 133099 89649 133118
rect 89263 133076 89329 133099
rect 89415 133076 89497 133099
rect 89583 133076 89649 133099
rect 89263 133036 89272 133076
rect 89312 133036 89329 133076
rect 89415 133036 89436 133076
rect 89476 133036 89497 133076
rect 89583 133036 89600 133076
rect 89640 133036 89649 133076
rect 89263 133013 89329 133036
rect 89415 133013 89497 133036
rect 89583 133013 89649 133036
rect 89263 132994 89649 133013
rect 104383 133099 104769 133118
rect 104383 133076 104449 133099
rect 104535 133076 104617 133099
rect 104703 133076 104769 133099
rect 104383 133036 104392 133076
rect 104432 133036 104449 133076
rect 104535 133036 104556 133076
rect 104596 133036 104617 133076
rect 104703 133036 104720 133076
rect 104760 133036 104769 133076
rect 104383 133013 104449 133036
rect 104535 133013 104617 133036
rect 104703 133013 104769 133036
rect 104383 132994 104769 133013
rect 119503 133099 119889 133118
rect 119503 133076 119569 133099
rect 119655 133076 119737 133099
rect 119823 133076 119889 133099
rect 119503 133036 119512 133076
rect 119552 133036 119569 133076
rect 119655 133036 119676 133076
rect 119716 133036 119737 133076
rect 119823 133036 119840 133076
rect 119880 133036 119889 133076
rect 119503 133013 119569 133036
rect 119655 133013 119737 133036
rect 119823 133013 119889 133036
rect 119503 132994 119889 133013
rect 134623 133099 135009 133118
rect 134623 133076 134689 133099
rect 134775 133076 134857 133099
rect 134943 133076 135009 133099
rect 134623 133036 134632 133076
rect 134672 133036 134689 133076
rect 134775 133036 134796 133076
rect 134836 133036 134857 133076
rect 134943 133036 134960 133076
rect 135000 133036 135009 133076
rect 134623 133013 134689 133036
rect 134775 133013 134857 133036
rect 134943 133013 135009 133036
rect 134623 132994 135009 133013
rect 149743 133099 150129 133118
rect 149743 133076 149809 133099
rect 149895 133076 149977 133099
rect 150063 133076 150129 133099
rect 149743 133036 149752 133076
rect 149792 133036 149809 133076
rect 149895 133036 149916 133076
rect 149956 133036 149977 133076
rect 150063 133036 150080 133076
rect 150120 133036 150129 133076
rect 149743 133013 149809 133036
rect 149895 133013 149977 133036
rect 150063 133013 150129 133036
rect 149743 132994 150129 133013
rect 75383 132343 75769 132362
rect 75383 132320 75449 132343
rect 75535 132320 75617 132343
rect 75703 132320 75769 132343
rect 75383 132280 75392 132320
rect 75432 132280 75449 132320
rect 75535 132280 75556 132320
rect 75596 132280 75617 132320
rect 75703 132280 75720 132320
rect 75760 132280 75769 132320
rect 75383 132257 75449 132280
rect 75535 132257 75617 132280
rect 75703 132257 75769 132280
rect 75383 132238 75769 132257
rect 90503 132343 90889 132362
rect 90503 132320 90569 132343
rect 90655 132320 90737 132343
rect 90823 132320 90889 132343
rect 90503 132280 90512 132320
rect 90552 132280 90569 132320
rect 90655 132280 90676 132320
rect 90716 132280 90737 132320
rect 90823 132280 90840 132320
rect 90880 132280 90889 132320
rect 90503 132257 90569 132280
rect 90655 132257 90737 132280
rect 90823 132257 90889 132280
rect 90503 132238 90889 132257
rect 105623 132343 106009 132362
rect 105623 132320 105689 132343
rect 105775 132320 105857 132343
rect 105943 132320 106009 132343
rect 105623 132280 105632 132320
rect 105672 132280 105689 132320
rect 105775 132280 105796 132320
rect 105836 132280 105857 132320
rect 105943 132280 105960 132320
rect 106000 132280 106009 132320
rect 105623 132257 105689 132280
rect 105775 132257 105857 132280
rect 105943 132257 106009 132280
rect 105623 132238 106009 132257
rect 120743 132343 121129 132362
rect 120743 132320 120809 132343
rect 120895 132320 120977 132343
rect 121063 132320 121129 132343
rect 120743 132280 120752 132320
rect 120792 132280 120809 132320
rect 120895 132280 120916 132320
rect 120956 132280 120977 132320
rect 121063 132280 121080 132320
rect 121120 132280 121129 132320
rect 120743 132257 120809 132280
rect 120895 132257 120977 132280
rect 121063 132257 121129 132280
rect 120743 132238 121129 132257
rect 135863 132343 136249 132362
rect 135863 132320 135929 132343
rect 136015 132320 136097 132343
rect 136183 132320 136249 132343
rect 135863 132280 135872 132320
rect 135912 132280 135929 132320
rect 136015 132280 136036 132320
rect 136076 132280 136097 132320
rect 136183 132280 136200 132320
rect 136240 132280 136249 132320
rect 135863 132257 135929 132280
rect 136015 132257 136097 132280
rect 136183 132257 136249 132280
rect 135863 132238 136249 132257
rect 150983 132343 151369 132362
rect 150983 132320 151049 132343
rect 151135 132320 151217 132343
rect 151303 132320 151369 132343
rect 150983 132280 150992 132320
rect 151032 132280 151049 132320
rect 151135 132280 151156 132320
rect 151196 132280 151217 132320
rect 151303 132280 151320 132320
rect 151360 132280 151369 132320
rect 150983 132257 151049 132280
rect 151135 132257 151217 132280
rect 151303 132257 151369 132280
rect 150983 132238 151369 132257
rect 74143 131587 74529 131606
rect 74143 131564 74209 131587
rect 74295 131564 74377 131587
rect 74463 131564 74529 131587
rect 74143 131524 74152 131564
rect 74192 131524 74209 131564
rect 74295 131524 74316 131564
rect 74356 131524 74377 131564
rect 74463 131524 74480 131564
rect 74520 131524 74529 131564
rect 74143 131501 74209 131524
rect 74295 131501 74377 131524
rect 74463 131501 74529 131524
rect 74143 131482 74529 131501
rect 89263 131587 89649 131606
rect 89263 131564 89329 131587
rect 89415 131564 89497 131587
rect 89583 131564 89649 131587
rect 89263 131524 89272 131564
rect 89312 131524 89329 131564
rect 89415 131524 89436 131564
rect 89476 131524 89497 131564
rect 89583 131524 89600 131564
rect 89640 131524 89649 131564
rect 89263 131501 89329 131524
rect 89415 131501 89497 131524
rect 89583 131501 89649 131524
rect 89263 131482 89649 131501
rect 104383 131587 104769 131606
rect 104383 131564 104449 131587
rect 104535 131564 104617 131587
rect 104703 131564 104769 131587
rect 104383 131524 104392 131564
rect 104432 131524 104449 131564
rect 104535 131524 104556 131564
rect 104596 131524 104617 131564
rect 104703 131524 104720 131564
rect 104760 131524 104769 131564
rect 104383 131501 104449 131524
rect 104535 131501 104617 131524
rect 104703 131501 104769 131524
rect 104383 131482 104769 131501
rect 119503 131587 119889 131606
rect 119503 131564 119569 131587
rect 119655 131564 119737 131587
rect 119823 131564 119889 131587
rect 119503 131524 119512 131564
rect 119552 131524 119569 131564
rect 119655 131524 119676 131564
rect 119716 131524 119737 131564
rect 119823 131524 119840 131564
rect 119880 131524 119889 131564
rect 119503 131501 119569 131524
rect 119655 131501 119737 131524
rect 119823 131501 119889 131524
rect 119503 131482 119889 131501
rect 134623 131587 135009 131606
rect 134623 131564 134689 131587
rect 134775 131564 134857 131587
rect 134943 131564 135009 131587
rect 134623 131524 134632 131564
rect 134672 131524 134689 131564
rect 134775 131524 134796 131564
rect 134836 131524 134857 131564
rect 134943 131524 134960 131564
rect 135000 131524 135009 131564
rect 134623 131501 134689 131524
rect 134775 131501 134857 131524
rect 134943 131501 135009 131524
rect 134623 131482 135009 131501
rect 149743 131587 150129 131606
rect 149743 131564 149809 131587
rect 149895 131564 149977 131587
rect 150063 131564 150129 131587
rect 149743 131524 149752 131564
rect 149792 131524 149809 131564
rect 149895 131524 149916 131564
rect 149956 131524 149977 131564
rect 150063 131524 150080 131564
rect 150120 131524 150129 131564
rect 149743 131501 149809 131524
rect 149895 131501 149977 131524
rect 150063 131501 150129 131524
rect 149743 131482 150129 131501
rect 75383 130831 75769 130850
rect 75383 130808 75449 130831
rect 75535 130808 75617 130831
rect 75703 130808 75769 130831
rect 75383 130768 75392 130808
rect 75432 130768 75449 130808
rect 75535 130768 75556 130808
rect 75596 130768 75617 130808
rect 75703 130768 75720 130808
rect 75760 130768 75769 130808
rect 75383 130745 75449 130768
rect 75535 130745 75617 130768
rect 75703 130745 75769 130768
rect 75383 130726 75769 130745
rect 90503 130831 90889 130850
rect 90503 130808 90569 130831
rect 90655 130808 90737 130831
rect 90823 130808 90889 130831
rect 90503 130768 90512 130808
rect 90552 130768 90569 130808
rect 90655 130768 90676 130808
rect 90716 130768 90737 130808
rect 90823 130768 90840 130808
rect 90880 130768 90889 130808
rect 90503 130745 90569 130768
rect 90655 130745 90737 130768
rect 90823 130745 90889 130768
rect 90503 130726 90889 130745
rect 105623 130831 106009 130850
rect 105623 130808 105689 130831
rect 105775 130808 105857 130831
rect 105943 130808 106009 130831
rect 105623 130768 105632 130808
rect 105672 130768 105689 130808
rect 105775 130768 105796 130808
rect 105836 130768 105857 130808
rect 105943 130768 105960 130808
rect 106000 130768 106009 130808
rect 105623 130745 105689 130768
rect 105775 130745 105857 130768
rect 105943 130745 106009 130768
rect 105623 130726 106009 130745
rect 120743 130831 121129 130850
rect 120743 130808 120809 130831
rect 120895 130808 120977 130831
rect 121063 130808 121129 130831
rect 120743 130768 120752 130808
rect 120792 130768 120809 130808
rect 120895 130768 120916 130808
rect 120956 130768 120977 130808
rect 121063 130768 121080 130808
rect 121120 130768 121129 130808
rect 120743 130745 120809 130768
rect 120895 130745 120977 130768
rect 121063 130745 121129 130768
rect 120743 130726 121129 130745
rect 135863 130831 136249 130850
rect 135863 130808 135929 130831
rect 136015 130808 136097 130831
rect 136183 130808 136249 130831
rect 135863 130768 135872 130808
rect 135912 130768 135929 130808
rect 136015 130768 136036 130808
rect 136076 130768 136097 130808
rect 136183 130768 136200 130808
rect 136240 130768 136249 130808
rect 135863 130745 135929 130768
rect 136015 130745 136097 130768
rect 136183 130745 136249 130768
rect 135863 130726 136249 130745
rect 150983 130831 151369 130850
rect 150983 130808 151049 130831
rect 151135 130808 151217 130831
rect 151303 130808 151369 130831
rect 150983 130768 150992 130808
rect 151032 130768 151049 130808
rect 151135 130768 151156 130808
rect 151196 130768 151217 130808
rect 151303 130768 151320 130808
rect 151360 130768 151369 130808
rect 150983 130745 151049 130768
rect 151135 130745 151217 130768
rect 151303 130745 151369 130768
rect 150983 130726 151369 130745
rect 74143 130075 74529 130094
rect 74143 130052 74209 130075
rect 74295 130052 74377 130075
rect 74463 130052 74529 130075
rect 74143 130012 74152 130052
rect 74192 130012 74209 130052
rect 74295 130012 74316 130052
rect 74356 130012 74377 130052
rect 74463 130012 74480 130052
rect 74520 130012 74529 130052
rect 74143 129989 74209 130012
rect 74295 129989 74377 130012
rect 74463 129989 74529 130012
rect 74143 129970 74529 129989
rect 89263 130075 89649 130094
rect 89263 130052 89329 130075
rect 89415 130052 89497 130075
rect 89583 130052 89649 130075
rect 89263 130012 89272 130052
rect 89312 130012 89329 130052
rect 89415 130012 89436 130052
rect 89476 130012 89497 130052
rect 89583 130012 89600 130052
rect 89640 130012 89649 130052
rect 89263 129989 89329 130012
rect 89415 129989 89497 130012
rect 89583 129989 89649 130012
rect 89263 129970 89649 129989
rect 104383 130075 104769 130094
rect 104383 130052 104449 130075
rect 104535 130052 104617 130075
rect 104703 130052 104769 130075
rect 104383 130012 104392 130052
rect 104432 130012 104449 130052
rect 104535 130012 104556 130052
rect 104596 130012 104617 130052
rect 104703 130012 104720 130052
rect 104760 130012 104769 130052
rect 104383 129989 104449 130012
rect 104535 129989 104617 130012
rect 104703 129989 104769 130012
rect 104383 129970 104769 129989
rect 119503 130075 119889 130094
rect 119503 130052 119569 130075
rect 119655 130052 119737 130075
rect 119823 130052 119889 130075
rect 119503 130012 119512 130052
rect 119552 130012 119569 130052
rect 119655 130012 119676 130052
rect 119716 130012 119737 130052
rect 119823 130012 119840 130052
rect 119880 130012 119889 130052
rect 119503 129989 119569 130012
rect 119655 129989 119737 130012
rect 119823 129989 119889 130012
rect 119503 129970 119889 129989
rect 134623 130075 135009 130094
rect 134623 130052 134689 130075
rect 134775 130052 134857 130075
rect 134943 130052 135009 130075
rect 134623 130012 134632 130052
rect 134672 130012 134689 130052
rect 134775 130012 134796 130052
rect 134836 130012 134857 130052
rect 134943 130012 134960 130052
rect 135000 130012 135009 130052
rect 134623 129989 134689 130012
rect 134775 129989 134857 130012
rect 134943 129989 135009 130012
rect 134623 129970 135009 129989
rect 149743 130075 150129 130094
rect 149743 130052 149809 130075
rect 149895 130052 149977 130075
rect 150063 130052 150129 130075
rect 149743 130012 149752 130052
rect 149792 130012 149809 130052
rect 149895 130012 149916 130052
rect 149956 130012 149977 130052
rect 150063 130012 150080 130052
rect 150120 130012 150129 130052
rect 149743 129989 149809 130012
rect 149895 129989 149977 130012
rect 150063 129989 150129 130012
rect 149743 129970 150129 129989
rect 75383 129319 75769 129338
rect 75383 129296 75449 129319
rect 75535 129296 75617 129319
rect 75703 129296 75769 129319
rect 75383 129256 75392 129296
rect 75432 129256 75449 129296
rect 75535 129256 75556 129296
rect 75596 129256 75617 129296
rect 75703 129256 75720 129296
rect 75760 129256 75769 129296
rect 75383 129233 75449 129256
rect 75535 129233 75617 129256
rect 75703 129233 75769 129256
rect 75383 129214 75769 129233
rect 90503 129319 90889 129338
rect 90503 129296 90569 129319
rect 90655 129296 90737 129319
rect 90823 129296 90889 129319
rect 90503 129256 90512 129296
rect 90552 129256 90569 129296
rect 90655 129256 90676 129296
rect 90716 129256 90737 129296
rect 90823 129256 90840 129296
rect 90880 129256 90889 129296
rect 90503 129233 90569 129256
rect 90655 129233 90737 129256
rect 90823 129233 90889 129256
rect 90503 129214 90889 129233
rect 105623 129319 106009 129338
rect 105623 129296 105689 129319
rect 105775 129296 105857 129319
rect 105943 129296 106009 129319
rect 105623 129256 105632 129296
rect 105672 129256 105689 129296
rect 105775 129256 105796 129296
rect 105836 129256 105857 129296
rect 105943 129256 105960 129296
rect 106000 129256 106009 129296
rect 105623 129233 105689 129256
rect 105775 129233 105857 129256
rect 105943 129233 106009 129256
rect 105623 129214 106009 129233
rect 120743 129319 121129 129338
rect 120743 129296 120809 129319
rect 120895 129296 120977 129319
rect 121063 129296 121129 129319
rect 120743 129256 120752 129296
rect 120792 129256 120809 129296
rect 120895 129256 120916 129296
rect 120956 129256 120977 129296
rect 121063 129256 121080 129296
rect 121120 129256 121129 129296
rect 120743 129233 120809 129256
rect 120895 129233 120977 129256
rect 121063 129233 121129 129256
rect 120743 129214 121129 129233
rect 135863 129319 136249 129338
rect 135863 129296 135929 129319
rect 136015 129296 136097 129319
rect 136183 129296 136249 129319
rect 135863 129256 135872 129296
rect 135912 129256 135929 129296
rect 136015 129256 136036 129296
rect 136076 129256 136097 129296
rect 136183 129256 136200 129296
rect 136240 129256 136249 129296
rect 135863 129233 135929 129256
rect 136015 129233 136097 129256
rect 136183 129233 136249 129256
rect 135863 129214 136249 129233
rect 150983 129319 151369 129338
rect 150983 129296 151049 129319
rect 151135 129296 151217 129319
rect 151303 129296 151369 129319
rect 150983 129256 150992 129296
rect 151032 129256 151049 129296
rect 151135 129256 151156 129296
rect 151196 129256 151217 129296
rect 151303 129256 151320 129296
rect 151360 129256 151369 129296
rect 150983 129233 151049 129256
rect 151135 129233 151217 129256
rect 151303 129233 151369 129256
rect 150983 129214 151369 129233
rect 74143 128563 74529 128582
rect 74143 128540 74209 128563
rect 74295 128540 74377 128563
rect 74463 128540 74529 128563
rect 74143 128500 74152 128540
rect 74192 128500 74209 128540
rect 74295 128500 74316 128540
rect 74356 128500 74377 128540
rect 74463 128500 74480 128540
rect 74520 128500 74529 128540
rect 74143 128477 74209 128500
rect 74295 128477 74377 128500
rect 74463 128477 74529 128500
rect 74143 128458 74529 128477
rect 89263 128563 89649 128582
rect 89263 128540 89329 128563
rect 89415 128540 89497 128563
rect 89583 128540 89649 128563
rect 89263 128500 89272 128540
rect 89312 128500 89329 128540
rect 89415 128500 89436 128540
rect 89476 128500 89497 128540
rect 89583 128500 89600 128540
rect 89640 128500 89649 128540
rect 89263 128477 89329 128500
rect 89415 128477 89497 128500
rect 89583 128477 89649 128500
rect 89263 128458 89649 128477
rect 104383 128563 104769 128582
rect 104383 128540 104449 128563
rect 104535 128540 104617 128563
rect 104703 128540 104769 128563
rect 104383 128500 104392 128540
rect 104432 128500 104449 128540
rect 104535 128500 104556 128540
rect 104596 128500 104617 128540
rect 104703 128500 104720 128540
rect 104760 128500 104769 128540
rect 104383 128477 104449 128500
rect 104535 128477 104617 128500
rect 104703 128477 104769 128500
rect 104383 128458 104769 128477
rect 119503 128563 119889 128582
rect 119503 128540 119569 128563
rect 119655 128540 119737 128563
rect 119823 128540 119889 128563
rect 119503 128500 119512 128540
rect 119552 128500 119569 128540
rect 119655 128500 119676 128540
rect 119716 128500 119737 128540
rect 119823 128500 119840 128540
rect 119880 128500 119889 128540
rect 119503 128477 119569 128500
rect 119655 128477 119737 128500
rect 119823 128477 119889 128500
rect 119503 128458 119889 128477
rect 134623 128563 135009 128582
rect 134623 128540 134689 128563
rect 134775 128540 134857 128563
rect 134943 128540 135009 128563
rect 134623 128500 134632 128540
rect 134672 128500 134689 128540
rect 134775 128500 134796 128540
rect 134836 128500 134857 128540
rect 134943 128500 134960 128540
rect 135000 128500 135009 128540
rect 134623 128477 134689 128500
rect 134775 128477 134857 128500
rect 134943 128477 135009 128500
rect 134623 128458 135009 128477
rect 149743 128563 150129 128582
rect 149743 128540 149809 128563
rect 149895 128540 149977 128563
rect 150063 128540 150129 128563
rect 149743 128500 149752 128540
rect 149792 128500 149809 128540
rect 149895 128500 149916 128540
rect 149956 128500 149977 128540
rect 150063 128500 150080 128540
rect 150120 128500 150129 128540
rect 149743 128477 149809 128500
rect 149895 128477 149977 128500
rect 150063 128477 150129 128500
rect 149743 128458 150129 128477
rect 75383 127807 75769 127826
rect 75383 127784 75449 127807
rect 75535 127784 75617 127807
rect 75703 127784 75769 127807
rect 75383 127744 75392 127784
rect 75432 127744 75449 127784
rect 75535 127744 75556 127784
rect 75596 127744 75617 127784
rect 75703 127744 75720 127784
rect 75760 127744 75769 127784
rect 75383 127721 75449 127744
rect 75535 127721 75617 127744
rect 75703 127721 75769 127744
rect 75383 127702 75769 127721
rect 90503 127807 90889 127826
rect 90503 127784 90569 127807
rect 90655 127784 90737 127807
rect 90823 127784 90889 127807
rect 90503 127744 90512 127784
rect 90552 127744 90569 127784
rect 90655 127744 90676 127784
rect 90716 127744 90737 127784
rect 90823 127744 90840 127784
rect 90880 127744 90889 127784
rect 90503 127721 90569 127744
rect 90655 127721 90737 127744
rect 90823 127721 90889 127744
rect 90503 127702 90889 127721
rect 105623 127807 106009 127826
rect 105623 127784 105689 127807
rect 105775 127784 105857 127807
rect 105943 127784 106009 127807
rect 105623 127744 105632 127784
rect 105672 127744 105689 127784
rect 105775 127744 105796 127784
rect 105836 127744 105857 127784
rect 105943 127744 105960 127784
rect 106000 127744 106009 127784
rect 105623 127721 105689 127744
rect 105775 127721 105857 127744
rect 105943 127721 106009 127744
rect 105623 127702 106009 127721
rect 120743 127807 121129 127826
rect 120743 127784 120809 127807
rect 120895 127784 120977 127807
rect 121063 127784 121129 127807
rect 120743 127744 120752 127784
rect 120792 127744 120809 127784
rect 120895 127744 120916 127784
rect 120956 127744 120977 127784
rect 121063 127744 121080 127784
rect 121120 127744 121129 127784
rect 120743 127721 120809 127744
rect 120895 127721 120977 127744
rect 121063 127721 121129 127744
rect 120743 127702 121129 127721
rect 135863 127807 136249 127826
rect 135863 127784 135929 127807
rect 136015 127784 136097 127807
rect 136183 127784 136249 127807
rect 135863 127744 135872 127784
rect 135912 127744 135929 127784
rect 136015 127744 136036 127784
rect 136076 127744 136097 127784
rect 136183 127744 136200 127784
rect 136240 127744 136249 127784
rect 135863 127721 135929 127744
rect 136015 127721 136097 127744
rect 136183 127721 136249 127744
rect 135863 127702 136249 127721
rect 150983 127807 151369 127826
rect 150983 127784 151049 127807
rect 151135 127784 151217 127807
rect 151303 127784 151369 127807
rect 150983 127744 150992 127784
rect 151032 127744 151049 127784
rect 151135 127744 151156 127784
rect 151196 127744 151217 127784
rect 151303 127744 151320 127784
rect 151360 127744 151369 127784
rect 150983 127721 151049 127744
rect 151135 127721 151217 127744
rect 151303 127721 151369 127744
rect 150983 127702 151369 127721
rect 74143 127051 74529 127070
rect 74143 127028 74209 127051
rect 74295 127028 74377 127051
rect 74463 127028 74529 127051
rect 74143 126988 74152 127028
rect 74192 126988 74209 127028
rect 74295 126988 74316 127028
rect 74356 126988 74377 127028
rect 74463 126988 74480 127028
rect 74520 126988 74529 127028
rect 74143 126965 74209 126988
rect 74295 126965 74377 126988
rect 74463 126965 74529 126988
rect 74143 126946 74529 126965
rect 89263 127051 89649 127070
rect 89263 127028 89329 127051
rect 89415 127028 89497 127051
rect 89583 127028 89649 127051
rect 89263 126988 89272 127028
rect 89312 126988 89329 127028
rect 89415 126988 89436 127028
rect 89476 126988 89497 127028
rect 89583 126988 89600 127028
rect 89640 126988 89649 127028
rect 89263 126965 89329 126988
rect 89415 126965 89497 126988
rect 89583 126965 89649 126988
rect 89263 126946 89649 126965
rect 104383 127051 104769 127070
rect 104383 127028 104449 127051
rect 104535 127028 104617 127051
rect 104703 127028 104769 127051
rect 104383 126988 104392 127028
rect 104432 126988 104449 127028
rect 104535 126988 104556 127028
rect 104596 126988 104617 127028
rect 104703 126988 104720 127028
rect 104760 126988 104769 127028
rect 104383 126965 104449 126988
rect 104535 126965 104617 126988
rect 104703 126965 104769 126988
rect 104383 126946 104769 126965
rect 119503 127051 119889 127070
rect 119503 127028 119569 127051
rect 119655 127028 119737 127051
rect 119823 127028 119889 127051
rect 119503 126988 119512 127028
rect 119552 126988 119569 127028
rect 119655 126988 119676 127028
rect 119716 126988 119737 127028
rect 119823 126988 119840 127028
rect 119880 126988 119889 127028
rect 119503 126965 119569 126988
rect 119655 126965 119737 126988
rect 119823 126965 119889 126988
rect 119503 126946 119889 126965
rect 134623 127051 135009 127070
rect 134623 127028 134689 127051
rect 134775 127028 134857 127051
rect 134943 127028 135009 127051
rect 134623 126988 134632 127028
rect 134672 126988 134689 127028
rect 134775 126988 134796 127028
rect 134836 126988 134857 127028
rect 134943 126988 134960 127028
rect 135000 126988 135009 127028
rect 134623 126965 134689 126988
rect 134775 126965 134857 126988
rect 134943 126965 135009 126988
rect 134623 126946 135009 126965
rect 149743 127051 150129 127070
rect 149743 127028 149809 127051
rect 149895 127028 149977 127051
rect 150063 127028 150129 127051
rect 149743 126988 149752 127028
rect 149792 126988 149809 127028
rect 149895 126988 149916 127028
rect 149956 126988 149977 127028
rect 150063 126988 150080 127028
rect 150120 126988 150129 127028
rect 149743 126965 149809 126988
rect 149895 126965 149977 126988
rect 150063 126965 150129 126988
rect 149743 126946 150129 126965
rect 75383 126295 75769 126314
rect 75383 126272 75449 126295
rect 75535 126272 75617 126295
rect 75703 126272 75769 126295
rect 75383 126232 75392 126272
rect 75432 126232 75449 126272
rect 75535 126232 75556 126272
rect 75596 126232 75617 126272
rect 75703 126232 75720 126272
rect 75760 126232 75769 126272
rect 75383 126209 75449 126232
rect 75535 126209 75617 126232
rect 75703 126209 75769 126232
rect 75383 126190 75769 126209
rect 90503 126295 90889 126314
rect 90503 126272 90569 126295
rect 90655 126272 90737 126295
rect 90823 126272 90889 126295
rect 90503 126232 90512 126272
rect 90552 126232 90569 126272
rect 90655 126232 90676 126272
rect 90716 126232 90737 126272
rect 90823 126232 90840 126272
rect 90880 126232 90889 126272
rect 90503 126209 90569 126232
rect 90655 126209 90737 126232
rect 90823 126209 90889 126232
rect 90503 126190 90889 126209
rect 105623 126295 106009 126314
rect 105623 126272 105689 126295
rect 105775 126272 105857 126295
rect 105943 126272 106009 126295
rect 105623 126232 105632 126272
rect 105672 126232 105689 126272
rect 105775 126232 105796 126272
rect 105836 126232 105857 126272
rect 105943 126232 105960 126272
rect 106000 126232 106009 126272
rect 105623 126209 105689 126232
rect 105775 126209 105857 126232
rect 105943 126209 106009 126232
rect 105623 126190 106009 126209
rect 120743 126295 121129 126314
rect 120743 126272 120809 126295
rect 120895 126272 120977 126295
rect 121063 126272 121129 126295
rect 120743 126232 120752 126272
rect 120792 126232 120809 126272
rect 120895 126232 120916 126272
rect 120956 126232 120977 126272
rect 121063 126232 121080 126272
rect 121120 126232 121129 126272
rect 120743 126209 120809 126232
rect 120895 126209 120977 126232
rect 121063 126209 121129 126232
rect 120743 126190 121129 126209
rect 135863 126295 136249 126314
rect 135863 126272 135929 126295
rect 136015 126272 136097 126295
rect 136183 126272 136249 126295
rect 135863 126232 135872 126272
rect 135912 126232 135929 126272
rect 136015 126232 136036 126272
rect 136076 126232 136097 126272
rect 136183 126232 136200 126272
rect 136240 126232 136249 126272
rect 135863 126209 135929 126232
rect 136015 126209 136097 126232
rect 136183 126209 136249 126232
rect 135863 126190 136249 126209
rect 150983 126295 151369 126314
rect 150983 126272 151049 126295
rect 151135 126272 151217 126295
rect 151303 126272 151369 126295
rect 150983 126232 150992 126272
rect 151032 126232 151049 126272
rect 151135 126232 151156 126272
rect 151196 126232 151217 126272
rect 151303 126232 151320 126272
rect 151360 126232 151369 126272
rect 150983 126209 151049 126232
rect 151135 126209 151217 126232
rect 151303 126209 151369 126232
rect 150983 126190 151369 126209
rect 74143 125539 74529 125558
rect 74143 125516 74209 125539
rect 74295 125516 74377 125539
rect 74463 125516 74529 125539
rect 74143 125476 74152 125516
rect 74192 125476 74209 125516
rect 74295 125476 74316 125516
rect 74356 125476 74377 125516
rect 74463 125476 74480 125516
rect 74520 125476 74529 125516
rect 74143 125453 74209 125476
rect 74295 125453 74377 125476
rect 74463 125453 74529 125476
rect 74143 125434 74529 125453
rect 89263 125539 89649 125558
rect 89263 125516 89329 125539
rect 89415 125516 89497 125539
rect 89583 125516 89649 125539
rect 89263 125476 89272 125516
rect 89312 125476 89329 125516
rect 89415 125476 89436 125516
rect 89476 125476 89497 125516
rect 89583 125476 89600 125516
rect 89640 125476 89649 125516
rect 89263 125453 89329 125476
rect 89415 125453 89497 125476
rect 89583 125453 89649 125476
rect 89263 125434 89649 125453
rect 104383 125539 104769 125558
rect 104383 125516 104449 125539
rect 104535 125516 104617 125539
rect 104703 125516 104769 125539
rect 104383 125476 104392 125516
rect 104432 125476 104449 125516
rect 104535 125476 104556 125516
rect 104596 125476 104617 125516
rect 104703 125476 104720 125516
rect 104760 125476 104769 125516
rect 104383 125453 104449 125476
rect 104535 125453 104617 125476
rect 104703 125453 104769 125476
rect 104383 125434 104769 125453
rect 119503 125539 119889 125558
rect 119503 125516 119569 125539
rect 119655 125516 119737 125539
rect 119823 125516 119889 125539
rect 119503 125476 119512 125516
rect 119552 125476 119569 125516
rect 119655 125476 119676 125516
rect 119716 125476 119737 125516
rect 119823 125476 119840 125516
rect 119880 125476 119889 125516
rect 119503 125453 119569 125476
rect 119655 125453 119737 125476
rect 119823 125453 119889 125476
rect 119503 125434 119889 125453
rect 134623 125539 135009 125558
rect 134623 125516 134689 125539
rect 134775 125516 134857 125539
rect 134943 125516 135009 125539
rect 134623 125476 134632 125516
rect 134672 125476 134689 125516
rect 134775 125476 134796 125516
rect 134836 125476 134857 125516
rect 134943 125476 134960 125516
rect 135000 125476 135009 125516
rect 134623 125453 134689 125476
rect 134775 125453 134857 125476
rect 134943 125453 135009 125476
rect 134623 125434 135009 125453
rect 149743 125539 150129 125558
rect 149743 125516 149809 125539
rect 149895 125516 149977 125539
rect 150063 125516 150129 125539
rect 149743 125476 149752 125516
rect 149792 125476 149809 125516
rect 149895 125476 149916 125516
rect 149956 125476 149977 125516
rect 150063 125476 150080 125516
rect 150120 125476 150129 125516
rect 149743 125453 149809 125476
rect 149895 125453 149977 125476
rect 150063 125453 150129 125476
rect 149743 125434 150129 125453
rect 75383 124783 75769 124802
rect 75383 124760 75449 124783
rect 75535 124760 75617 124783
rect 75703 124760 75769 124783
rect 75383 124720 75392 124760
rect 75432 124720 75449 124760
rect 75535 124720 75556 124760
rect 75596 124720 75617 124760
rect 75703 124720 75720 124760
rect 75760 124720 75769 124760
rect 75383 124697 75449 124720
rect 75535 124697 75617 124720
rect 75703 124697 75769 124720
rect 75383 124678 75769 124697
rect 90503 124783 90889 124802
rect 90503 124760 90569 124783
rect 90655 124760 90737 124783
rect 90823 124760 90889 124783
rect 90503 124720 90512 124760
rect 90552 124720 90569 124760
rect 90655 124720 90676 124760
rect 90716 124720 90737 124760
rect 90823 124720 90840 124760
rect 90880 124720 90889 124760
rect 90503 124697 90569 124720
rect 90655 124697 90737 124720
rect 90823 124697 90889 124720
rect 90503 124678 90889 124697
rect 105623 124783 106009 124802
rect 105623 124760 105689 124783
rect 105775 124760 105857 124783
rect 105943 124760 106009 124783
rect 105623 124720 105632 124760
rect 105672 124720 105689 124760
rect 105775 124720 105796 124760
rect 105836 124720 105857 124760
rect 105943 124720 105960 124760
rect 106000 124720 106009 124760
rect 105623 124697 105689 124720
rect 105775 124697 105857 124720
rect 105943 124697 106009 124720
rect 105623 124678 106009 124697
rect 120743 124783 121129 124802
rect 120743 124760 120809 124783
rect 120895 124760 120977 124783
rect 121063 124760 121129 124783
rect 120743 124720 120752 124760
rect 120792 124720 120809 124760
rect 120895 124720 120916 124760
rect 120956 124720 120977 124760
rect 121063 124720 121080 124760
rect 121120 124720 121129 124760
rect 120743 124697 120809 124720
rect 120895 124697 120977 124720
rect 121063 124697 121129 124720
rect 120743 124678 121129 124697
rect 135863 124783 136249 124802
rect 135863 124760 135929 124783
rect 136015 124760 136097 124783
rect 136183 124760 136249 124783
rect 135863 124720 135872 124760
rect 135912 124720 135929 124760
rect 136015 124720 136036 124760
rect 136076 124720 136097 124760
rect 136183 124720 136200 124760
rect 136240 124720 136249 124760
rect 135863 124697 135929 124720
rect 136015 124697 136097 124720
rect 136183 124697 136249 124720
rect 135863 124678 136249 124697
rect 150983 124783 151369 124802
rect 150983 124760 151049 124783
rect 151135 124760 151217 124783
rect 151303 124760 151369 124783
rect 150983 124720 150992 124760
rect 151032 124720 151049 124760
rect 151135 124720 151156 124760
rect 151196 124720 151217 124760
rect 151303 124720 151320 124760
rect 151360 124720 151369 124760
rect 150983 124697 151049 124720
rect 151135 124697 151217 124720
rect 151303 124697 151369 124720
rect 150983 124678 151369 124697
rect 74143 124027 74529 124046
rect 74143 124004 74209 124027
rect 74295 124004 74377 124027
rect 74463 124004 74529 124027
rect 74143 123964 74152 124004
rect 74192 123964 74209 124004
rect 74295 123964 74316 124004
rect 74356 123964 74377 124004
rect 74463 123964 74480 124004
rect 74520 123964 74529 124004
rect 74143 123941 74209 123964
rect 74295 123941 74377 123964
rect 74463 123941 74529 123964
rect 74143 123922 74529 123941
rect 89263 124027 89649 124046
rect 89263 124004 89329 124027
rect 89415 124004 89497 124027
rect 89583 124004 89649 124027
rect 89263 123964 89272 124004
rect 89312 123964 89329 124004
rect 89415 123964 89436 124004
rect 89476 123964 89497 124004
rect 89583 123964 89600 124004
rect 89640 123964 89649 124004
rect 89263 123941 89329 123964
rect 89415 123941 89497 123964
rect 89583 123941 89649 123964
rect 89263 123922 89649 123941
rect 104383 124027 104769 124046
rect 104383 124004 104449 124027
rect 104535 124004 104617 124027
rect 104703 124004 104769 124027
rect 104383 123964 104392 124004
rect 104432 123964 104449 124004
rect 104535 123964 104556 124004
rect 104596 123964 104617 124004
rect 104703 123964 104720 124004
rect 104760 123964 104769 124004
rect 104383 123941 104449 123964
rect 104535 123941 104617 123964
rect 104703 123941 104769 123964
rect 104383 123922 104769 123941
rect 119503 124027 119889 124046
rect 119503 124004 119569 124027
rect 119655 124004 119737 124027
rect 119823 124004 119889 124027
rect 119503 123964 119512 124004
rect 119552 123964 119569 124004
rect 119655 123964 119676 124004
rect 119716 123964 119737 124004
rect 119823 123964 119840 124004
rect 119880 123964 119889 124004
rect 119503 123941 119569 123964
rect 119655 123941 119737 123964
rect 119823 123941 119889 123964
rect 119503 123922 119889 123941
rect 134623 124027 135009 124046
rect 134623 124004 134689 124027
rect 134775 124004 134857 124027
rect 134943 124004 135009 124027
rect 134623 123964 134632 124004
rect 134672 123964 134689 124004
rect 134775 123964 134796 124004
rect 134836 123964 134857 124004
rect 134943 123964 134960 124004
rect 135000 123964 135009 124004
rect 134623 123941 134689 123964
rect 134775 123941 134857 123964
rect 134943 123941 135009 123964
rect 134623 123922 135009 123941
rect 149743 124027 150129 124046
rect 149743 124004 149809 124027
rect 149895 124004 149977 124027
rect 150063 124004 150129 124027
rect 149743 123964 149752 124004
rect 149792 123964 149809 124004
rect 149895 123964 149916 124004
rect 149956 123964 149977 124004
rect 150063 123964 150080 124004
rect 150120 123964 150129 124004
rect 149743 123941 149809 123964
rect 149895 123941 149977 123964
rect 150063 123941 150129 123964
rect 149743 123922 150129 123941
rect 75383 123271 75769 123290
rect 75383 123248 75449 123271
rect 75535 123248 75617 123271
rect 75703 123248 75769 123271
rect 75383 123208 75392 123248
rect 75432 123208 75449 123248
rect 75535 123208 75556 123248
rect 75596 123208 75617 123248
rect 75703 123208 75720 123248
rect 75760 123208 75769 123248
rect 75383 123185 75449 123208
rect 75535 123185 75617 123208
rect 75703 123185 75769 123208
rect 75383 123166 75769 123185
rect 90503 123271 90889 123290
rect 90503 123248 90569 123271
rect 90655 123248 90737 123271
rect 90823 123248 90889 123271
rect 90503 123208 90512 123248
rect 90552 123208 90569 123248
rect 90655 123208 90676 123248
rect 90716 123208 90737 123248
rect 90823 123208 90840 123248
rect 90880 123208 90889 123248
rect 90503 123185 90569 123208
rect 90655 123185 90737 123208
rect 90823 123185 90889 123208
rect 90503 123166 90889 123185
rect 105623 123271 106009 123290
rect 105623 123248 105689 123271
rect 105775 123248 105857 123271
rect 105943 123248 106009 123271
rect 105623 123208 105632 123248
rect 105672 123208 105689 123248
rect 105775 123208 105796 123248
rect 105836 123208 105857 123248
rect 105943 123208 105960 123248
rect 106000 123208 106009 123248
rect 105623 123185 105689 123208
rect 105775 123185 105857 123208
rect 105943 123185 106009 123208
rect 105623 123166 106009 123185
rect 120743 123271 121129 123290
rect 120743 123248 120809 123271
rect 120895 123248 120977 123271
rect 121063 123248 121129 123271
rect 120743 123208 120752 123248
rect 120792 123208 120809 123248
rect 120895 123208 120916 123248
rect 120956 123208 120977 123248
rect 121063 123208 121080 123248
rect 121120 123208 121129 123248
rect 120743 123185 120809 123208
rect 120895 123185 120977 123208
rect 121063 123185 121129 123208
rect 120743 123166 121129 123185
rect 135863 123271 136249 123290
rect 135863 123248 135929 123271
rect 136015 123248 136097 123271
rect 136183 123248 136249 123271
rect 135863 123208 135872 123248
rect 135912 123208 135929 123248
rect 136015 123208 136036 123248
rect 136076 123208 136097 123248
rect 136183 123208 136200 123248
rect 136240 123208 136249 123248
rect 135863 123185 135929 123208
rect 136015 123185 136097 123208
rect 136183 123185 136249 123208
rect 135863 123166 136249 123185
rect 150983 123271 151369 123290
rect 150983 123248 151049 123271
rect 151135 123248 151217 123271
rect 151303 123248 151369 123271
rect 150983 123208 150992 123248
rect 151032 123208 151049 123248
rect 151135 123208 151156 123248
rect 151196 123208 151217 123248
rect 151303 123208 151320 123248
rect 151360 123208 151369 123248
rect 150983 123185 151049 123208
rect 151135 123185 151217 123208
rect 151303 123185 151369 123208
rect 150983 123166 151369 123185
rect 74143 122515 74529 122534
rect 74143 122492 74209 122515
rect 74295 122492 74377 122515
rect 74463 122492 74529 122515
rect 74143 122452 74152 122492
rect 74192 122452 74209 122492
rect 74295 122452 74316 122492
rect 74356 122452 74377 122492
rect 74463 122452 74480 122492
rect 74520 122452 74529 122492
rect 74143 122429 74209 122452
rect 74295 122429 74377 122452
rect 74463 122429 74529 122452
rect 74143 122410 74529 122429
rect 89263 122515 89649 122534
rect 89263 122492 89329 122515
rect 89415 122492 89497 122515
rect 89583 122492 89649 122515
rect 89263 122452 89272 122492
rect 89312 122452 89329 122492
rect 89415 122452 89436 122492
rect 89476 122452 89497 122492
rect 89583 122452 89600 122492
rect 89640 122452 89649 122492
rect 89263 122429 89329 122452
rect 89415 122429 89497 122452
rect 89583 122429 89649 122452
rect 89263 122410 89649 122429
rect 104383 122515 104769 122534
rect 104383 122492 104449 122515
rect 104535 122492 104617 122515
rect 104703 122492 104769 122515
rect 104383 122452 104392 122492
rect 104432 122452 104449 122492
rect 104535 122452 104556 122492
rect 104596 122452 104617 122492
rect 104703 122452 104720 122492
rect 104760 122452 104769 122492
rect 104383 122429 104449 122452
rect 104535 122429 104617 122452
rect 104703 122429 104769 122452
rect 104383 122410 104769 122429
rect 119503 122515 119889 122534
rect 119503 122492 119569 122515
rect 119655 122492 119737 122515
rect 119823 122492 119889 122515
rect 119503 122452 119512 122492
rect 119552 122452 119569 122492
rect 119655 122452 119676 122492
rect 119716 122452 119737 122492
rect 119823 122452 119840 122492
rect 119880 122452 119889 122492
rect 119503 122429 119569 122452
rect 119655 122429 119737 122452
rect 119823 122429 119889 122452
rect 119503 122410 119889 122429
rect 134623 122515 135009 122534
rect 134623 122492 134689 122515
rect 134775 122492 134857 122515
rect 134943 122492 135009 122515
rect 134623 122452 134632 122492
rect 134672 122452 134689 122492
rect 134775 122452 134796 122492
rect 134836 122452 134857 122492
rect 134943 122452 134960 122492
rect 135000 122452 135009 122492
rect 134623 122429 134689 122452
rect 134775 122429 134857 122452
rect 134943 122429 135009 122452
rect 134623 122410 135009 122429
rect 149743 122515 150129 122534
rect 149743 122492 149809 122515
rect 149895 122492 149977 122515
rect 150063 122492 150129 122515
rect 149743 122452 149752 122492
rect 149792 122452 149809 122492
rect 149895 122452 149916 122492
rect 149956 122452 149977 122492
rect 150063 122452 150080 122492
rect 150120 122452 150129 122492
rect 149743 122429 149809 122452
rect 149895 122429 149977 122452
rect 150063 122429 150129 122452
rect 149743 122410 150129 122429
rect 75383 121759 75769 121778
rect 75383 121736 75449 121759
rect 75535 121736 75617 121759
rect 75703 121736 75769 121759
rect 75383 121696 75392 121736
rect 75432 121696 75449 121736
rect 75535 121696 75556 121736
rect 75596 121696 75617 121736
rect 75703 121696 75720 121736
rect 75760 121696 75769 121736
rect 75383 121673 75449 121696
rect 75535 121673 75617 121696
rect 75703 121673 75769 121696
rect 75383 121654 75769 121673
rect 90503 121759 90889 121778
rect 90503 121736 90569 121759
rect 90655 121736 90737 121759
rect 90823 121736 90889 121759
rect 90503 121696 90512 121736
rect 90552 121696 90569 121736
rect 90655 121696 90676 121736
rect 90716 121696 90737 121736
rect 90823 121696 90840 121736
rect 90880 121696 90889 121736
rect 90503 121673 90569 121696
rect 90655 121673 90737 121696
rect 90823 121673 90889 121696
rect 90503 121654 90889 121673
rect 105623 121759 106009 121778
rect 105623 121736 105689 121759
rect 105775 121736 105857 121759
rect 105943 121736 106009 121759
rect 105623 121696 105632 121736
rect 105672 121696 105689 121736
rect 105775 121696 105796 121736
rect 105836 121696 105857 121736
rect 105943 121696 105960 121736
rect 106000 121696 106009 121736
rect 105623 121673 105689 121696
rect 105775 121673 105857 121696
rect 105943 121673 106009 121696
rect 105623 121654 106009 121673
rect 120743 121759 121129 121778
rect 120743 121736 120809 121759
rect 120895 121736 120977 121759
rect 121063 121736 121129 121759
rect 120743 121696 120752 121736
rect 120792 121696 120809 121736
rect 120895 121696 120916 121736
rect 120956 121696 120977 121736
rect 121063 121696 121080 121736
rect 121120 121696 121129 121736
rect 120743 121673 120809 121696
rect 120895 121673 120977 121696
rect 121063 121673 121129 121696
rect 120743 121654 121129 121673
rect 135863 121759 136249 121778
rect 135863 121736 135929 121759
rect 136015 121736 136097 121759
rect 136183 121736 136249 121759
rect 135863 121696 135872 121736
rect 135912 121696 135929 121736
rect 136015 121696 136036 121736
rect 136076 121696 136097 121736
rect 136183 121696 136200 121736
rect 136240 121696 136249 121736
rect 135863 121673 135929 121696
rect 136015 121673 136097 121696
rect 136183 121673 136249 121696
rect 135863 121654 136249 121673
rect 150983 121759 151369 121778
rect 150983 121736 151049 121759
rect 151135 121736 151217 121759
rect 151303 121736 151369 121759
rect 150983 121696 150992 121736
rect 151032 121696 151049 121736
rect 151135 121696 151156 121736
rect 151196 121696 151217 121736
rect 151303 121696 151320 121736
rect 151360 121696 151369 121736
rect 150983 121673 151049 121696
rect 151135 121673 151217 121696
rect 151303 121673 151369 121696
rect 150983 121654 151369 121673
rect 74143 121003 74529 121022
rect 74143 120980 74209 121003
rect 74295 120980 74377 121003
rect 74463 120980 74529 121003
rect 74143 120940 74152 120980
rect 74192 120940 74209 120980
rect 74295 120940 74316 120980
rect 74356 120940 74377 120980
rect 74463 120940 74480 120980
rect 74520 120940 74529 120980
rect 74143 120917 74209 120940
rect 74295 120917 74377 120940
rect 74463 120917 74529 120940
rect 74143 120898 74529 120917
rect 89263 121003 89649 121022
rect 89263 120980 89329 121003
rect 89415 120980 89497 121003
rect 89583 120980 89649 121003
rect 89263 120940 89272 120980
rect 89312 120940 89329 120980
rect 89415 120940 89436 120980
rect 89476 120940 89497 120980
rect 89583 120940 89600 120980
rect 89640 120940 89649 120980
rect 89263 120917 89329 120940
rect 89415 120917 89497 120940
rect 89583 120917 89649 120940
rect 89263 120898 89649 120917
rect 104383 121003 104769 121022
rect 104383 120980 104449 121003
rect 104535 120980 104617 121003
rect 104703 120980 104769 121003
rect 104383 120940 104392 120980
rect 104432 120940 104449 120980
rect 104535 120940 104556 120980
rect 104596 120940 104617 120980
rect 104703 120940 104720 120980
rect 104760 120940 104769 120980
rect 104383 120917 104449 120940
rect 104535 120917 104617 120940
rect 104703 120917 104769 120940
rect 104383 120898 104769 120917
rect 119503 121003 119889 121022
rect 119503 120980 119569 121003
rect 119655 120980 119737 121003
rect 119823 120980 119889 121003
rect 119503 120940 119512 120980
rect 119552 120940 119569 120980
rect 119655 120940 119676 120980
rect 119716 120940 119737 120980
rect 119823 120940 119840 120980
rect 119880 120940 119889 120980
rect 119503 120917 119569 120940
rect 119655 120917 119737 120940
rect 119823 120917 119889 120940
rect 119503 120898 119889 120917
rect 134623 121003 135009 121022
rect 134623 120980 134689 121003
rect 134775 120980 134857 121003
rect 134943 120980 135009 121003
rect 134623 120940 134632 120980
rect 134672 120940 134689 120980
rect 134775 120940 134796 120980
rect 134836 120940 134857 120980
rect 134943 120940 134960 120980
rect 135000 120940 135009 120980
rect 134623 120917 134689 120940
rect 134775 120917 134857 120940
rect 134943 120917 135009 120940
rect 134623 120898 135009 120917
rect 149743 121003 150129 121022
rect 149743 120980 149809 121003
rect 149895 120980 149977 121003
rect 150063 120980 150129 121003
rect 149743 120940 149752 120980
rect 149792 120940 149809 120980
rect 149895 120940 149916 120980
rect 149956 120940 149977 120980
rect 150063 120940 150080 120980
rect 150120 120940 150129 120980
rect 149743 120917 149809 120940
rect 149895 120917 149977 120940
rect 150063 120917 150129 120940
rect 149743 120898 150129 120917
rect 75383 120247 75769 120266
rect 75383 120224 75449 120247
rect 75535 120224 75617 120247
rect 75703 120224 75769 120247
rect 75383 120184 75392 120224
rect 75432 120184 75449 120224
rect 75535 120184 75556 120224
rect 75596 120184 75617 120224
rect 75703 120184 75720 120224
rect 75760 120184 75769 120224
rect 75383 120161 75449 120184
rect 75535 120161 75617 120184
rect 75703 120161 75769 120184
rect 75383 120142 75769 120161
rect 90503 120247 90889 120266
rect 90503 120224 90569 120247
rect 90655 120224 90737 120247
rect 90823 120224 90889 120247
rect 90503 120184 90512 120224
rect 90552 120184 90569 120224
rect 90655 120184 90676 120224
rect 90716 120184 90737 120224
rect 90823 120184 90840 120224
rect 90880 120184 90889 120224
rect 90503 120161 90569 120184
rect 90655 120161 90737 120184
rect 90823 120161 90889 120184
rect 90503 120142 90889 120161
rect 105623 120247 106009 120266
rect 105623 120224 105689 120247
rect 105775 120224 105857 120247
rect 105943 120224 106009 120247
rect 105623 120184 105632 120224
rect 105672 120184 105689 120224
rect 105775 120184 105796 120224
rect 105836 120184 105857 120224
rect 105943 120184 105960 120224
rect 106000 120184 106009 120224
rect 105623 120161 105689 120184
rect 105775 120161 105857 120184
rect 105943 120161 106009 120184
rect 105623 120142 106009 120161
rect 120743 120247 121129 120266
rect 120743 120224 120809 120247
rect 120895 120224 120977 120247
rect 121063 120224 121129 120247
rect 120743 120184 120752 120224
rect 120792 120184 120809 120224
rect 120895 120184 120916 120224
rect 120956 120184 120977 120224
rect 121063 120184 121080 120224
rect 121120 120184 121129 120224
rect 120743 120161 120809 120184
rect 120895 120161 120977 120184
rect 121063 120161 121129 120184
rect 120743 120142 121129 120161
rect 135863 120247 136249 120266
rect 135863 120224 135929 120247
rect 136015 120224 136097 120247
rect 136183 120224 136249 120247
rect 135863 120184 135872 120224
rect 135912 120184 135929 120224
rect 136015 120184 136036 120224
rect 136076 120184 136097 120224
rect 136183 120184 136200 120224
rect 136240 120184 136249 120224
rect 135863 120161 135929 120184
rect 136015 120161 136097 120184
rect 136183 120161 136249 120184
rect 135863 120142 136249 120161
rect 150983 120247 151369 120266
rect 150983 120224 151049 120247
rect 151135 120224 151217 120247
rect 151303 120224 151369 120247
rect 150983 120184 150992 120224
rect 151032 120184 151049 120224
rect 151135 120184 151156 120224
rect 151196 120184 151217 120224
rect 151303 120184 151320 120224
rect 151360 120184 151369 120224
rect 150983 120161 151049 120184
rect 151135 120161 151217 120184
rect 151303 120161 151369 120184
rect 150983 120142 151369 120161
rect 74143 119491 74529 119510
rect 74143 119468 74209 119491
rect 74295 119468 74377 119491
rect 74463 119468 74529 119491
rect 74143 119428 74152 119468
rect 74192 119428 74209 119468
rect 74295 119428 74316 119468
rect 74356 119428 74377 119468
rect 74463 119428 74480 119468
rect 74520 119428 74529 119468
rect 74143 119405 74209 119428
rect 74295 119405 74377 119428
rect 74463 119405 74529 119428
rect 74143 119386 74529 119405
rect 89263 119491 89649 119510
rect 89263 119468 89329 119491
rect 89415 119468 89497 119491
rect 89583 119468 89649 119491
rect 89263 119428 89272 119468
rect 89312 119428 89329 119468
rect 89415 119428 89436 119468
rect 89476 119428 89497 119468
rect 89583 119428 89600 119468
rect 89640 119428 89649 119468
rect 89263 119405 89329 119428
rect 89415 119405 89497 119428
rect 89583 119405 89649 119428
rect 89263 119386 89649 119405
rect 104383 119491 104769 119510
rect 104383 119468 104449 119491
rect 104535 119468 104617 119491
rect 104703 119468 104769 119491
rect 104383 119428 104392 119468
rect 104432 119428 104449 119468
rect 104535 119428 104556 119468
rect 104596 119428 104617 119468
rect 104703 119428 104720 119468
rect 104760 119428 104769 119468
rect 104383 119405 104449 119428
rect 104535 119405 104617 119428
rect 104703 119405 104769 119428
rect 104383 119386 104769 119405
rect 119503 119491 119889 119510
rect 119503 119468 119569 119491
rect 119655 119468 119737 119491
rect 119823 119468 119889 119491
rect 119503 119428 119512 119468
rect 119552 119428 119569 119468
rect 119655 119428 119676 119468
rect 119716 119428 119737 119468
rect 119823 119428 119840 119468
rect 119880 119428 119889 119468
rect 119503 119405 119569 119428
rect 119655 119405 119737 119428
rect 119823 119405 119889 119428
rect 119503 119386 119889 119405
rect 134623 119491 135009 119510
rect 134623 119468 134689 119491
rect 134775 119468 134857 119491
rect 134943 119468 135009 119491
rect 134623 119428 134632 119468
rect 134672 119428 134689 119468
rect 134775 119428 134796 119468
rect 134836 119428 134857 119468
rect 134943 119428 134960 119468
rect 135000 119428 135009 119468
rect 134623 119405 134689 119428
rect 134775 119405 134857 119428
rect 134943 119405 135009 119428
rect 134623 119386 135009 119405
rect 149743 119491 150129 119510
rect 149743 119468 149809 119491
rect 149895 119468 149977 119491
rect 150063 119468 150129 119491
rect 149743 119428 149752 119468
rect 149792 119428 149809 119468
rect 149895 119428 149916 119468
rect 149956 119428 149977 119468
rect 150063 119428 150080 119468
rect 150120 119428 150129 119468
rect 149743 119405 149809 119428
rect 149895 119405 149977 119428
rect 150063 119405 150129 119428
rect 149743 119386 150129 119405
rect 75383 118735 75769 118754
rect 75383 118712 75449 118735
rect 75535 118712 75617 118735
rect 75703 118712 75769 118735
rect 75383 118672 75392 118712
rect 75432 118672 75449 118712
rect 75535 118672 75556 118712
rect 75596 118672 75617 118712
rect 75703 118672 75720 118712
rect 75760 118672 75769 118712
rect 75383 118649 75449 118672
rect 75535 118649 75617 118672
rect 75703 118649 75769 118672
rect 75383 118630 75769 118649
rect 90503 118735 90889 118754
rect 90503 118712 90569 118735
rect 90655 118712 90737 118735
rect 90823 118712 90889 118735
rect 90503 118672 90512 118712
rect 90552 118672 90569 118712
rect 90655 118672 90676 118712
rect 90716 118672 90737 118712
rect 90823 118672 90840 118712
rect 90880 118672 90889 118712
rect 90503 118649 90569 118672
rect 90655 118649 90737 118672
rect 90823 118649 90889 118672
rect 90503 118630 90889 118649
rect 105623 118735 106009 118754
rect 105623 118712 105689 118735
rect 105775 118712 105857 118735
rect 105943 118712 106009 118735
rect 105623 118672 105632 118712
rect 105672 118672 105689 118712
rect 105775 118672 105796 118712
rect 105836 118672 105857 118712
rect 105943 118672 105960 118712
rect 106000 118672 106009 118712
rect 105623 118649 105689 118672
rect 105775 118649 105857 118672
rect 105943 118649 106009 118672
rect 105623 118630 106009 118649
rect 120743 118735 121129 118754
rect 120743 118712 120809 118735
rect 120895 118712 120977 118735
rect 121063 118712 121129 118735
rect 120743 118672 120752 118712
rect 120792 118672 120809 118712
rect 120895 118672 120916 118712
rect 120956 118672 120977 118712
rect 121063 118672 121080 118712
rect 121120 118672 121129 118712
rect 120743 118649 120809 118672
rect 120895 118649 120977 118672
rect 121063 118649 121129 118672
rect 120743 118630 121129 118649
rect 135863 118735 136249 118754
rect 135863 118712 135929 118735
rect 136015 118712 136097 118735
rect 136183 118712 136249 118735
rect 135863 118672 135872 118712
rect 135912 118672 135929 118712
rect 136015 118672 136036 118712
rect 136076 118672 136097 118712
rect 136183 118672 136200 118712
rect 136240 118672 136249 118712
rect 135863 118649 135929 118672
rect 136015 118649 136097 118672
rect 136183 118649 136249 118672
rect 135863 118630 136249 118649
rect 150983 118735 151369 118754
rect 150983 118712 151049 118735
rect 151135 118712 151217 118735
rect 151303 118712 151369 118735
rect 150983 118672 150992 118712
rect 151032 118672 151049 118712
rect 151135 118672 151156 118712
rect 151196 118672 151217 118712
rect 151303 118672 151320 118712
rect 151360 118672 151369 118712
rect 150983 118649 151049 118672
rect 151135 118649 151217 118672
rect 151303 118649 151369 118672
rect 150983 118630 151369 118649
rect 74143 117979 74529 117998
rect 74143 117956 74209 117979
rect 74295 117956 74377 117979
rect 74463 117956 74529 117979
rect 74143 117916 74152 117956
rect 74192 117916 74209 117956
rect 74295 117916 74316 117956
rect 74356 117916 74377 117956
rect 74463 117916 74480 117956
rect 74520 117916 74529 117956
rect 74143 117893 74209 117916
rect 74295 117893 74377 117916
rect 74463 117893 74529 117916
rect 74143 117874 74529 117893
rect 89263 117979 89649 117998
rect 89263 117956 89329 117979
rect 89415 117956 89497 117979
rect 89583 117956 89649 117979
rect 89263 117916 89272 117956
rect 89312 117916 89329 117956
rect 89415 117916 89436 117956
rect 89476 117916 89497 117956
rect 89583 117916 89600 117956
rect 89640 117916 89649 117956
rect 89263 117893 89329 117916
rect 89415 117893 89497 117916
rect 89583 117893 89649 117916
rect 89263 117874 89649 117893
rect 104383 117979 104769 117998
rect 104383 117956 104449 117979
rect 104535 117956 104617 117979
rect 104703 117956 104769 117979
rect 104383 117916 104392 117956
rect 104432 117916 104449 117956
rect 104535 117916 104556 117956
rect 104596 117916 104617 117956
rect 104703 117916 104720 117956
rect 104760 117916 104769 117956
rect 104383 117893 104449 117916
rect 104535 117893 104617 117916
rect 104703 117893 104769 117916
rect 104383 117874 104769 117893
rect 119503 117979 119889 117998
rect 119503 117956 119569 117979
rect 119655 117956 119737 117979
rect 119823 117956 119889 117979
rect 119503 117916 119512 117956
rect 119552 117916 119569 117956
rect 119655 117916 119676 117956
rect 119716 117916 119737 117956
rect 119823 117916 119840 117956
rect 119880 117916 119889 117956
rect 119503 117893 119569 117916
rect 119655 117893 119737 117916
rect 119823 117893 119889 117916
rect 119503 117874 119889 117893
rect 134623 117979 135009 117998
rect 134623 117956 134689 117979
rect 134775 117956 134857 117979
rect 134943 117956 135009 117979
rect 134623 117916 134632 117956
rect 134672 117916 134689 117956
rect 134775 117916 134796 117956
rect 134836 117916 134857 117956
rect 134943 117916 134960 117956
rect 135000 117916 135009 117956
rect 134623 117893 134689 117916
rect 134775 117893 134857 117916
rect 134943 117893 135009 117916
rect 134623 117874 135009 117893
rect 149743 117979 150129 117998
rect 149743 117956 149809 117979
rect 149895 117956 149977 117979
rect 150063 117956 150129 117979
rect 149743 117916 149752 117956
rect 149792 117916 149809 117956
rect 149895 117916 149916 117956
rect 149956 117916 149977 117956
rect 150063 117916 150080 117956
rect 150120 117916 150129 117956
rect 149743 117893 149809 117916
rect 149895 117893 149977 117916
rect 150063 117893 150129 117916
rect 149743 117874 150129 117893
rect 75383 117223 75769 117242
rect 75383 117200 75449 117223
rect 75535 117200 75617 117223
rect 75703 117200 75769 117223
rect 75383 117160 75392 117200
rect 75432 117160 75449 117200
rect 75535 117160 75556 117200
rect 75596 117160 75617 117200
rect 75703 117160 75720 117200
rect 75760 117160 75769 117200
rect 75383 117137 75449 117160
rect 75535 117137 75617 117160
rect 75703 117137 75769 117160
rect 75383 117118 75769 117137
rect 90503 117223 90889 117242
rect 90503 117200 90569 117223
rect 90655 117200 90737 117223
rect 90823 117200 90889 117223
rect 90503 117160 90512 117200
rect 90552 117160 90569 117200
rect 90655 117160 90676 117200
rect 90716 117160 90737 117200
rect 90823 117160 90840 117200
rect 90880 117160 90889 117200
rect 90503 117137 90569 117160
rect 90655 117137 90737 117160
rect 90823 117137 90889 117160
rect 90503 117118 90889 117137
rect 105623 117223 106009 117242
rect 105623 117200 105689 117223
rect 105775 117200 105857 117223
rect 105943 117200 106009 117223
rect 105623 117160 105632 117200
rect 105672 117160 105689 117200
rect 105775 117160 105796 117200
rect 105836 117160 105857 117200
rect 105943 117160 105960 117200
rect 106000 117160 106009 117200
rect 105623 117137 105689 117160
rect 105775 117137 105857 117160
rect 105943 117137 106009 117160
rect 105623 117118 106009 117137
rect 120743 117223 121129 117242
rect 120743 117200 120809 117223
rect 120895 117200 120977 117223
rect 121063 117200 121129 117223
rect 120743 117160 120752 117200
rect 120792 117160 120809 117200
rect 120895 117160 120916 117200
rect 120956 117160 120977 117200
rect 121063 117160 121080 117200
rect 121120 117160 121129 117200
rect 120743 117137 120809 117160
rect 120895 117137 120977 117160
rect 121063 117137 121129 117160
rect 120743 117118 121129 117137
rect 135863 117223 136249 117242
rect 135863 117200 135929 117223
rect 136015 117200 136097 117223
rect 136183 117200 136249 117223
rect 135863 117160 135872 117200
rect 135912 117160 135929 117200
rect 136015 117160 136036 117200
rect 136076 117160 136097 117200
rect 136183 117160 136200 117200
rect 136240 117160 136249 117200
rect 135863 117137 135929 117160
rect 136015 117137 136097 117160
rect 136183 117137 136249 117160
rect 135863 117118 136249 117137
rect 150983 117223 151369 117242
rect 150983 117200 151049 117223
rect 151135 117200 151217 117223
rect 151303 117200 151369 117223
rect 150983 117160 150992 117200
rect 151032 117160 151049 117200
rect 151135 117160 151156 117200
rect 151196 117160 151217 117200
rect 151303 117160 151320 117200
rect 151360 117160 151369 117200
rect 150983 117137 151049 117160
rect 151135 117137 151217 117160
rect 151303 117137 151369 117160
rect 150983 117118 151369 117137
rect 74143 116467 74529 116486
rect 74143 116444 74209 116467
rect 74295 116444 74377 116467
rect 74463 116444 74529 116467
rect 74143 116404 74152 116444
rect 74192 116404 74209 116444
rect 74295 116404 74316 116444
rect 74356 116404 74377 116444
rect 74463 116404 74480 116444
rect 74520 116404 74529 116444
rect 74143 116381 74209 116404
rect 74295 116381 74377 116404
rect 74463 116381 74529 116404
rect 74143 116362 74529 116381
rect 89263 116467 89649 116486
rect 89263 116444 89329 116467
rect 89415 116444 89497 116467
rect 89583 116444 89649 116467
rect 89263 116404 89272 116444
rect 89312 116404 89329 116444
rect 89415 116404 89436 116444
rect 89476 116404 89497 116444
rect 89583 116404 89600 116444
rect 89640 116404 89649 116444
rect 89263 116381 89329 116404
rect 89415 116381 89497 116404
rect 89583 116381 89649 116404
rect 89263 116362 89649 116381
rect 104383 116467 104769 116486
rect 104383 116444 104449 116467
rect 104535 116444 104617 116467
rect 104703 116444 104769 116467
rect 104383 116404 104392 116444
rect 104432 116404 104449 116444
rect 104535 116404 104556 116444
rect 104596 116404 104617 116444
rect 104703 116404 104720 116444
rect 104760 116404 104769 116444
rect 104383 116381 104449 116404
rect 104535 116381 104617 116404
rect 104703 116381 104769 116404
rect 104383 116362 104769 116381
rect 119503 116467 119889 116486
rect 119503 116444 119569 116467
rect 119655 116444 119737 116467
rect 119823 116444 119889 116467
rect 119503 116404 119512 116444
rect 119552 116404 119569 116444
rect 119655 116404 119676 116444
rect 119716 116404 119737 116444
rect 119823 116404 119840 116444
rect 119880 116404 119889 116444
rect 119503 116381 119569 116404
rect 119655 116381 119737 116404
rect 119823 116381 119889 116404
rect 119503 116362 119889 116381
rect 134623 116467 135009 116486
rect 134623 116444 134689 116467
rect 134775 116444 134857 116467
rect 134943 116444 135009 116467
rect 134623 116404 134632 116444
rect 134672 116404 134689 116444
rect 134775 116404 134796 116444
rect 134836 116404 134857 116444
rect 134943 116404 134960 116444
rect 135000 116404 135009 116444
rect 134623 116381 134689 116404
rect 134775 116381 134857 116404
rect 134943 116381 135009 116404
rect 134623 116362 135009 116381
rect 149743 116467 150129 116486
rect 149743 116444 149809 116467
rect 149895 116444 149977 116467
rect 150063 116444 150129 116467
rect 149743 116404 149752 116444
rect 149792 116404 149809 116444
rect 149895 116404 149916 116444
rect 149956 116404 149977 116444
rect 150063 116404 150080 116444
rect 150120 116404 150129 116444
rect 149743 116381 149809 116404
rect 149895 116381 149977 116404
rect 150063 116381 150129 116404
rect 149743 116362 150129 116381
rect 75383 115711 75769 115730
rect 75383 115688 75449 115711
rect 75535 115688 75617 115711
rect 75703 115688 75769 115711
rect 75383 115648 75392 115688
rect 75432 115648 75449 115688
rect 75535 115648 75556 115688
rect 75596 115648 75617 115688
rect 75703 115648 75720 115688
rect 75760 115648 75769 115688
rect 75383 115625 75449 115648
rect 75535 115625 75617 115648
rect 75703 115625 75769 115648
rect 75383 115606 75769 115625
rect 90503 115711 90889 115730
rect 90503 115688 90569 115711
rect 90655 115688 90737 115711
rect 90823 115688 90889 115711
rect 90503 115648 90512 115688
rect 90552 115648 90569 115688
rect 90655 115648 90676 115688
rect 90716 115648 90737 115688
rect 90823 115648 90840 115688
rect 90880 115648 90889 115688
rect 90503 115625 90569 115648
rect 90655 115625 90737 115648
rect 90823 115625 90889 115648
rect 90503 115606 90889 115625
rect 105623 115711 106009 115730
rect 105623 115688 105689 115711
rect 105775 115688 105857 115711
rect 105943 115688 106009 115711
rect 105623 115648 105632 115688
rect 105672 115648 105689 115688
rect 105775 115648 105796 115688
rect 105836 115648 105857 115688
rect 105943 115648 105960 115688
rect 106000 115648 106009 115688
rect 105623 115625 105689 115648
rect 105775 115625 105857 115648
rect 105943 115625 106009 115648
rect 105623 115606 106009 115625
rect 120743 115711 121129 115730
rect 120743 115688 120809 115711
rect 120895 115688 120977 115711
rect 121063 115688 121129 115711
rect 120743 115648 120752 115688
rect 120792 115648 120809 115688
rect 120895 115648 120916 115688
rect 120956 115648 120977 115688
rect 121063 115648 121080 115688
rect 121120 115648 121129 115688
rect 120743 115625 120809 115648
rect 120895 115625 120977 115648
rect 121063 115625 121129 115648
rect 120743 115606 121129 115625
rect 135863 115711 136249 115730
rect 135863 115688 135929 115711
rect 136015 115688 136097 115711
rect 136183 115688 136249 115711
rect 135863 115648 135872 115688
rect 135912 115648 135929 115688
rect 136015 115648 136036 115688
rect 136076 115648 136097 115688
rect 136183 115648 136200 115688
rect 136240 115648 136249 115688
rect 135863 115625 135929 115648
rect 136015 115625 136097 115648
rect 136183 115625 136249 115648
rect 135863 115606 136249 115625
rect 150983 115711 151369 115730
rect 150983 115688 151049 115711
rect 151135 115688 151217 115711
rect 151303 115688 151369 115711
rect 150983 115648 150992 115688
rect 151032 115648 151049 115688
rect 151135 115648 151156 115688
rect 151196 115648 151217 115688
rect 151303 115648 151320 115688
rect 151360 115648 151369 115688
rect 150983 115625 151049 115648
rect 151135 115625 151217 115648
rect 151303 115625 151369 115648
rect 150983 115606 151369 115625
rect 74143 114955 74529 114974
rect 74143 114932 74209 114955
rect 74295 114932 74377 114955
rect 74463 114932 74529 114955
rect 74143 114892 74152 114932
rect 74192 114892 74209 114932
rect 74295 114892 74316 114932
rect 74356 114892 74377 114932
rect 74463 114892 74480 114932
rect 74520 114892 74529 114932
rect 74143 114869 74209 114892
rect 74295 114869 74377 114892
rect 74463 114869 74529 114892
rect 74143 114850 74529 114869
rect 89263 114955 89649 114974
rect 89263 114932 89329 114955
rect 89415 114932 89497 114955
rect 89583 114932 89649 114955
rect 89263 114892 89272 114932
rect 89312 114892 89329 114932
rect 89415 114892 89436 114932
rect 89476 114892 89497 114932
rect 89583 114892 89600 114932
rect 89640 114892 89649 114932
rect 89263 114869 89329 114892
rect 89415 114869 89497 114892
rect 89583 114869 89649 114892
rect 89263 114850 89649 114869
rect 104383 114955 104769 114974
rect 104383 114932 104449 114955
rect 104535 114932 104617 114955
rect 104703 114932 104769 114955
rect 104383 114892 104392 114932
rect 104432 114892 104449 114932
rect 104535 114892 104556 114932
rect 104596 114892 104617 114932
rect 104703 114892 104720 114932
rect 104760 114892 104769 114932
rect 104383 114869 104449 114892
rect 104535 114869 104617 114892
rect 104703 114869 104769 114892
rect 104383 114850 104769 114869
rect 119503 114955 119889 114974
rect 119503 114932 119569 114955
rect 119655 114932 119737 114955
rect 119823 114932 119889 114955
rect 119503 114892 119512 114932
rect 119552 114892 119569 114932
rect 119655 114892 119676 114932
rect 119716 114892 119737 114932
rect 119823 114892 119840 114932
rect 119880 114892 119889 114932
rect 119503 114869 119569 114892
rect 119655 114869 119737 114892
rect 119823 114869 119889 114892
rect 119503 114850 119889 114869
rect 134623 114955 135009 114974
rect 134623 114932 134689 114955
rect 134775 114932 134857 114955
rect 134943 114932 135009 114955
rect 134623 114892 134632 114932
rect 134672 114892 134689 114932
rect 134775 114892 134796 114932
rect 134836 114892 134857 114932
rect 134943 114892 134960 114932
rect 135000 114892 135009 114932
rect 134623 114869 134689 114892
rect 134775 114869 134857 114892
rect 134943 114869 135009 114892
rect 134623 114850 135009 114869
rect 149743 114955 150129 114974
rect 149743 114932 149809 114955
rect 149895 114932 149977 114955
rect 150063 114932 150129 114955
rect 149743 114892 149752 114932
rect 149792 114892 149809 114932
rect 149895 114892 149916 114932
rect 149956 114892 149977 114932
rect 150063 114892 150080 114932
rect 150120 114892 150129 114932
rect 149743 114869 149809 114892
rect 149895 114869 149977 114892
rect 150063 114869 150129 114892
rect 149743 114850 150129 114869
rect 75383 114199 75769 114218
rect 75383 114176 75449 114199
rect 75535 114176 75617 114199
rect 75703 114176 75769 114199
rect 75383 114136 75392 114176
rect 75432 114136 75449 114176
rect 75535 114136 75556 114176
rect 75596 114136 75617 114176
rect 75703 114136 75720 114176
rect 75760 114136 75769 114176
rect 75383 114113 75449 114136
rect 75535 114113 75617 114136
rect 75703 114113 75769 114136
rect 75383 114094 75769 114113
rect 90503 114199 90889 114218
rect 90503 114176 90569 114199
rect 90655 114176 90737 114199
rect 90823 114176 90889 114199
rect 90503 114136 90512 114176
rect 90552 114136 90569 114176
rect 90655 114136 90676 114176
rect 90716 114136 90737 114176
rect 90823 114136 90840 114176
rect 90880 114136 90889 114176
rect 90503 114113 90569 114136
rect 90655 114113 90737 114136
rect 90823 114113 90889 114136
rect 90503 114094 90889 114113
rect 105623 114199 106009 114218
rect 105623 114176 105689 114199
rect 105775 114176 105857 114199
rect 105943 114176 106009 114199
rect 105623 114136 105632 114176
rect 105672 114136 105689 114176
rect 105775 114136 105796 114176
rect 105836 114136 105857 114176
rect 105943 114136 105960 114176
rect 106000 114136 106009 114176
rect 105623 114113 105689 114136
rect 105775 114113 105857 114136
rect 105943 114113 106009 114136
rect 105623 114094 106009 114113
rect 120743 114199 121129 114218
rect 120743 114176 120809 114199
rect 120895 114176 120977 114199
rect 121063 114176 121129 114199
rect 120743 114136 120752 114176
rect 120792 114136 120809 114176
rect 120895 114136 120916 114176
rect 120956 114136 120977 114176
rect 121063 114136 121080 114176
rect 121120 114136 121129 114176
rect 120743 114113 120809 114136
rect 120895 114113 120977 114136
rect 121063 114113 121129 114136
rect 120743 114094 121129 114113
rect 135863 114199 136249 114218
rect 135863 114176 135929 114199
rect 136015 114176 136097 114199
rect 136183 114176 136249 114199
rect 135863 114136 135872 114176
rect 135912 114136 135929 114176
rect 136015 114136 136036 114176
rect 136076 114136 136097 114176
rect 136183 114136 136200 114176
rect 136240 114136 136249 114176
rect 135863 114113 135929 114136
rect 136015 114113 136097 114136
rect 136183 114113 136249 114136
rect 135863 114094 136249 114113
rect 150983 114199 151369 114218
rect 150983 114176 151049 114199
rect 151135 114176 151217 114199
rect 151303 114176 151369 114199
rect 150983 114136 150992 114176
rect 151032 114136 151049 114176
rect 151135 114136 151156 114176
rect 151196 114136 151217 114176
rect 151303 114136 151320 114176
rect 151360 114136 151369 114176
rect 150983 114113 151049 114136
rect 151135 114113 151217 114136
rect 151303 114113 151369 114136
rect 150983 114094 151369 114113
rect 74143 113443 74529 113462
rect 74143 113420 74209 113443
rect 74295 113420 74377 113443
rect 74463 113420 74529 113443
rect 74143 113380 74152 113420
rect 74192 113380 74209 113420
rect 74295 113380 74316 113420
rect 74356 113380 74377 113420
rect 74463 113380 74480 113420
rect 74520 113380 74529 113420
rect 74143 113357 74209 113380
rect 74295 113357 74377 113380
rect 74463 113357 74529 113380
rect 74143 113338 74529 113357
rect 89263 113443 89649 113462
rect 89263 113420 89329 113443
rect 89415 113420 89497 113443
rect 89583 113420 89649 113443
rect 89263 113380 89272 113420
rect 89312 113380 89329 113420
rect 89415 113380 89436 113420
rect 89476 113380 89497 113420
rect 89583 113380 89600 113420
rect 89640 113380 89649 113420
rect 89263 113357 89329 113380
rect 89415 113357 89497 113380
rect 89583 113357 89649 113380
rect 89263 113338 89649 113357
rect 104383 113443 104769 113462
rect 104383 113420 104449 113443
rect 104535 113420 104617 113443
rect 104703 113420 104769 113443
rect 104383 113380 104392 113420
rect 104432 113380 104449 113420
rect 104535 113380 104556 113420
rect 104596 113380 104617 113420
rect 104703 113380 104720 113420
rect 104760 113380 104769 113420
rect 104383 113357 104449 113380
rect 104535 113357 104617 113380
rect 104703 113357 104769 113380
rect 104383 113338 104769 113357
rect 119503 113443 119889 113462
rect 119503 113420 119569 113443
rect 119655 113420 119737 113443
rect 119823 113420 119889 113443
rect 119503 113380 119512 113420
rect 119552 113380 119569 113420
rect 119655 113380 119676 113420
rect 119716 113380 119737 113420
rect 119823 113380 119840 113420
rect 119880 113380 119889 113420
rect 119503 113357 119569 113380
rect 119655 113357 119737 113380
rect 119823 113357 119889 113380
rect 119503 113338 119889 113357
rect 134623 113443 135009 113462
rect 134623 113420 134689 113443
rect 134775 113420 134857 113443
rect 134943 113420 135009 113443
rect 134623 113380 134632 113420
rect 134672 113380 134689 113420
rect 134775 113380 134796 113420
rect 134836 113380 134857 113420
rect 134943 113380 134960 113420
rect 135000 113380 135009 113420
rect 134623 113357 134689 113380
rect 134775 113357 134857 113380
rect 134943 113357 135009 113380
rect 134623 113338 135009 113357
rect 149743 113443 150129 113462
rect 149743 113420 149809 113443
rect 149895 113420 149977 113443
rect 150063 113420 150129 113443
rect 149743 113380 149752 113420
rect 149792 113380 149809 113420
rect 149895 113380 149916 113420
rect 149956 113380 149977 113420
rect 150063 113380 150080 113420
rect 150120 113380 150129 113420
rect 149743 113357 149809 113380
rect 149895 113357 149977 113380
rect 150063 113357 150129 113380
rect 149743 113338 150129 113357
rect 75383 112687 75769 112706
rect 75383 112664 75449 112687
rect 75535 112664 75617 112687
rect 75703 112664 75769 112687
rect 75383 112624 75392 112664
rect 75432 112624 75449 112664
rect 75535 112624 75556 112664
rect 75596 112624 75617 112664
rect 75703 112624 75720 112664
rect 75760 112624 75769 112664
rect 75383 112601 75449 112624
rect 75535 112601 75617 112624
rect 75703 112601 75769 112624
rect 75383 112582 75769 112601
rect 90503 112687 90889 112706
rect 90503 112664 90569 112687
rect 90655 112664 90737 112687
rect 90823 112664 90889 112687
rect 90503 112624 90512 112664
rect 90552 112624 90569 112664
rect 90655 112624 90676 112664
rect 90716 112624 90737 112664
rect 90823 112624 90840 112664
rect 90880 112624 90889 112664
rect 90503 112601 90569 112624
rect 90655 112601 90737 112624
rect 90823 112601 90889 112624
rect 90503 112582 90889 112601
rect 105623 112687 106009 112706
rect 105623 112664 105689 112687
rect 105775 112664 105857 112687
rect 105943 112664 106009 112687
rect 105623 112624 105632 112664
rect 105672 112624 105689 112664
rect 105775 112624 105796 112664
rect 105836 112624 105857 112664
rect 105943 112624 105960 112664
rect 106000 112624 106009 112664
rect 105623 112601 105689 112624
rect 105775 112601 105857 112624
rect 105943 112601 106009 112624
rect 105623 112582 106009 112601
rect 120743 112687 121129 112706
rect 120743 112664 120809 112687
rect 120895 112664 120977 112687
rect 121063 112664 121129 112687
rect 120743 112624 120752 112664
rect 120792 112624 120809 112664
rect 120895 112624 120916 112664
rect 120956 112624 120977 112664
rect 121063 112624 121080 112664
rect 121120 112624 121129 112664
rect 120743 112601 120809 112624
rect 120895 112601 120977 112624
rect 121063 112601 121129 112624
rect 120743 112582 121129 112601
rect 135863 112687 136249 112706
rect 135863 112664 135929 112687
rect 136015 112664 136097 112687
rect 136183 112664 136249 112687
rect 135863 112624 135872 112664
rect 135912 112624 135929 112664
rect 136015 112624 136036 112664
rect 136076 112624 136097 112664
rect 136183 112624 136200 112664
rect 136240 112624 136249 112664
rect 135863 112601 135929 112624
rect 136015 112601 136097 112624
rect 136183 112601 136249 112624
rect 135863 112582 136249 112601
rect 150983 112687 151369 112706
rect 150983 112664 151049 112687
rect 151135 112664 151217 112687
rect 151303 112664 151369 112687
rect 150983 112624 150992 112664
rect 151032 112624 151049 112664
rect 151135 112624 151156 112664
rect 151196 112624 151217 112664
rect 151303 112624 151320 112664
rect 151360 112624 151369 112664
rect 150983 112601 151049 112624
rect 151135 112601 151217 112624
rect 151303 112601 151369 112624
rect 150983 112582 151369 112601
rect 74143 111931 74529 111950
rect 74143 111908 74209 111931
rect 74295 111908 74377 111931
rect 74463 111908 74529 111931
rect 74143 111868 74152 111908
rect 74192 111868 74209 111908
rect 74295 111868 74316 111908
rect 74356 111868 74377 111908
rect 74463 111868 74480 111908
rect 74520 111868 74529 111908
rect 74143 111845 74209 111868
rect 74295 111845 74377 111868
rect 74463 111845 74529 111868
rect 74143 111826 74529 111845
rect 89263 111931 89649 111950
rect 89263 111908 89329 111931
rect 89415 111908 89497 111931
rect 89583 111908 89649 111931
rect 89263 111868 89272 111908
rect 89312 111868 89329 111908
rect 89415 111868 89436 111908
rect 89476 111868 89497 111908
rect 89583 111868 89600 111908
rect 89640 111868 89649 111908
rect 89263 111845 89329 111868
rect 89415 111845 89497 111868
rect 89583 111845 89649 111868
rect 89263 111826 89649 111845
rect 104383 111931 104769 111950
rect 104383 111908 104449 111931
rect 104535 111908 104617 111931
rect 104703 111908 104769 111931
rect 104383 111868 104392 111908
rect 104432 111868 104449 111908
rect 104535 111868 104556 111908
rect 104596 111868 104617 111908
rect 104703 111868 104720 111908
rect 104760 111868 104769 111908
rect 104383 111845 104449 111868
rect 104535 111845 104617 111868
rect 104703 111845 104769 111868
rect 104383 111826 104769 111845
rect 119503 111931 119889 111950
rect 119503 111908 119569 111931
rect 119655 111908 119737 111931
rect 119823 111908 119889 111931
rect 119503 111868 119512 111908
rect 119552 111868 119569 111908
rect 119655 111868 119676 111908
rect 119716 111868 119737 111908
rect 119823 111868 119840 111908
rect 119880 111868 119889 111908
rect 119503 111845 119569 111868
rect 119655 111845 119737 111868
rect 119823 111845 119889 111868
rect 119503 111826 119889 111845
rect 134623 111931 135009 111950
rect 134623 111908 134689 111931
rect 134775 111908 134857 111931
rect 134943 111908 135009 111931
rect 134623 111868 134632 111908
rect 134672 111868 134689 111908
rect 134775 111868 134796 111908
rect 134836 111868 134857 111908
rect 134943 111868 134960 111908
rect 135000 111868 135009 111908
rect 134623 111845 134689 111868
rect 134775 111845 134857 111868
rect 134943 111845 135009 111868
rect 134623 111826 135009 111845
rect 149743 111931 150129 111950
rect 149743 111908 149809 111931
rect 149895 111908 149977 111931
rect 150063 111908 150129 111931
rect 149743 111868 149752 111908
rect 149792 111868 149809 111908
rect 149895 111868 149916 111908
rect 149956 111868 149977 111908
rect 150063 111868 150080 111908
rect 150120 111868 150129 111908
rect 149743 111845 149809 111868
rect 149895 111845 149977 111868
rect 150063 111845 150129 111868
rect 149743 111826 150129 111845
rect 75383 111175 75769 111194
rect 75383 111152 75449 111175
rect 75535 111152 75617 111175
rect 75703 111152 75769 111175
rect 75383 111112 75392 111152
rect 75432 111112 75449 111152
rect 75535 111112 75556 111152
rect 75596 111112 75617 111152
rect 75703 111112 75720 111152
rect 75760 111112 75769 111152
rect 75383 111089 75449 111112
rect 75535 111089 75617 111112
rect 75703 111089 75769 111112
rect 75383 111070 75769 111089
rect 90503 111175 90889 111194
rect 90503 111152 90569 111175
rect 90655 111152 90737 111175
rect 90823 111152 90889 111175
rect 90503 111112 90512 111152
rect 90552 111112 90569 111152
rect 90655 111112 90676 111152
rect 90716 111112 90737 111152
rect 90823 111112 90840 111152
rect 90880 111112 90889 111152
rect 90503 111089 90569 111112
rect 90655 111089 90737 111112
rect 90823 111089 90889 111112
rect 90503 111070 90889 111089
rect 105623 111175 106009 111194
rect 105623 111152 105689 111175
rect 105775 111152 105857 111175
rect 105943 111152 106009 111175
rect 105623 111112 105632 111152
rect 105672 111112 105689 111152
rect 105775 111112 105796 111152
rect 105836 111112 105857 111152
rect 105943 111112 105960 111152
rect 106000 111112 106009 111152
rect 105623 111089 105689 111112
rect 105775 111089 105857 111112
rect 105943 111089 106009 111112
rect 105623 111070 106009 111089
rect 120743 111175 121129 111194
rect 120743 111152 120809 111175
rect 120895 111152 120977 111175
rect 121063 111152 121129 111175
rect 120743 111112 120752 111152
rect 120792 111112 120809 111152
rect 120895 111112 120916 111152
rect 120956 111112 120977 111152
rect 121063 111112 121080 111152
rect 121120 111112 121129 111152
rect 120743 111089 120809 111112
rect 120895 111089 120977 111112
rect 121063 111089 121129 111112
rect 120743 111070 121129 111089
rect 135863 111175 136249 111194
rect 135863 111152 135929 111175
rect 136015 111152 136097 111175
rect 136183 111152 136249 111175
rect 135863 111112 135872 111152
rect 135912 111112 135929 111152
rect 136015 111112 136036 111152
rect 136076 111112 136097 111152
rect 136183 111112 136200 111152
rect 136240 111112 136249 111152
rect 135863 111089 135929 111112
rect 136015 111089 136097 111112
rect 136183 111089 136249 111112
rect 135863 111070 136249 111089
rect 150983 111175 151369 111194
rect 150983 111152 151049 111175
rect 151135 111152 151217 111175
rect 151303 111152 151369 111175
rect 150983 111112 150992 111152
rect 151032 111112 151049 111152
rect 151135 111112 151156 111152
rect 151196 111112 151217 111152
rect 151303 111112 151320 111152
rect 151360 111112 151369 111152
rect 150983 111089 151049 111112
rect 151135 111089 151217 111112
rect 151303 111089 151369 111112
rect 150983 111070 151369 111089
rect 74143 110419 74529 110438
rect 74143 110396 74209 110419
rect 74295 110396 74377 110419
rect 74463 110396 74529 110419
rect 74143 110356 74152 110396
rect 74192 110356 74209 110396
rect 74295 110356 74316 110396
rect 74356 110356 74377 110396
rect 74463 110356 74480 110396
rect 74520 110356 74529 110396
rect 74143 110333 74209 110356
rect 74295 110333 74377 110356
rect 74463 110333 74529 110356
rect 74143 110314 74529 110333
rect 89263 110419 89649 110438
rect 89263 110396 89329 110419
rect 89415 110396 89497 110419
rect 89583 110396 89649 110419
rect 89263 110356 89272 110396
rect 89312 110356 89329 110396
rect 89415 110356 89436 110396
rect 89476 110356 89497 110396
rect 89583 110356 89600 110396
rect 89640 110356 89649 110396
rect 89263 110333 89329 110356
rect 89415 110333 89497 110356
rect 89583 110333 89649 110356
rect 89263 110314 89649 110333
rect 104383 110419 104769 110438
rect 104383 110396 104449 110419
rect 104535 110396 104617 110419
rect 104703 110396 104769 110419
rect 104383 110356 104392 110396
rect 104432 110356 104449 110396
rect 104535 110356 104556 110396
rect 104596 110356 104617 110396
rect 104703 110356 104720 110396
rect 104760 110356 104769 110396
rect 104383 110333 104449 110356
rect 104535 110333 104617 110356
rect 104703 110333 104769 110356
rect 104383 110314 104769 110333
rect 119503 110419 119889 110438
rect 119503 110396 119569 110419
rect 119655 110396 119737 110419
rect 119823 110396 119889 110419
rect 119503 110356 119512 110396
rect 119552 110356 119569 110396
rect 119655 110356 119676 110396
rect 119716 110356 119737 110396
rect 119823 110356 119840 110396
rect 119880 110356 119889 110396
rect 119503 110333 119569 110356
rect 119655 110333 119737 110356
rect 119823 110333 119889 110356
rect 119503 110314 119889 110333
rect 134623 110419 135009 110438
rect 134623 110396 134689 110419
rect 134775 110396 134857 110419
rect 134943 110396 135009 110419
rect 134623 110356 134632 110396
rect 134672 110356 134689 110396
rect 134775 110356 134796 110396
rect 134836 110356 134857 110396
rect 134943 110356 134960 110396
rect 135000 110356 135009 110396
rect 134623 110333 134689 110356
rect 134775 110333 134857 110356
rect 134943 110333 135009 110356
rect 134623 110314 135009 110333
rect 149743 110419 150129 110438
rect 149743 110396 149809 110419
rect 149895 110396 149977 110419
rect 150063 110396 150129 110419
rect 149743 110356 149752 110396
rect 149792 110356 149809 110396
rect 149895 110356 149916 110396
rect 149956 110356 149977 110396
rect 150063 110356 150080 110396
rect 150120 110356 150129 110396
rect 149743 110333 149809 110356
rect 149895 110333 149977 110356
rect 150063 110333 150129 110356
rect 149743 110314 150129 110333
rect 75383 109663 75769 109682
rect 75383 109640 75449 109663
rect 75535 109640 75617 109663
rect 75703 109640 75769 109663
rect 75383 109600 75392 109640
rect 75432 109600 75449 109640
rect 75535 109600 75556 109640
rect 75596 109600 75617 109640
rect 75703 109600 75720 109640
rect 75760 109600 75769 109640
rect 75383 109577 75449 109600
rect 75535 109577 75617 109600
rect 75703 109577 75769 109600
rect 75383 109558 75769 109577
rect 90503 109663 90889 109682
rect 90503 109640 90569 109663
rect 90655 109640 90737 109663
rect 90823 109640 90889 109663
rect 90503 109600 90512 109640
rect 90552 109600 90569 109640
rect 90655 109600 90676 109640
rect 90716 109600 90737 109640
rect 90823 109600 90840 109640
rect 90880 109600 90889 109640
rect 90503 109577 90569 109600
rect 90655 109577 90737 109600
rect 90823 109577 90889 109600
rect 90503 109558 90889 109577
rect 105623 109663 106009 109682
rect 105623 109640 105689 109663
rect 105775 109640 105857 109663
rect 105943 109640 106009 109663
rect 105623 109600 105632 109640
rect 105672 109600 105689 109640
rect 105775 109600 105796 109640
rect 105836 109600 105857 109640
rect 105943 109600 105960 109640
rect 106000 109600 106009 109640
rect 105623 109577 105689 109600
rect 105775 109577 105857 109600
rect 105943 109577 106009 109600
rect 105623 109558 106009 109577
rect 120743 109663 121129 109682
rect 120743 109640 120809 109663
rect 120895 109640 120977 109663
rect 121063 109640 121129 109663
rect 120743 109600 120752 109640
rect 120792 109600 120809 109640
rect 120895 109600 120916 109640
rect 120956 109600 120977 109640
rect 121063 109600 121080 109640
rect 121120 109600 121129 109640
rect 120743 109577 120809 109600
rect 120895 109577 120977 109600
rect 121063 109577 121129 109600
rect 120743 109558 121129 109577
rect 135863 109663 136249 109682
rect 135863 109640 135929 109663
rect 136015 109640 136097 109663
rect 136183 109640 136249 109663
rect 135863 109600 135872 109640
rect 135912 109600 135929 109640
rect 136015 109600 136036 109640
rect 136076 109600 136097 109640
rect 136183 109600 136200 109640
rect 136240 109600 136249 109640
rect 135863 109577 135929 109600
rect 136015 109577 136097 109600
rect 136183 109577 136249 109600
rect 135863 109558 136249 109577
rect 150983 109663 151369 109682
rect 150983 109640 151049 109663
rect 151135 109640 151217 109663
rect 151303 109640 151369 109663
rect 150983 109600 150992 109640
rect 151032 109600 151049 109640
rect 151135 109600 151156 109640
rect 151196 109600 151217 109640
rect 151303 109600 151320 109640
rect 151360 109600 151369 109640
rect 150983 109577 151049 109600
rect 151135 109577 151217 109600
rect 151303 109577 151369 109600
rect 150983 109558 151369 109577
rect 74143 108907 74529 108926
rect 74143 108884 74209 108907
rect 74295 108884 74377 108907
rect 74463 108884 74529 108907
rect 74143 108844 74152 108884
rect 74192 108844 74209 108884
rect 74295 108844 74316 108884
rect 74356 108844 74377 108884
rect 74463 108844 74480 108884
rect 74520 108844 74529 108884
rect 74143 108821 74209 108844
rect 74295 108821 74377 108844
rect 74463 108821 74529 108844
rect 74143 108802 74529 108821
rect 89263 108907 89649 108926
rect 89263 108884 89329 108907
rect 89415 108884 89497 108907
rect 89583 108884 89649 108907
rect 89263 108844 89272 108884
rect 89312 108844 89329 108884
rect 89415 108844 89436 108884
rect 89476 108844 89497 108884
rect 89583 108844 89600 108884
rect 89640 108844 89649 108884
rect 89263 108821 89329 108844
rect 89415 108821 89497 108844
rect 89583 108821 89649 108844
rect 89263 108802 89649 108821
rect 104383 108907 104769 108926
rect 104383 108884 104449 108907
rect 104535 108884 104617 108907
rect 104703 108884 104769 108907
rect 104383 108844 104392 108884
rect 104432 108844 104449 108884
rect 104535 108844 104556 108884
rect 104596 108844 104617 108884
rect 104703 108844 104720 108884
rect 104760 108844 104769 108884
rect 104383 108821 104449 108844
rect 104535 108821 104617 108844
rect 104703 108821 104769 108844
rect 104383 108802 104769 108821
rect 119503 108907 119889 108926
rect 119503 108884 119569 108907
rect 119655 108884 119737 108907
rect 119823 108884 119889 108907
rect 119503 108844 119512 108884
rect 119552 108844 119569 108884
rect 119655 108844 119676 108884
rect 119716 108844 119737 108884
rect 119823 108844 119840 108884
rect 119880 108844 119889 108884
rect 119503 108821 119569 108844
rect 119655 108821 119737 108844
rect 119823 108821 119889 108844
rect 119503 108802 119889 108821
rect 134623 108907 135009 108926
rect 134623 108884 134689 108907
rect 134775 108884 134857 108907
rect 134943 108884 135009 108907
rect 134623 108844 134632 108884
rect 134672 108844 134689 108884
rect 134775 108844 134796 108884
rect 134836 108844 134857 108884
rect 134943 108844 134960 108884
rect 135000 108844 135009 108884
rect 134623 108821 134689 108844
rect 134775 108821 134857 108844
rect 134943 108821 135009 108844
rect 134623 108802 135009 108821
rect 149743 108907 150129 108926
rect 149743 108884 149809 108907
rect 149895 108884 149977 108907
rect 150063 108884 150129 108907
rect 149743 108844 149752 108884
rect 149792 108844 149809 108884
rect 149895 108844 149916 108884
rect 149956 108844 149977 108884
rect 150063 108844 150080 108884
rect 150120 108844 150129 108884
rect 149743 108821 149809 108844
rect 149895 108821 149977 108844
rect 150063 108821 150129 108844
rect 149743 108802 150129 108821
rect 75383 108151 75769 108170
rect 75383 108128 75449 108151
rect 75535 108128 75617 108151
rect 75703 108128 75769 108151
rect 75383 108088 75392 108128
rect 75432 108088 75449 108128
rect 75535 108088 75556 108128
rect 75596 108088 75617 108128
rect 75703 108088 75720 108128
rect 75760 108088 75769 108128
rect 75383 108065 75449 108088
rect 75535 108065 75617 108088
rect 75703 108065 75769 108088
rect 75383 108046 75769 108065
rect 90503 108151 90889 108170
rect 90503 108128 90569 108151
rect 90655 108128 90737 108151
rect 90823 108128 90889 108151
rect 90503 108088 90512 108128
rect 90552 108088 90569 108128
rect 90655 108088 90676 108128
rect 90716 108088 90737 108128
rect 90823 108088 90840 108128
rect 90880 108088 90889 108128
rect 90503 108065 90569 108088
rect 90655 108065 90737 108088
rect 90823 108065 90889 108088
rect 90503 108046 90889 108065
rect 105623 108151 106009 108170
rect 105623 108128 105689 108151
rect 105775 108128 105857 108151
rect 105943 108128 106009 108151
rect 105623 108088 105632 108128
rect 105672 108088 105689 108128
rect 105775 108088 105796 108128
rect 105836 108088 105857 108128
rect 105943 108088 105960 108128
rect 106000 108088 106009 108128
rect 105623 108065 105689 108088
rect 105775 108065 105857 108088
rect 105943 108065 106009 108088
rect 105623 108046 106009 108065
rect 120743 108151 121129 108170
rect 120743 108128 120809 108151
rect 120895 108128 120977 108151
rect 121063 108128 121129 108151
rect 120743 108088 120752 108128
rect 120792 108088 120809 108128
rect 120895 108088 120916 108128
rect 120956 108088 120977 108128
rect 121063 108088 121080 108128
rect 121120 108088 121129 108128
rect 120743 108065 120809 108088
rect 120895 108065 120977 108088
rect 121063 108065 121129 108088
rect 120743 108046 121129 108065
rect 135863 108151 136249 108170
rect 135863 108128 135929 108151
rect 136015 108128 136097 108151
rect 136183 108128 136249 108151
rect 135863 108088 135872 108128
rect 135912 108088 135929 108128
rect 136015 108088 136036 108128
rect 136076 108088 136097 108128
rect 136183 108088 136200 108128
rect 136240 108088 136249 108128
rect 135863 108065 135929 108088
rect 136015 108065 136097 108088
rect 136183 108065 136249 108088
rect 135863 108046 136249 108065
rect 150983 108151 151369 108170
rect 150983 108128 151049 108151
rect 151135 108128 151217 108151
rect 151303 108128 151369 108151
rect 150983 108088 150992 108128
rect 151032 108088 151049 108128
rect 151135 108088 151156 108128
rect 151196 108088 151217 108128
rect 151303 108088 151320 108128
rect 151360 108088 151369 108128
rect 150983 108065 151049 108088
rect 151135 108065 151217 108088
rect 151303 108065 151369 108088
rect 150983 108046 151369 108065
rect 74143 107395 74529 107414
rect 74143 107372 74209 107395
rect 74295 107372 74377 107395
rect 74463 107372 74529 107395
rect 74143 107332 74152 107372
rect 74192 107332 74209 107372
rect 74295 107332 74316 107372
rect 74356 107332 74377 107372
rect 74463 107332 74480 107372
rect 74520 107332 74529 107372
rect 74143 107309 74209 107332
rect 74295 107309 74377 107332
rect 74463 107309 74529 107332
rect 74143 107290 74529 107309
rect 89263 107395 89649 107414
rect 89263 107372 89329 107395
rect 89415 107372 89497 107395
rect 89583 107372 89649 107395
rect 89263 107332 89272 107372
rect 89312 107332 89329 107372
rect 89415 107332 89436 107372
rect 89476 107332 89497 107372
rect 89583 107332 89600 107372
rect 89640 107332 89649 107372
rect 89263 107309 89329 107332
rect 89415 107309 89497 107332
rect 89583 107309 89649 107332
rect 89263 107290 89649 107309
rect 104383 107395 104769 107414
rect 104383 107372 104449 107395
rect 104535 107372 104617 107395
rect 104703 107372 104769 107395
rect 104383 107332 104392 107372
rect 104432 107332 104449 107372
rect 104535 107332 104556 107372
rect 104596 107332 104617 107372
rect 104703 107332 104720 107372
rect 104760 107332 104769 107372
rect 104383 107309 104449 107332
rect 104535 107309 104617 107332
rect 104703 107309 104769 107332
rect 104383 107290 104769 107309
rect 119503 107395 119889 107414
rect 119503 107372 119569 107395
rect 119655 107372 119737 107395
rect 119823 107372 119889 107395
rect 119503 107332 119512 107372
rect 119552 107332 119569 107372
rect 119655 107332 119676 107372
rect 119716 107332 119737 107372
rect 119823 107332 119840 107372
rect 119880 107332 119889 107372
rect 119503 107309 119569 107332
rect 119655 107309 119737 107332
rect 119823 107309 119889 107332
rect 119503 107290 119889 107309
rect 134623 107395 135009 107414
rect 134623 107372 134689 107395
rect 134775 107372 134857 107395
rect 134943 107372 135009 107395
rect 134623 107332 134632 107372
rect 134672 107332 134689 107372
rect 134775 107332 134796 107372
rect 134836 107332 134857 107372
rect 134943 107332 134960 107372
rect 135000 107332 135009 107372
rect 134623 107309 134689 107332
rect 134775 107309 134857 107332
rect 134943 107309 135009 107332
rect 134623 107290 135009 107309
rect 149743 107395 150129 107414
rect 149743 107372 149809 107395
rect 149895 107372 149977 107395
rect 150063 107372 150129 107395
rect 149743 107332 149752 107372
rect 149792 107332 149809 107372
rect 149895 107332 149916 107372
rect 149956 107332 149977 107372
rect 150063 107332 150080 107372
rect 150120 107332 150129 107372
rect 149743 107309 149809 107332
rect 149895 107309 149977 107332
rect 150063 107309 150129 107332
rect 149743 107290 150129 107309
rect 75383 106639 75769 106658
rect 75383 106616 75449 106639
rect 75535 106616 75617 106639
rect 75703 106616 75769 106639
rect 75383 106576 75392 106616
rect 75432 106576 75449 106616
rect 75535 106576 75556 106616
rect 75596 106576 75617 106616
rect 75703 106576 75720 106616
rect 75760 106576 75769 106616
rect 75383 106553 75449 106576
rect 75535 106553 75617 106576
rect 75703 106553 75769 106576
rect 75383 106534 75769 106553
rect 90503 106639 90889 106658
rect 90503 106616 90569 106639
rect 90655 106616 90737 106639
rect 90823 106616 90889 106639
rect 90503 106576 90512 106616
rect 90552 106576 90569 106616
rect 90655 106576 90676 106616
rect 90716 106576 90737 106616
rect 90823 106576 90840 106616
rect 90880 106576 90889 106616
rect 90503 106553 90569 106576
rect 90655 106553 90737 106576
rect 90823 106553 90889 106576
rect 90503 106534 90889 106553
rect 105623 106639 106009 106658
rect 105623 106616 105689 106639
rect 105775 106616 105857 106639
rect 105943 106616 106009 106639
rect 105623 106576 105632 106616
rect 105672 106576 105689 106616
rect 105775 106576 105796 106616
rect 105836 106576 105857 106616
rect 105943 106576 105960 106616
rect 106000 106576 106009 106616
rect 105623 106553 105689 106576
rect 105775 106553 105857 106576
rect 105943 106553 106009 106576
rect 105623 106534 106009 106553
rect 120743 106639 121129 106658
rect 120743 106616 120809 106639
rect 120895 106616 120977 106639
rect 121063 106616 121129 106639
rect 120743 106576 120752 106616
rect 120792 106576 120809 106616
rect 120895 106576 120916 106616
rect 120956 106576 120977 106616
rect 121063 106576 121080 106616
rect 121120 106576 121129 106616
rect 120743 106553 120809 106576
rect 120895 106553 120977 106576
rect 121063 106553 121129 106576
rect 120743 106534 121129 106553
rect 135863 106639 136249 106658
rect 135863 106616 135929 106639
rect 136015 106616 136097 106639
rect 136183 106616 136249 106639
rect 135863 106576 135872 106616
rect 135912 106576 135929 106616
rect 136015 106576 136036 106616
rect 136076 106576 136097 106616
rect 136183 106576 136200 106616
rect 136240 106576 136249 106616
rect 135863 106553 135929 106576
rect 136015 106553 136097 106576
rect 136183 106553 136249 106576
rect 135863 106534 136249 106553
rect 150983 106639 151369 106658
rect 150983 106616 151049 106639
rect 151135 106616 151217 106639
rect 151303 106616 151369 106639
rect 150983 106576 150992 106616
rect 151032 106576 151049 106616
rect 151135 106576 151156 106616
rect 151196 106576 151217 106616
rect 151303 106576 151320 106616
rect 151360 106576 151369 106616
rect 150983 106553 151049 106576
rect 151135 106553 151217 106576
rect 151303 106553 151369 106576
rect 150983 106534 151369 106553
rect 74143 105883 74529 105902
rect 74143 105860 74209 105883
rect 74295 105860 74377 105883
rect 74463 105860 74529 105883
rect 74143 105820 74152 105860
rect 74192 105820 74209 105860
rect 74295 105820 74316 105860
rect 74356 105820 74377 105860
rect 74463 105820 74480 105860
rect 74520 105820 74529 105860
rect 74143 105797 74209 105820
rect 74295 105797 74377 105820
rect 74463 105797 74529 105820
rect 74143 105778 74529 105797
rect 89263 105883 89649 105902
rect 89263 105860 89329 105883
rect 89415 105860 89497 105883
rect 89583 105860 89649 105883
rect 89263 105820 89272 105860
rect 89312 105820 89329 105860
rect 89415 105820 89436 105860
rect 89476 105820 89497 105860
rect 89583 105820 89600 105860
rect 89640 105820 89649 105860
rect 89263 105797 89329 105820
rect 89415 105797 89497 105820
rect 89583 105797 89649 105820
rect 89263 105778 89649 105797
rect 104383 105883 104769 105902
rect 104383 105860 104449 105883
rect 104535 105860 104617 105883
rect 104703 105860 104769 105883
rect 104383 105820 104392 105860
rect 104432 105820 104449 105860
rect 104535 105820 104556 105860
rect 104596 105820 104617 105860
rect 104703 105820 104720 105860
rect 104760 105820 104769 105860
rect 104383 105797 104449 105820
rect 104535 105797 104617 105820
rect 104703 105797 104769 105820
rect 104383 105778 104769 105797
rect 119503 105883 119889 105902
rect 119503 105860 119569 105883
rect 119655 105860 119737 105883
rect 119823 105860 119889 105883
rect 119503 105820 119512 105860
rect 119552 105820 119569 105860
rect 119655 105820 119676 105860
rect 119716 105820 119737 105860
rect 119823 105820 119840 105860
rect 119880 105820 119889 105860
rect 119503 105797 119569 105820
rect 119655 105797 119737 105820
rect 119823 105797 119889 105820
rect 119503 105778 119889 105797
rect 134623 105883 135009 105902
rect 134623 105860 134689 105883
rect 134775 105860 134857 105883
rect 134943 105860 135009 105883
rect 134623 105820 134632 105860
rect 134672 105820 134689 105860
rect 134775 105820 134796 105860
rect 134836 105820 134857 105860
rect 134943 105820 134960 105860
rect 135000 105820 135009 105860
rect 134623 105797 134689 105820
rect 134775 105797 134857 105820
rect 134943 105797 135009 105820
rect 134623 105778 135009 105797
rect 149743 105883 150129 105902
rect 149743 105860 149809 105883
rect 149895 105860 149977 105883
rect 150063 105860 150129 105883
rect 149743 105820 149752 105860
rect 149792 105820 149809 105860
rect 149895 105820 149916 105860
rect 149956 105820 149977 105860
rect 150063 105820 150080 105860
rect 150120 105820 150129 105860
rect 149743 105797 149809 105820
rect 149895 105797 149977 105820
rect 150063 105797 150129 105820
rect 149743 105778 150129 105797
rect 75383 105127 75769 105146
rect 75383 105104 75449 105127
rect 75535 105104 75617 105127
rect 75703 105104 75769 105127
rect 75383 105064 75392 105104
rect 75432 105064 75449 105104
rect 75535 105064 75556 105104
rect 75596 105064 75617 105104
rect 75703 105064 75720 105104
rect 75760 105064 75769 105104
rect 75383 105041 75449 105064
rect 75535 105041 75617 105064
rect 75703 105041 75769 105064
rect 75383 105022 75769 105041
rect 90503 105127 90889 105146
rect 90503 105104 90569 105127
rect 90655 105104 90737 105127
rect 90823 105104 90889 105127
rect 90503 105064 90512 105104
rect 90552 105064 90569 105104
rect 90655 105064 90676 105104
rect 90716 105064 90737 105104
rect 90823 105064 90840 105104
rect 90880 105064 90889 105104
rect 90503 105041 90569 105064
rect 90655 105041 90737 105064
rect 90823 105041 90889 105064
rect 90503 105022 90889 105041
rect 105623 105127 106009 105146
rect 105623 105104 105689 105127
rect 105775 105104 105857 105127
rect 105943 105104 106009 105127
rect 105623 105064 105632 105104
rect 105672 105064 105689 105104
rect 105775 105064 105796 105104
rect 105836 105064 105857 105104
rect 105943 105064 105960 105104
rect 106000 105064 106009 105104
rect 105623 105041 105689 105064
rect 105775 105041 105857 105064
rect 105943 105041 106009 105064
rect 105623 105022 106009 105041
rect 120743 105127 121129 105146
rect 120743 105104 120809 105127
rect 120895 105104 120977 105127
rect 121063 105104 121129 105127
rect 120743 105064 120752 105104
rect 120792 105064 120809 105104
rect 120895 105064 120916 105104
rect 120956 105064 120977 105104
rect 121063 105064 121080 105104
rect 121120 105064 121129 105104
rect 120743 105041 120809 105064
rect 120895 105041 120977 105064
rect 121063 105041 121129 105064
rect 120743 105022 121129 105041
rect 135863 105127 136249 105146
rect 135863 105104 135929 105127
rect 136015 105104 136097 105127
rect 136183 105104 136249 105127
rect 135863 105064 135872 105104
rect 135912 105064 135929 105104
rect 136015 105064 136036 105104
rect 136076 105064 136097 105104
rect 136183 105064 136200 105104
rect 136240 105064 136249 105104
rect 135863 105041 135929 105064
rect 136015 105041 136097 105064
rect 136183 105041 136249 105064
rect 135863 105022 136249 105041
rect 150983 105127 151369 105146
rect 150983 105104 151049 105127
rect 151135 105104 151217 105127
rect 151303 105104 151369 105127
rect 150983 105064 150992 105104
rect 151032 105064 151049 105104
rect 151135 105064 151156 105104
rect 151196 105064 151217 105104
rect 151303 105064 151320 105104
rect 151360 105064 151369 105104
rect 150983 105041 151049 105064
rect 151135 105041 151217 105064
rect 151303 105041 151369 105064
rect 150983 105022 151369 105041
rect 74143 104371 74529 104390
rect 74143 104348 74209 104371
rect 74295 104348 74377 104371
rect 74463 104348 74529 104371
rect 74143 104308 74152 104348
rect 74192 104308 74209 104348
rect 74295 104308 74316 104348
rect 74356 104308 74377 104348
rect 74463 104308 74480 104348
rect 74520 104308 74529 104348
rect 74143 104285 74209 104308
rect 74295 104285 74377 104308
rect 74463 104285 74529 104308
rect 74143 104266 74529 104285
rect 89263 104371 89649 104390
rect 89263 104348 89329 104371
rect 89415 104348 89497 104371
rect 89583 104348 89649 104371
rect 89263 104308 89272 104348
rect 89312 104308 89329 104348
rect 89415 104308 89436 104348
rect 89476 104308 89497 104348
rect 89583 104308 89600 104348
rect 89640 104308 89649 104348
rect 89263 104285 89329 104308
rect 89415 104285 89497 104308
rect 89583 104285 89649 104308
rect 89263 104266 89649 104285
rect 104383 104371 104769 104390
rect 104383 104348 104449 104371
rect 104535 104348 104617 104371
rect 104703 104348 104769 104371
rect 104383 104308 104392 104348
rect 104432 104308 104449 104348
rect 104535 104308 104556 104348
rect 104596 104308 104617 104348
rect 104703 104308 104720 104348
rect 104760 104308 104769 104348
rect 104383 104285 104449 104308
rect 104535 104285 104617 104308
rect 104703 104285 104769 104308
rect 104383 104266 104769 104285
rect 119503 104371 119889 104390
rect 119503 104348 119569 104371
rect 119655 104348 119737 104371
rect 119823 104348 119889 104371
rect 119503 104308 119512 104348
rect 119552 104308 119569 104348
rect 119655 104308 119676 104348
rect 119716 104308 119737 104348
rect 119823 104308 119840 104348
rect 119880 104308 119889 104348
rect 119503 104285 119569 104308
rect 119655 104285 119737 104308
rect 119823 104285 119889 104308
rect 119503 104266 119889 104285
rect 134623 104371 135009 104390
rect 134623 104348 134689 104371
rect 134775 104348 134857 104371
rect 134943 104348 135009 104371
rect 134623 104308 134632 104348
rect 134672 104308 134689 104348
rect 134775 104308 134796 104348
rect 134836 104308 134857 104348
rect 134943 104308 134960 104348
rect 135000 104308 135009 104348
rect 134623 104285 134689 104308
rect 134775 104285 134857 104308
rect 134943 104285 135009 104308
rect 134623 104266 135009 104285
rect 149743 104371 150129 104390
rect 149743 104348 149809 104371
rect 149895 104348 149977 104371
rect 150063 104348 150129 104371
rect 149743 104308 149752 104348
rect 149792 104308 149809 104348
rect 149895 104308 149916 104348
rect 149956 104308 149977 104348
rect 150063 104308 150080 104348
rect 150120 104308 150129 104348
rect 149743 104285 149809 104308
rect 149895 104285 149977 104308
rect 150063 104285 150129 104308
rect 149743 104266 150129 104285
rect 75383 103615 75769 103634
rect 75383 103592 75449 103615
rect 75535 103592 75617 103615
rect 75703 103592 75769 103615
rect 75383 103552 75392 103592
rect 75432 103552 75449 103592
rect 75535 103552 75556 103592
rect 75596 103552 75617 103592
rect 75703 103552 75720 103592
rect 75760 103552 75769 103592
rect 75383 103529 75449 103552
rect 75535 103529 75617 103552
rect 75703 103529 75769 103552
rect 75383 103510 75769 103529
rect 90503 103615 90889 103634
rect 90503 103592 90569 103615
rect 90655 103592 90737 103615
rect 90823 103592 90889 103615
rect 90503 103552 90512 103592
rect 90552 103552 90569 103592
rect 90655 103552 90676 103592
rect 90716 103552 90737 103592
rect 90823 103552 90840 103592
rect 90880 103552 90889 103592
rect 90503 103529 90569 103552
rect 90655 103529 90737 103552
rect 90823 103529 90889 103552
rect 90503 103510 90889 103529
rect 105623 103615 106009 103634
rect 105623 103592 105689 103615
rect 105775 103592 105857 103615
rect 105943 103592 106009 103615
rect 105623 103552 105632 103592
rect 105672 103552 105689 103592
rect 105775 103552 105796 103592
rect 105836 103552 105857 103592
rect 105943 103552 105960 103592
rect 106000 103552 106009 103592
rect 105623 103529 105689 103552
rect 105775 103529 105857 103552
rect 105943 103529 106009 103552
rect 105623 103510 106009 103529
rect 120743 103615 121129 103634
rect 120743 103592 120809 103615
rect 120895 103592 120977 103615
rect 121063 103592 121129 103615
rect 120743 103552 120752 103592
rect 120792 103552 120809 103592
rect 120895 103552 120916 103592
rect 120956 103552 120977 103592
rect 121063 103552 121080 103592
rect 121120 103552 121129 103592
rect 120743 103529 120809 103552
rect 120895 103529 120977 103552
rect 121063 103529 121129 103552
rect 120743 103510 121129 103529
rect 135863 103615 136249 103634
rect 135863 103592 135929 103615
rect 136015 103592 136097 103615
rect 136183 103592 136249 103615
rect 135863 103552 135872 103592
rect 135912 103552 135929 103592
rect 136015 103552 136036 103592
rect 136076 103552 136097 103592
rect 136183 103552 136200 103592
rect 136240 103552 136249 103592
rect 135863 103529 135929 103552
rect 136015 103529 136097 103552
rect 136183 103529 136249 103552
rect 135863 103510 136249 103529
rect 150983 103615 151369 103634
rect 150983 103592 151049 103615
rect 151135 103592 151217 103615
rect 151303 103592 151369 103615
rect 150983 103552 150992 103592
rect 151032 103552 151049 103592
rect 151135 103552 151156 103592
rect 151196 103552 151217 103592
rect 151303 103552 151320 103592
rect 151360 103552 151369 103592
rect 150983 103529 151049 103552
rect 151135 103529 151217 103552
rect 151303 103529 151369 103552
rect 150983 103510 151369 103529
rect 74143 102859 74529 102878
rect 74143 102836 74209 102859
rect 74295 102836 74377 102859
rect 74463 102836 74529 102859
rect 74143 102796 74152 102836
rect 74192 102796 74209 102836
rect 74295 102796 74316 102836
rect 74356 102796 74377 102836
rect 74463 102796 74480 102836
rect 74520 102796 74529 102836
rect 74143 102773 74209 102796
rect 74295 102773 74377 102796
rect 74463 102773 74529 102796
rect 74143 102754 74529 102773
rect 89263 102859 89649 102878
rect 89263 102836 89329 102859
rect 89415 102836 89497 102859
rect 89583 102836 89649 102859
rect 89263 102796 89272 102836
rect 89312 102796 89329 102836
rect 89415 102796 89436 102836
rect 89476 102796 89497 102836
rect 89583 102796 89600 102836
rect 89640 102796 89649 102836
rect 89263 102773 89329 102796
rect 89415 102773 89497 102796
rect 89583 102773 89649 102796
rect 89263 102754 89649 102773
rect 104383 102859 104769 102878
rect 104383 102836 104449 102859
rect 104535 102836 104617 102859
rect 104703 102836 104769 102859
rect 104383 102796 104392 102836
rect 104432 102796 104449 102836
rect 104535 102796 104556 102836
rect 104596 102796 104617 102836
rect 104703 102796 104720 102836
rect 104760 102796 104769 102836
rect 104383 102773 104449 102796
rect 104535 102773 104617 102796
rect 104703 102773 104769 102796
rect 104383 102754 104769 102773
rect 119503 102859 119889 102878
rect 119503 102836 119569 102859
rect 119655 102836 119737 102859
rect 119823 102836 119889 102859
rect 119503 102796 119512 102836
rect 119552 102796 119569 102836
rect 119655 102796 119676 102836
rect 119716 102796 119737 102836
rect 119823 102796 119840 102836
rect 119880 102796 119889 102836
rect 119503 102773 119569 102796
rect 119655 102773 119737 102796
rect 119823 102773 119889 102796
rect 119503 102754 119889 102773
rect 134623 102859 135009 102878
rect 134623 102836 134689 102859
rect 134775 102836 134857 102859
rect 134943 102836 135009 102859
rect 134623 102796 134632 102836
rect 134672 102796 134689 102836
rect 134775 102796 134796 102836
rect 134836 102796 134857 102836
rect 134943 102796 134960 102836
rect 135000 102796 135009 102836
rect 134623 102773 134689 102796
rect 134775 102773 134857 102796
rect 134943 102773 135009 102796
rect 134623 102754 135009 102773
rect 149743 102859 150129 102878
rect 149743 102836 149809 102859
rect 149895 102836 149977 102859
rect 150063 102836 150129 102859
rect 149743 102796 149752 102836
rect 149792 102796 149809 102836
rect 149895 102796 149916 102836
rect 149956 102796 149977 102836
rect 150063 102796 150080 102836
rect 150120 102796 150129 102836
rect 149743 102773 149809 102796
rect 149895 102773 149977 102796
rect 150063 102773 150129 102796
rect 149743 102754 150129 102773
rect 75383 102103 75769 102122
rect 75383 102080 75449 102103
rect 75535 102080 75617 102103
rect 75703 102080 75769 102103
rect 75383 102040 75392 102080
rect 75432 102040 75449 102080
rect 75535 102040 75556 102080
rect 75596 102040 75617 102080
rect 75703 102040 75720 102080
rect 75760 102040 75769 102080
rect 75383 102017 75449 102040
rect 75535 102017 75617 102040
rect 75703 102017 75769 102040
rect 75383 101998 75769 102017
rect 90503 102103 90889 102122
rect 90503 102080 90569 102103
rect 90655 102080 90737 102103
rect 90823 102080 90889 102103
rect 90503 102040 90512 102080
rect 90552 102040 90569 102080
rect 90655 102040 90676 102080
rect 90716 102040 90737 102080
rect 90823 102040 90840 102080
rect 90880 102040 90889 102080
rect 90503 102017 90569 102040
rect 90655 102017 90737 102040
rect 90823 102017 90889 102040
rect 90503 101998 90889 102017
rect 105623 102103 106009 102122
rect 105623 102080 105689 102103
rect 105775 102080 105857 102103
rect 105943 102080 106009 102103
rect 105623 102040 105632 102080
rect 105672 102040 105689 102080
rect 105775 102040 105796 102080
rect 105836 102040 105857 102080
rect 105943 102040 105960 102080
rect 106000 102040 106009 102080
rect 105623 102017 105689 102040
rect 105775 102017 105857 102040
rect 105943 102017 106009 102040
rect 105623 101998 106009 102017
rect 120743 102103 121129 102122
rect 120743 102080 120809 102103
rect 120895 102080 120977 102103
rect 121063 102080 121129 102103
rect 120743 102040 120752 102080
rect 120792 102040 120809 102080
rect 120895 102040 120916 102080
rect 120956 102040 120977 102080
rect 121063 102040 121080 102080
rect 121120 102040 121129 102080
rect 120743 102017 120809 102040
rect 120895 102017 120977 102040
rect 121063 102017 121129 102040
rect 120743 101998 121129 102017
rect 135863 102103 136249 102122
rect 135863 102080 135929 102103
rect 136015 102080 136097 102103
rect 136183 102080 136249 102103
rect 135863 102040 135872 102080
rect 135912 102040 135929 102080
rect 136015 102040 136036 102080
rect 136076 102040 136097 102080
rect 136183 102040 136200 102080
rect 136240 102040 136249 102080
rect 135863 102017 135929 102040
rect 136015 102017 136097 102040
rect 136183 102017 136249 102040
rect 135863 101998 136249 102017
rect 150983 102103 151369 102122
rect 150983 102080 151049 102103
rect 151135 102080 151217 102103
rect 151303 102080 151369 102103
rect 150983 102040 150992 102080
rect 151032 102040 151049 102080
rect 151135 102040 151156 102080
rect 151196 102040 151217 102080
rect 151303 102040 151320 102080
rect 151360 102040 151369 102080
rect 150983 102017 151049 102040
rect 151135 102017 151217 102040
rect 151303 102017 151369 102040
rect 150983 101998 151369 102017
rect 74143 101347 74529 101366
rect 74143 101324 74209 101347
rect 74295 101324 74377 101347
rect 74463 101324 74529 101347
rect 74143 101284 74152 101324
rect 74192 101284 74209 101324
rect 74295 101284 74316 101324
rect 74356 101284 74377 101324
rect 74463 101284 74480 101324
rect 74520 101284 74529 101324
rect 74143 101261 74209 101284
rect 74295 101261 74377 101284
rect 74463 101261 74529 101284
rect 74143 101242 74529 101261
rect 89263 101347 89649 101366
rect 89263 101324 89329 101347
rect 89415 101324 89497 101347
rect 89583 101324 89649 101347
rect 89263 101284 89272 101324
rect 89312 101284 89329 101324
rect 89415 101284 89436 101324
rect 89476 101284 89497 101324
rect 89583 101284 89600 101324
rect 89640 101284 89649 101324
rect 89263 101261 89329 101284
rect 89415 101261 89497 101284
rect 89583 101261 89649 101284
rect 89263 101242 89649 101261
rect 104383 101347 104769 101366
rect 104383 101324 104449 101347
rect 104535 101324 104617 101347
rect 104703 101324 104769 101347
rect 104383 101284 104392 101324
rect 104432 101284 104449 101324
rect 104535 101284 104556 101324
rect 104596 101284 104617 101324
rect 104703 101284 104720 101324
rect 104760 101284 104769 101324
rect 104383 101261 104449 101284
rect 104535 101261 104617 101284
rect 104703 101261 104769 101284
rect 104383 101242 104769 101261
rect 119503 101347 119889 101366
rect 119503 101324 119569 101347
rect 119655 101324 119737 101347
rect 119823 101324 119889 101347
rect 119503 101284 119512 101324
rect 119552 101284 119569 101324
rect 119655 101284 119676 101324
rect 119716 101284 119737 101324
rect 119823 101284 119840 101324
rect 119880 101284 119889 101324
rect 119503 101261 119569 101284
rect 119655 101261 119737 101284
rect 119823 101261 119889 101284
rect 119503 101242 119889 101261
rect 134623 101347 135009 101366
rect 134623 101324 134689 101347
rect 134775 101324 134857 101347
rect 134943 101324 135009 101347
rect 134623 101284 134632 101324
rect 134672 101284 134689 101324
rect 134775 101284 134796 101324
rect 134836 101284 134857 101324
rect 134943 101284 134960 101324
rect 135000 101284 135009 101324
rect 134623 101261 134689 101284
rect 134775 101261 134857 101284
rect 134943 101261 135009 101284
rect 134623 101242 135009 101261
rect 149743 101347 150129 101366
rect 149743 101324 149809 101347
rect 149895 101324 149977 101347
rect 150063 101324 150129 101347
rect 149743 101284 149752 101324
rect 149792 101284 149809 101324
rect 149895 101284 149916 101324
rect 149956 101284 149977 101324
rect 150063 101284 150080 101324
rect 150120 101284 150129 101324
rect 149743 101261 149809 101284
rect 149895 101261 149977 101284
rect 150063 101261 150129 101284
rect 149743 101242 150129 101261
rect 75383 100591 75769 100610
rect 75383 100568 75449 100591
rect 75535 100568 75617 100591
rect 75703 100568 75769 100591
rect 75383 100528 75392 100568
rect 75432 100528 75449 100568
rect 75535 100528 75556 100568
rect 75596 100528 75617 100568
rect 75703 100528 75720 100568
rect 75760 100528 75769 100568
rect 75383 100505 75449 100528
rect 75535 100505 75617 100528
rect 75703 100505 75769 100528
rect 75383 100486 75769 100505
rect 90503 100591 90889 100610
rect 90503 100568 90569 100591
rect 90655 100568 90737 100591
rect 90823 100568 90889 100591
rect 90503 100528 90512 100568
rect 90552 100528 90569 100568
rect 90655 100528 90676 100568
rect 90716 100528 90737 100568
rect 90823 100528 90840 100568
rect 90880 100528 90889 100568
rect 90503 100505 90569 100528
rect 90655 100505 90737 100528
rect 90823 100505 90889 100528
rect 90503 100486 90889 100505
rect 105623 100591 106009 100610
rect 105623 100568 105689 100591
rect 105775 100568 105857 100591
rect 105943 100568 106009 100591
rect 105623 100528 105632 100568
rect 105672 100528 105689 100568
rect 105775 100528 105796 100568
rect 105836 100528 105857 100568
rect 105943 100528 105960 100568
rect 106000 100528 106009 100568
rect 105623 100505 105689 100528
rect 105775 100505 105857 100528
rect 105943 100505 106009 100528
rect 105623 100486 106009 100505
rect 120743 100591 121129 100610
rect 120743 100568 120809 100591
rect 120895 100568 120977 100591
rect 121063 100568 121129 100591
rect 120743 100528 120752 100568
rect 120792 100528 120809 100568
rect 120895 100528 120916 100568
rect 120956 100528 120977 100568
rect 121063 100528 121080 100568
rect 121120 100528 121129 100568
rect 120743 100505 120809 100528
rect 120895 100505 120977 100528
rect 121063 100505 121129 100528
rect 120743 100486 121129 100505
rect 135863 100591 136249 100610
rect 135863 100568 135929 100591
rect 136015 100568 136097 100591
rect 136183 100568 136249 100591
rect 135863 100528 135872 100568
rect 135912 100528 135929 100568
rect 136015 100528 136036 100568
rect 136076 100528 136097 100568
rect 136183 100528 136200 100568
rect 136240 100528 136249 100568
rect 135863 100505 135929 100528
rect 136015 100505 136097 100528
rect 136183 100505 136249 100528
rect 135863 100486 136249 100505
rect 150983 100591 151369 100610
rect 150983 100568 151049 100591
rect 151135 100568 151217 100591
rect 151303 100568 151369 100591
rect 150983 100528 150992 100568
rect 151032 100528 151049 100568
rect 151135 100528 151156 100568
rect 151196 100528 151217 100568
rect 151303 100528 151320 100568
rect 151360 100528 151369 100568
rect 150983 100505 151049 100528
rect 151135 100505 151217 100528
rect 151303 100505 151369 100528
rect 150983 100486 151369 100505
rect 74143 99835 74529 99854
rect 74143 99812 74209 99835
rect 74295 99812 74377 99835
rect 74463 99812 74529 99835
rect 74143 99772 74152 99812
rect 74192 99772 74209 99812
rect 74295 99772 74316 99812
rect 74356 99772 74377 99812
rect 74463 99772 74480 99812
rect 74520 99772 74529 99812
rect 74143 99749 74209 99772
rect 74295 99749 74377 99772
rect 74463 99749 74529 99772
rect 74143 99730 74529 99749
rect 89263 99835 89649 99854
rect 89263 99812 89329 99835
rect 89415 99812 89497 99835
rect 89583 99812 89649 99835
rect 89263 99772 89272 99812
rect 89312 99772 89329 99812
rect 89415 99772 89436 99812
rect 89476 99772 89497 99812
rect 89583 99772 89600 99812
rect 89640 99772 89649 99812
rect 89263 99749 89329 99772
rect 89415 99749 89497 99772
rect 89583 99749 89649 99772
rect 89263 99730 89649 99749
rect 104383 99835 104769 99854
rect 104383 99812 104449 99835
rect 104535 99812 104617 99835
rect 104703 99812 104769 99835
rect 104383 99772 104392 99812
rect 104432 99772 104449 99812
rect 104535 99772 104556 99812
rect 104596 99772 104617 99812
rect 104703 99772 104720 99812
rect 104760 99772 104769 99812
rect 104383 99749 104449 99772
rect 104535 99749 104617 99772
rect 104703 99749 104769 99772
rect 104383 99730 104769 99749
rect 119503 99835 119889 99854
rect 119503 99812 119569 99835
rect 119655 99812 119737 99835
rect 119823 99812 119889 99835
rect 119503 99772 119512 99812
rect 119552 99772 119569 99812
rect 119655 99772 119676 99812
rect 119716 99772 119737 99812
rect 119823 99772 119840 99812
rect 119880 99772 119889 99812
rect 119503 99749 119569 99772
rect 119655 99749 119737 99772
rect 119823 99749 119889 99772
rect 119503 99730 119889 99749
rect 134623 99835 135009 99854
rect 134623 99812 134689 99835
rect 134775 99812 134857 99835
rect 134943 99812 135009 99835
rect 134623 99772 134632 99812
rect 134672 99772 134689 99812
rect 134775 99772 134796 99812
rect 134836 99772 134857 99812
rect 134943 99772 134960 99812
rect 135000 99772 135009 99812
rect 134623 99749 134689 99772
rect 134775 99749 134857 99772
rect 134943 99749 135009 99772
rect 134623 99730 135009 99749
rect 149743 99835 150129 99854
rect 149743 99812 149809 99835
rect 149895 99812 149977 99835
rect 150063 99812 150129 99835
rect 149743 99772 149752 99812
rect 149792 99772 149809 99812
rect 149895 99772 149916 99812
rect 149956 99772 149977 99812
rect 150063 99772 150080 99812
rect 150120 99772 150129 99812
rect 149743 99749 149809 99772
rect 149895 99749 149977 99772
rect 150063 99749 150129 99772
rect 149743 99730 150129 99749
rect 75383 99079 75769 99098
rect 75383 99056 75449 99079
rect 75535 99056 75617 99079
rect 75703 99056 75769 99079
rect 75383 99016 75392 99056
rect 75432 99016 75449 99056
rect 75535 99016 75556 99056
rect 75596 99016 75617 99056
rect 75703 99016 75720 99056
rect 75760 99016 75769 99056
rect 75383 98993 75449 99016
rect 75535 98993 75617 99016
rect 75703 98993 75769 99016
rect 75383 98974 75769 98993
rect 90503 99079 90889 99098
rect 90503 99056 90569 99079
rect 90655 99056 90737 99079
rect 90823 99056 90889 99079
rect 90503 99016 90512 99056
rect 90552 99016 90569 99056
rect 90655 99016 90676 99056
rect 90716 99016 90737 99056
rect 90823 99016 90840 99056
rect 90880 99016 90889 99056
rect 90503 98993 90569 99016
rect 90655 98993 90737 99016
rect 90823 98993 90889 99016
rect 90503 98974 90889 98993
rect 105623 99079 106009 99098
rect 105623 99056 105689 99079
rect 105775 99056 105857 99079
rect 105943 99056 106009 99079
rect 105623 99016 105632 99056
rect 105672 99016 105689 99056
rect 105775 99016 105796 99056
rect 105836 99016 105857 99056
rect 105943 99016 105960 99056
rect 106000 99016 106009 99056
rect 105623 98993 105689 99016
rect 105775 98993 105857 99016
rect 105943 98993 106009 99016
rect 105623 98974 106009 98993
rect 120743 99079 121129 99098
rect 120743 99056 120809 99079
rect 120895 99056 120977 99079
rect 121063 99056 121129 99079
rect 120743 99016 120752 99056
rect 120792 99016 120809 99056
rect 120895 99016 120916 99056
rect 120956 99016 120977 99056
rect 121063 99016 121080 99056
rect 121120 99016 121129 99056
rect 120743 98993 120809 99016
rect 120895 98993 120977 99016
rect 121063 98993 121129 99016
rect 120743 98974 121129 98993
rect 135863 99079 136249 99098
rect 135863 99056 135929 99079
rect 136015 99056 136097 99079
rect 136183 99056 136249 99079
rect 135863 99016 135872 99056
rect 135912 99016 135929 99056
rect 136015 99016 136036 99056
rect 136076 99016 136097 99056
rect 136183 99016 136200 99056
rect 136240 99016 136249 99056
rect 135863 98993 135929 99016
rect 136015 98993 136097 99016
rect 136183 98993 136249 99016
rect 135863 98974 136249 98993
rect 150983 99079 151369 99098
rect 150983 99056 151049 99079
rect 151135 99056 151217 99079
rect 151303 99056 151369 99079
rect 150983 99016 150992 99056
rect 151032 99016 151049 99056
rect 151135 99016 151156 99056
rect 151196 99016 151217 99056
rect 151303 99016 151320 99056
rect 151360 99016 151369 99056
rect 150983 98993 151049 99016
rect 151135 98993 151217 99016
rect 151303 98993 151369 99016
rect 150983 98974 151369 98993
rect 74143 98323 74529 98342
rect 74143 98300 74209 98323
rect 74295 98300 74377 98323
rect 74463 98300 74529 98323
rect 74143 98260 74152 98300
rect 74192 98260 74209 98300
rect 74295 98260 74316 98300
rect 74356 98260 74377 98300
rect 74463 98260 74480 98300
rect 74520 98260 74529 98300
rect 74143 98237 74209 98260
rect 74295 98237 74377 98260
rect 74463 98237 74529 98260
rect 74143 98218 74529 98237
rect 89263 98323 89649 98342
rect 89263 98300 89329 98323
rect 89415 98300 89497 98323
rect 89583 98300 89649 98323
rect 89263 98260 89272 98300
rect 89312 98260 89329 98300
rect 89415 98260 89436 98300
rect 89476 98260 89497 98300
rect 89583 98260 89600 98300
rect 89640 98260 89649 98300
rect 89263 98237 89329 98260
rect 89415 98237 89497 98260
rect 89583 98237 89649 98260
rect 89263 98218 89649 98237
rect 104383 98323 104769 98342
rect 104383 98300 104449 98323
rect 104535 98300 104617 98323
rect 104703 98300 104769 98323
rect 104383 98260 104392 98300
rect 104432 98260 104449 98300
rect 104535 98260 104556 98300
rect 104596 98260 104617 98300
rect 104703 98260 104720 98300
rect 104760 98260 104769 98300
rect 104383 98237 104449 98260
rect 104535 98237 104617 98260
rect 104703 98237 104769 98260
rect 104383 98218 104769 98237
rect 119503 98323 119889 98342
rect 119503 98300 119569 98323
rect 119655 98300 119737 98323
rect 119823 98300 119889 98323
rect 119503 98260 119512 98300
rect 119552 98260 119569 98300
rect 119655 98260 119676 98300
rect 119716 98260 119737 98300
rect 119823 98260 119840 98300
rect 119880 98260 119889 98300
rect 119503 98237 119569 98260
rect 119655 98237 119737 98260
rect 119823 98237 119889 98260
rect 119503 98218 119889 98237
rect 134623 98323 135009 98342
rect 134623 98300 134689 98323
rect 134775 98300 134857 98323
rect 134943 98300 135009 98323
rect 134623 98260 134632 98300
rect 134672 98260 134689 98300
rect 134775 98260 134796 98300
rect 134836 98260 134857 98300
rect 134943 98260 134960 98300
rect 135000 98260 135009 98300
rect 134623 98237 134689 98260
rect 134775 98237 134857 98260
rect 134943 98237 135009 98260
rect 134623 98218 135009 98237
rect 149743 98323 150129 98342
rect 149743 98300 149809 98323
rect 149895 98300 149977 98323
rect 150063 98300 150129 98323
rect 149743 98260 149752 98300
rect 149792 98260 149809 98300
rect 149895 98260 149916 98300
rect 149956 98260 149977 98300
rect 150063 98260 150080 98300
rect 150120 98260 150129 98300
rect 149743 98237 149809 98260
rect 149895 98237 149977 98260
rect 150063 98237 150129 98260
rect 149743 98218 150129 98237
rect 75383 97567 75769 97586
rect 75383 97544 75449 97567
rect 75535 97544 75617 97567
rect 75703 97544 75769 97567
rect 75383 97504 75392 97544
rect 75432 97504 75449 97544
rect 75535 97504 75556 97544
rect 75596 97504 75617 97544
rect 75703 97504 75720 97544
rect 75760 97504 75769 97544
rect 75383 97481 75449 97504
rect 75535 97481 75617 97504
rect 75703 97481 75769 97504
rect 75383 97462 75769 97481
rect 90503 97567 90889 97586
rect 90503 97544 90569 97567
rect 90655 97544 90737 97567
rect 90823 97544 90889 97567
rect 90503 97504 90512 97544
rect 90552 97504 90569 97544
rect 90655 97504 90676 97544
rect 90716 97504 90737 97544
rect 90823 97504 90840 97544
rect 90880 97504 90889 97544
rect 90503 97481 90569 97504
rect 90655 97481 90737 97504
rect 90823 97481 90889 97504
rect 90503 97462 90889 97481
rect 105623 97567 106009 97586
rect 105623 97544 105689 97567
rect 105775 97544 105857 97567
rect 105943 97544 106009 97567
rect 105623 97504 105632 97544
rect 105672 97504 105689 97544
rect 105775 97504 105796 97544
rect 105836 97504 105857 97544
rect 105943 97504 105960 97544
rect 106000 97504 106009 97544
rect 105623 97481 105689 97504
rect 105775 97481 105857 97504
rect 105943 97481 106009 97504
rect 105623 97462 106009 97481
rect 120743 97567 121129 97586
rect 120743 97544 120809 97567
rect 120895 97544 120977 97567
rect 121063 97544 121129 97567
rect 120743 97504 120752 97544
rect 120792 97504 120809 97544
rect 120895 97504 120916 97544
rect 120956 97504 120977 97544
rect 121063 97504 121080 97544
rect 121120 97504 121129 97544
rect 120743 97481 120809 97504
rect 120895 97481 120977 97504
rect 121063 97481 121129 97504
rect 120743 97462 121129 97481
rect 135863 97567 136249 97586
rect 135863 97544 135929 97567
rect 136015 97544 136097 97567
rect 136183 97544 136249 97567
rect 135863 97504 135872 97544
rect 135912 97504 135929 97544
rect 136015 97504 136036 97544
rect 136076 97504 136097 97544
rect 136183 97504 136200 97544
rect 136240 97504 136249 97544
rect 135863 97481 135929 97504
rect 136015 97481 136097 97504
rect 136183 97481 136249 97504
rect 135863 97462 136249 97481
rect 150983 97567 151369 97586
rect 150983 97544 151049 97567
rect 151135 97544 151217 97567
rect 151303 97544 151369 97567
rect 150983 97504 150992 97544
rect 151032 97504 151049 97544
rect 151135 97504 151156 97544
rect 151196 97504 151217 97544
rect 151303 97504 151320 97544
rect 151360 97504 151369 97544
rect 150983 97481 151049 97504
rect 151135 97481 151217 97504
rect 151303 97481 151369 97504
rect 150983 97462 151369 97481
rect 74143 96811 74529 96830
rect 74143 96788 74209 96811
rect 74295 96788 74377 96811
rect 74463 96788 74529 96811
rect 74143 96748 74152 96788
rect 74192 96748 74209 96788
rect 74295 96748 74316 96788
rect 74356 96748 74377 96788
rect 74463 96748 74480 96788
rect 74520 96748 74529 96788
rect 74143 96725 74209 96748
rect 74295 96725 74377 96748
rect 74463 96725 74529 96748
rect 74143 96706 74529 96725
rect 89263 96811 89649 96830
rect 89263 96788 89329 96811
rect 89415 96788 89497 96811
rect 89583 96788 89649 96811
rect 89263 96748 89272 96788
rect 89312 96748 89329 96788
rect 89415 96748 89436 96788
rect 89476 96748 89497 96788
rect 89583 96748 89600 96788
rect 89640 96748 89649 96788
rect 89263 96725 89329 96748
rect 89415 96725 89497 96748
rect 89583 96725 89649 96748
rect 89263 96706 89649 96725
rect 104383 96811 104769 96830
rect 104383 96788 104449 96811
rect 104535 96788 104617 96811
rect 104703 96788 104769 96811
rect 104383 96748 104392 96788
rect 104432 96748 104449 96788
rect 104535 96748 104556 96788
rect 104596 96748 104617 96788
rect 104703 96748 104720 96788
rect 104760 96748 104769 96788
rect 104383 96725 104449 96748
rect 104535 96725 104617 96748
rect 104703 96725 104769 96748
rect 104383 96706 104769 96725
rect 119503 96811 119889 96830
rect 119503 96788 119569 96811
rect 119655 96788 119737 96811
rect 119823 96788 119889 96811
rect 119503 96748 119512 96788
rect 119552 96748 119569 96788
rect 119655 96748 119676 96788
rect 119716 96748 119737 96788
rect 119823 96748 119840 96788
rect 119880 96748 119889 96788
rect 119503 96725 119569 96748
rect 119655 96725 119737 96748
rect 119823 96725 119889 96748
rect 119503 96706 119889 96725
rect 134623 96811 135009 96830
rect 134623 96788 134689 96811
rect 134775 96788 134857 96811
rect 134943 96788 135009 96811
rect 134623 96748 134632 96788
rect 134672 96748 134689 96788
rect 134775 96748 134796 96788
rect 134836 96748 134857 96788
rect 134943 96748 134960 96788
rect 135000 96748 135009 96788
rect 134623 96725 134689 96748
rect 134775 96725 134857 96748
rect 134943 96725 135009 96748
rect 134623 96706 135009 96725
rect 149743 96811 150129 96830
rect 149743 96788 149809 96811
rect 149895 96788 149977 96811
rect 150063 96788 150129 96811
rect 149743 96748 149752 96788
rect 149792 96748 149809 96788
rect 149895 96748 149916 96788
rect 149956 96748 149977 96788
rect 150063 96748 150080 96788
rect 150120 96748 150129 96788
rect 149743 96725 149809 96748
rect 149895 96725 149977 96748
rect 150063 96725 150129 96748
rect 149743 96706 150129 96725
rect 75383 96055 75769 96074
rect 75383 96032 75449 96055
rect 75535 96032 75617 96055
rect 75703 96032 75769 96055
rect 75383 95992 75392 96032
rect 75432 95992 75449 96032
rect 75535 95992 75556 96032
rect 75596 95992 75617 96032
rect 75703 95992 75720 96032
rect 75760 95992 75769 96032
rect 75383 95969 75449 95992
rect 75535 95969 75617 95992
rect 75703 95969 75769 95992
rect 75383 95950 75769 95969
rect 90503 96055 90889 96074
rect 90503 96032 90569 96055
rect 90655 96032 90737 96055
rect 90823 96032 90889 96055
rect 90503 95992 90512 96032
rect 90552 95992 90569 96032
rect 90655 95992 90676 96032
rect 90716 95992 90737 96032
rect 90823 95992 90840 96032
rect 90880 95992 90889 96032
rect 90503 95969 90569 95992
rect 90655 95969 90737 95992
rect 90823 95969 90889 95992
rect 90503 95950 90889 95969
rect 105623 96055 106009 96074
rect 105623 96032 105689 96055
rect 105775 96032 105857 96055
rect 105943 96032 106009 96055
rect 105623 95992 105632 96032
rect 105672 95992 105689 96032
rect 105775 95992 105796 96032
rect 105836 95992 105857 96032
rect 105943 95992 105960 96032
rect 106000 95992 106009 96032
rect 105623 95969 105689 95992
rect 105775 95969 105857 95992
rect 105943 95969 106009 95992
rect 105623 95950 106009 95969
rect 120743 96055 121129 96074
rect 120743 96032 120809 96055
rect 120895 96032 120977 96055
rect 121063 96032 121129 96055
rect 120743 95992 120752 96032
rect 120792 95992 120809 96032
rect 120895 95992 120916 96032
rect 120956 95992 120977 96032
rect 121063 95992 121080 96032
rect 121120 95992 121129 96032
rect 120743 95969 120809 95992
rect 120895 95969 120977 95992
rect 121063 95969 121129 95992
rect 120743 95950 121129 95969
rect 135863 96055 136249 96074
rect 135863 96032 135929 96055
rect 136015 96032 136097 96055
rect 136183 96032 136249 96055
rect 135863 95992 135872 96032
rect 135912 95992 135929 96032
rect 136015 95992 136036 96032
rect 136076 95992 136097 96032
rect 136183 95992 136200 96032
rect 136240 95992 136249 96032
rect 135863 95969 135929 95992
rect 136015 95969 136097 95992
rect 136183 95969 136249 95992
rect 135863 95950 136249 95969
rect 150983 96055 151369 96074
rect 150983 96032 151049 96055
rect 151135 96032 151217 96055
rect 151303 96032 151369 96055
rect 150983 95992 150992 96032
rect 151032 95992 151049 96032
rect 151135 95992 151156 96032
rect 151196 95992 151217 96032
rect 151303 95992 151320 96032
rect 151360 95992 151369 96032
rect 150983 95969 151049 95992
rect 151135 95969 151217 95992
rect 151303 95969 151369 95992
rect 150983 95950 151369 95969
rect 74143 95299 74529 95318
rect 74143 95276 74209 95299
rect 74295 95276 74377 95299
rect 74463 95276 74529 95299
rect 74143 95236 74152 95276
rect 74192 95236 74209 95276
rect 74295 95236 74316 95276
rect 74356 95236 74377 95276
rect 74463 95236 74480 95276
rect 74520 95236 74529 95276
rect 74143 95213 74209 95236
rect 74295 95213 74377 95236
rect 74463 95213 74529 95236
rect 74143 95194 74529 95213
rect 89263 95299 89649 95318
rect 89263 95276 89329 95299
rect 89415 95276 89497 95299
rect 89583 95276 89649 95299
rect 89263 95236 89272 95276
rect 89312 95236 89329 95276
rect 89415 95236 89436 95276
rect 89476 95236 89497 95276
rect 89583 95236 89600 95276
rect 89640 95236 89649 95276
rect 89263 95213 89329 95236
rect 89415 95213 89497 95236
rect 89583 95213 89649 95236
rect 89263 95194 89649 95213
rect 104383 95299 104769 95318
rect 104383 95276 104449 95299
rect 104535 95276 104617 95299
rect 104703 95276 104769 95299
rect 104383 95236 104392 95276
rect 104432 95236 104449 95276
rect 104535 95236 104556 95276
rect 104596 95236 104617 95276
rect 104703 95236 104720 95276
rect 104760 95236 104769 95276
rect 104383 95213 104449 95236
rect 104535 95213 104617 95236
rect 104703 95213 104769 95236
rect 104383 95194 104769 95213
rect 119503 95299 119889 95318
rect 119503 95276 119569 95299
rect 119655 95276 119737 95299
rect 119823 95276 119889 95299
rect 119503 95236 119512 95276
rect 119552 95236 119569 95276
rect 119655 95236 119676 95276
rect 119716 95236 119737 95276
rect 119823 95236 119840 95276
rect 119880 95236 119889 95276
rect 119503 95213 119569 95236
rect 119655 95213 119737 95236
rect 119823 95213 119889 95236
rect 119503 95194 119889 95213
rect 134623 95299 135009 95318
rect 134623 95276 134689 95299
rect 134775 95276 134857 95299
rect 134943 95276 135009 95299
rect 134623 95236 134632 95276
rect 134672 95236 134689 95276
rect 134775 95236 134796 95276
rect 134836 95236 134857 95276
rect 134943 95236 134960 95276
rect 135000 95236 135009 95276
rect 134623 95213 134689 95236
rect 134775 95213 134857 95236
rect 134943 95213 135009 95236
rect 134623 95194 135009 95213
rect 149743 95299 150129 95318
rect 149743 95276 149809 95299
rect 149895 95276 149977 95299
rect 150063 95276 150129 95299
rect 149743 95236 149752 95276
rect 149792 95236 149809 95276
rect 149895 95236 149916 95276
rect 149956 95236 149977 95276
rect 150063 95236 150080 95276
rect 150120 95236 150129 95276
rect 149743 95213 149809 95236
rect 149895 95213 149977 95236
rect 150063 95213 150129 95236
rect 149743 95194 150129 95213
rect 75383 94543 75769 94562
rect 75383 94520 75449 94543
rect 75535 94520 75617 94543
rect 75703 94520 75769 94543
rect 75383 94480 75392 94520
rect 75432 94480 75449 94520
rect 75535 94480 75556 94520
rect 75596 94480 75617 94520
rect 75703 94480 75720 94520
rect 75760 94480 75769 94520
rect 75383 94457 75449 94480
rect 75535 94457 75617 94480
rect 75703 94457 75769 94480
rect 75383 94438 75769 94457
rect 90503 94543 90889 94562
rect 90503 94520 90569 94543
rect 90655 94520 90737 94543
rect 90823 94520 90889 94543
rect 90503 94480 90512 94520
rect 90552 94480 90569 94520
rect 90655 94480 90676 94520
rect 90716 94480 90737 94520
rect 90823 94480 90840 94520
rect 90880 94480 90889 94520
rect 90503 94457 90569 94480
rect 90655 94457 90737 94480
rect 90823 94457 90889 94480
rect 90503 94438 90889 94457
rect 105623 94543 106009 94562
rect 105623 94520 105689 94543
rect 105775 94520 105857 94543
rect 105943 94520 106009 94543
rect 105623 94480 105632 94520
rect 105672 94480 105689 94520
rect 105775 94480 105796 94520
rect 105836 94480 105857 94520
rect 105943 94480 105960 94520
rect 106000 94480 106009 94520
rect 105623 94457 105689 94480
rect 105775 94457 105857 94480
rect 105943 94457 106009 94480
rect 105623 94438 106009 94457
rect 120743 94543 121129 94562
rect 120743 94520 120809 94543
rect 120895 94520 120977 94543
rect 121063 94520 121129 94543
rect 120743 94480 120752 94520
rect 120792 94480 120809 94520
rect 120895 94480 120916 94520
rect 120956 94480 120977 94520
rect 121063 94480 121080 94520
rect 121120 94480 121129 94520
rect 120743 94457 120809 94480
rect 120895 94457 120977 94480
rect 121063 94457 121129 94480
rect 120743 94438 121129 94457
rect 135863 94543 136249 94562
rect 135863 94520 135929 94543
rect 136015 94520 136097 94543
rect 136183 94520 136249 94543
rect 135863 94480 135872 94520
rect 135912 94480 135929 94520
rect 136015 94480 136036 94520
rect 136076 94480 136097 94520
rect 136183 94480 136200 94520
rect 136240 94480 136249 94520
rect 135863 94457 135929 94480
rect 136015 94457 136097 94480
rect 136183 94457 136249 94480
rect 135863 94438 136249 94457
rect 150983 94543 151369 94562
rect 150983 94520 151049 94543
rect 151135 94520 151217 94543
rect 151303 94520 151369 94543
rect 150983 94480 150992 94520
rect 151032 94480 151049 94520
rect 151135 94480 151156 94520
rect 151196 94480 151217 94520
rect 151303 94480 151320 94520
rect 151360 94480 151369 94520
rect 150983 94457 151049 94480
rect 151135 94457 151217 94480
rect 151303 94457 151369 94480
rect 150983 94438 151369 94457
rect 74143 93787 74529 93806
rect 74143 93764 74209 93787
rect 74295 93764 74377 93787
rect 74463 93764 74529 93787
rect 74143 93724 74152 93764
rect 74192 93724 74209 93764
rect 74295 93724 74316 93764
rect 74356 93724 74377 93764
rect 74463 93724 74480 93764
rect 74520 93724 74529 93764
rect 74143 93701 74209 93724
rect 74295 93701 74377 93724
rect 74463 93701 74529 93724
rect 74143 93682 74529 93701
rect 89263 93787 89649 93806
rect 89263 93764 89329 93787
rect 89415 93764 89497 93787
rect 89583 93764 89649 93787
rect 89263 93724 89272 93764
rect 89312 93724 89329 93764
rect 89415 93724 89436 93764
rect 89476 93724 89497 93764
rect 89583 93724 89600 93764
rect 89640 93724 89649 93764
rect 89263 93701 89329 93724
rect 89415 93701 89497 93724
rect 89583 93701 89649 93724
rect 89263 93682 89649 93701
rect 104383 93787 104769 93806
rect 104383 93764 104449 93787
rect 104535 93764 104617 93787
rect 104703 93764 104769 93787
rect 104383 93724 104392 93764
rect 104432 93724 104449 93764
rect 104535 93724 104556 93764
rect 104596 93724 104617 93764
rect 104703 93724 104720 93764
rect 104760 93724 104769 93764
rect 104383 93701 104449 93724
rect 104535 93701 104617 93724
rect 104703 93701 104769 93724
rect 104383 93682 104769 93701
rect 119503 93787 119889 93806
rect 119503 93764 119569 93787
rect 119655 93764 119737 93787
rect 119823 93764 119889 93787
rect 119503 93724 119512 93764
rect 119552 93724 119569 93764
rect 119655 93724 119676 93764
rect 119716 93724 119737 93764
rect 119823 93724 119840 93764
rect 119880 93724 119889 93764
rect 119503 93701 119569 93724
rect 119655 93701 119737 93724
rect 119823 93701 119889 93724
rect 119503 93682 119889 93701
rect 134623 93787 135009 93806
rect 134623 93764 134689 93787
rect 134775 93764 134857 93787
rect 134943 93764 135009 93787
rect 134623 93724 134632 93764
rect 134672 93724 134689 93764
rect 134775 93724 134796 93764
rect 134836 93724 134857 93764
rect 134943 93724 134960 93764
rect 135000 93724 135009 93764
rect 134623 93701 134689 93724
rect 134775 93701 134857 93724
rect 134943 93701 135009 93724
rect 134623 93682 135009 93701
rect 149743 93787 150129 93806
rect 149743 93764 149809 93787
rect 149895 93764 149977 93787
rect 150063 93764 150129 93787
rect 149743 93724 149752 93764
rect 149792 93724 149809 93764
rect 149895 93724 149916 93764
rect 149956 93724 149977 93764
rect 150063 93724 150080 93764
rect 150120 93724 150129 93764
rect 149743 93701 149809 93724
rect 149895 93701 149977 93724
rect 150063 93701 150129 93724
rect 149743 93682 150129 93701
rect 75383 93031 75769 93050
rect 75383 93008 75449 93031
rect 75535 93008 75617 93031
rect 75703 93008 75769 93031
rect 75383 92968 75392 93008
rect 75432 92968 75449 93008
rect 75535 92968 75556 93008
rect 75596 92968 75617 93008
rect 75703 92968 75720 93008
rect 75760 92968 75769 93008
rect 75383 92945 75449 92968
rect 75535 92945 75617 92968
rect 75703 92945 75769 92968
rect 75383 92926 75769 92945
rect 90503 93031 90889 93050
rect 90503 93008 90569 93031
rect 90655 93008 90737 93031
rect 90823 93008 90889 93031
rect 90503 92968 90512 93008
rect 90552 92968 90569 93008
rect 90655 92968 90676 93008
rect 90716 92968 90737 93008
rect 90823 92968 90840 93008
rect 90880 92968 90889 93008
rect 90503 92945 90569 92968
rect 90655 92945 90737 92968
rect 90823 92945 90889 92968
rect 90503 92926 90889 92945
rect 105623 93031 106009 93050
rect 105623 93008 105689 93031
rect 105775 93008 105857 93031
rect 105943 93008 106009 93031
rect 105623 92968 105632 93008
rect 105672 92968 105689 93008
rect 105775 92968 105796 93008
rect 105836 92968 105857 93008
rect 105943 92968 105960 93008
rect 106000 92968 106009 93008
rect 105623 92945 105689 92968
rect 105775 92945 105857 92968
rect 105943 92945 106009 92968
rect 105623 92926 106009 92945
rect 120743 93031 121129 93050
rect 120743 93008 120809 93031
rect 120895 93008 120977 93031
rect 121063 93008 121129 93031
rect 120743 92968 120752 93008
rect 120792 92968 120809 93008
rect 120895 92968 120916 93008
rect 120956 92968 120977 93008
rect 121063 92968 121080 93008
rect 121120 92968 121129 93008
rect 120743 92945 120809 92968
rect 120895 92945 120977 92968
rect 121063 92945 121129 92968
rect 120743 92926 121129 92945
rect 135863 93031 136249 93050
rect 135863 93008 135929 93031
rect 136015 93008 136097 93031
rect 136183 93008 136249 93031
rect 135863 92968 135872 93008
rect 135912 92968 135929 93008
rect 136015 92968 136036 93008
rect 136076 92968 136097 93008
rect 136183 92968 136200 93008
rect 136240 92968 136249 93008
rect 135863 92945 135929 92968
rect 136015 92945 136097 92968
rect 136183 92945 136249 92968
rect 135863 92926 136249 92945
rect 150983 93031 151369 93050
rect 150983 93008 151049 93031
rect 151135 93008 151217 93031
rect 151303 93008 151369 93031
rect 150983 92968 150992 93008
rect 151032 92968 151049 93008
rect 151135 92968 151156 93008
rect 151196 92968 151217 93008
rect 151303 92968 151320 93008
rect 151360 92968 151369 93008
rect 150983 92945 151049 92968
rect 151135 92945 151217 92968
rect 151303 92945 151369 92968
rect 150983 92926 151369 92945
rect 74143 92275 74529 92294
rect 74143 92252 74209 92275
rect 74295 92252 74377 92275
rect 74463 92252 74529 92275
rect 74143 92212 74152 92252
rect 74192 92212 74209 92252
rect 74295 92212 74316 92252
rect 74356 92212 74377 92252
rect 74463 92212 74480 92252
rect 74520 92212 74529 92252
rect 74143 92189 74209 92212
rect 74295 92189 74377 92212
rect 74463 92189 74529 92212
rect 74143 92170 74529 92189
rect 89263 92275 89649 92294
rect 89263 92252 89329 92275
rect 89415 92252 89497 92275
rect 89583 92252 89649 92275
rect 89263 92212 89272 92252
rect 89312 92212 89329 92252
rect 89415 92212 89436 92252
rect 89476 92212 89497 92252
rect 89583 92212 89600 92252
rect 89640 92212 89649 92252
rect 89263 92189 89329 92212
rect 89415 92189 89497 92212
rect 89583 92189 89649 92212
rect 89263 92170 89649 92189
rect 104383 92275 104769 92294
rect 104383 92252 104449 92275
rect 104535 92252 104617 92275
rect 104703 92252 104769 92275
rect 104383 92212 104392 92252
rect 104432 92212 104449 92252
rect 104535 92212 104556 92252
rect 104596 92212 104617 92252
rect 104703 92212 104720 92252
rect 104760 92212 104769 92252
rect 104383 92189 104449 92212
rect 104535 92189 104617 92212
rect 104703 92189 104769 92212
rect 104383 92170 104769 92189
rect 119503 92275 119889 92294
rect 119503 92252 119569 92275
rect 119655 92252 119737 92275
rect 119823 92252 119889 92275
rect 119503 92212 119512 92252
rect 119552 92212 119569 92252
rect 119655 92212 119676 92252
rect 119716 92212 119737 92252
rect 119823 92212 119840 92252
rect 119880 92212 119889 92252
rect 119503 92189 119569 92212
rect 119655 92189 119737 92212
rect 119823 92189 119889 92212
rect 119503 92170 119889 92189
rect 134623 92275 135009 92294
rect 134623 92252 134689 92275
rect 134775 92252 134857 92275
rect 134943 92252 135009 92275
rect 134623 92212 134632 92252
rect 134672 92212 134689 92252
rect 134775 92212 134796 92252
rect 134836 92212 134857 92252
rect 134943 92212 134960 92252
rect 135000 92212 135009 92252
rect 134623 92189 134689 92212
rect 134775 92189 134857 92212
rect 134943 92189 135009 92212
rect 134623 92170 135009 92189
rect 149743 92275 150129 92294
rect 149743 92252 149809 92275
rect 149895 92252 149977 92275
rect 150063 92252 150129 92275
rect 149743 92212 149752 92252
rect 149792 92212 149809 92252
rect 149895 92212 149916 92252
rect 149956 92212 149977 92252
rect 150063 92212 150080 92252
rect 150120 92212 150129 92252
rect 149743 92189 149809 92212
rect 149895 92189 149977 92212
rect 150063 92189 150129 92212
rect 149743 92170 150129 92189
rect 75383 91519 75769 91538
rect 75383 91496 75449 91519
rect 75535 91496 75617 91519
rect 75703 91496 75769 91519
rect 75383 91456 75392 91496
rect 75432 91456 75449 91496
rect 75535 91456 75556 91496
rect 75596 91456 75617 91496
rect 75703 91456 75720 91496
rect 75760 91456 75769 91496
rect 75383 91433 75449 91456
rect 75535 91433 75617 91456
rect 75703 91433 75769 91456
rect 75383 91414 75769 91433
rect 90503 91519 90889 91538
rect 90503 91496 90569 91519
rect 90655 91496 90737 91519
rect 90823 91496 90889 91519
rect 90503 91456 90512 91496
rect 90552 91456 90569 91496
rect 90655 91456 90676 91496
rect 90716 91456 90737 91496
rect 90823 91456 90840 91496
rect 90880 91456 90889 91496
rect 90503 91433 90569 91456
rect 90655 91433 90737 91456
rect 90823 91433 90889 91456
rect 90503 91414 90889 91433
rect 105623 91519 106009 91538
rect 105623 91496 105689 91519
rect 105775 91496 105857 91519
rect 105943 91496 106009 91519
rect 105623 91456 105632 91496
rect 105672 91456 105689 91496
rect 105775 91456 105796 91496
rect 105836 91456 105857 91496
rect 105943 91456 105960 91496
rect 106000 91456 106009 91496
rect 105623 91433 105689 91456
rect 105775 91433 105857 91456
rect 105943 91433 106009 91456
rect 105623 91414 106009 91433
rect 120743 91519 121129 91538
rect 120743 91496 120809 91519
rect 120895 91496 120977 91519
rect 121063 91496 121129 91519
rect 120743 91456 120752 91496
rect 120792 91456 120809 91496
rect 120895 91456 120916 91496
rect 120956 91456 120977 91496
rect 121063 91456 121080 91496
rect 121120 91456 121129 91496
rect 120743 91433 120809 91456
rect 120895 91433 120977 91456
rect 121063 91433 121129 91456
rect 120743 91414 121129 91433
rect 135863 91519 136249 91538
rect 135863 91496 135929 91519
rect 136015 91496 136097 91519
rect 136183 91496 136249 91519
rect 135863 91456 135872 91496
rect 135912 91456 135929 91496
rect 136015 91456 136036 91496
rect 136076 91456 136097 91496
rect 136183 91456 136200 91496
rect 136240 91456 136249 91496
rect 135863 91433 135929 91456
rect 136015 91433 136097 91456
rect 136183 91433 136249 91456
rect 135863 91414 136249 91433
rect 150983 91519 151369 91538
rect 150983 91496 151049 91519
rect 151135 91496 151217 91519
rect 151303 91496 151369 91519
rect 150983 91456 150992 91496
rect 151032 91456 151049 91496
rect 151135 91456 151156 91496
rect 151196 91456 151217 91496
rect 151303 91456 151320 91496
rect 151360 91456 151369 91496
rect 150983 91433 151049 91456
rect 151135 91433 151217 91456
rect 151303 91433 151369 91456
rect 150983 91414 151369 91433
rect 74143 90763 74529 90782
rect 74143 90740 74209 90763
rect 74295 90740 74377 90763
rect 74463 90740 74529 90763
rect 74143 90700 74152 90740
rect 74192 90700 74209 90740
rect 74295 90700 74316 90740
rect 74356 90700 74377 90740
rect 74463 90700 74480 90740
rect 74520 90700 74529 90740
rect 74143 90677 74209 90700
rect 74295 90677 74377 90700
rect 74463 90677 74529 90700
rect 74143 90658 74529 90677
rect 89263 90763 89649 90782
rect 89263 90740 89329 90763
rect 89415 90740 89497 90763
rect 89583 90740 89649 90763
rect 89263 90700 89272 90740
rect 89312 90700 89329 90740
rect 89415 90700 89436 90740
rect 89476 90700 89497 90740
rect 89583 90700 89600 90740
rect 89640 90700 89649 90740
rect 89263 90677 89329 90700
rect 89415 90677 89497 90700
rect 89583 90677 89649 90700
rect 89263 90658 89649 90677
rect 104383 90763 104769 90782
rect 104383 90740 104449 90763
rect 104535 90740 104617 90763
rect 104703 90740 104769 90763
rect 104383 90700 104392 90740
rect 104432 90700 104449 90740
rect 104535 90700 104556 90740
rect 104596 90700 104617 90740
rect 104703 90700 104720 90740
rect 104760 90700 104769 90740
rect 104383 90677 104449 90700
rect 104535 90677 104617 90700
rect 104703 90677 104769 90700
rect 104383 90658 104769 90677
rect 119503 90763 119889 90782
rect 119503 90740 119569 90763
rect 119655 90740 119737 90763
rect 119823 90740 119889 90763
rect 119503 90700 119512 90740
rect 119552 90700 119569 90740
rect 119655 90700 119676 90740
rect 119716 90700 119737 90740
rect 119823 90700 119840 90740
rect 119880 90700 119889 90740
rect 119503 90677 119569 90700
rect 119655 90677 119737 90700
rect 119823 90677 119889 90700
rect 119503 90658 119889 90677
rect 134623 90763 135009 90782
rect 134623 90740 134689 90763
rect 134775 90740 134857 90763
rect 134943 90740 135009 90763
rect 134623 90700 134632 90740
rect 134672 90700 134689 90740
rect 134775 90700 134796 90740
rect 134836 90700 134857 90740
rect 134943 90700 134960 90740
rect 135000 90700 135009 90740
rect 134623 90677 134689 90700
rect 134775 90677 134857 90700
rect 134943 90677 135009 90700
rect 134623 90658 135009 90677
rect 149743 90763 150129 90782
rect 149743 90740 149809 90763
rect 149895 90740 149977 90763
rect 150063 90740 150129 90763
rect 149743 90700 149752 90740
rect 149792 90700 149809 90740
rect 149895 90700 149916 90740
rect 149956 90700 149977 90740
rect 150063 90700 150080 90740
rect 150120 90700 150129 90740
rect 149743 90677 149809 90700
rect 149895 90677 149977 90700
rect 150063 90677 150129 90700
rect 149743 90658 150129 90677
rect 75383 90007 75769 90026
rect 75383 89984 75449 90007
rect 75535 89984 75617 90007
rect 75703 89984 75769 90007
rect 75383 89944 75392 89984
rect 75432 89944 75449 89984
rect 75535 89944 75556 89984
rect 75596 89944 75617 89984
rect 75703 89944 75720 89984
rect 75760 89944 75769 89984
rect 75383 89921 75449 89944
rect 75535 89921 75617 89944
rect 75703 89921 75769 89944
rect 75383 89902 75769 89921
rect 90503 90007 90889 90026
rect 90503 89984 90569 90007
rect 90655 89984 90737 90007
rect 90823 89984 90889 90007
rect 90503 89944 90512 89984
rect 90552 89944 90569 89984
rect 90655 89944 90676 89984
rect 90716 89944 90737 89984
rect 90823 89944 90840 89984
rect 90880 89944 90889 89984
rect 90503 89921 90569 89944
rect 90655 89921 90737 89944
rect 90823 89921 90889 89944
rect 90503 89902 90889 89921
rect 105623 90007 106009 90026
rect 105623 89984 105689 90007
rect 105775 89984 105857 90007
rect 105943 89984 106009 90007
rect 105623 89944 105632 89984
rect 105672 89944 105689 89984
rect 105775 89944 105796 89984
rect 105836 89944 105857 89984
rect 105943 89944 105960 89984
rect 106000 89944 106009 89984
rect 105623 89921 105689 89944
rect 105775 89921 105857 89944
rect 105943 89921 106009 89944
rect 105623 89902 106009 89921
rect 120743 90007 121129 90026
rect 120743 89984 120809 90007
rect 120895 89984 120977 90007
rect 121063 89984 121129 90007
rect 120743 89944 120752 89984
rect 120792 89944 120809 89984
rect 120895 89944 120916 89984
rect 120956 89944 120977 89984
rect 121063 89944 121080 89984
rect 121120 89944 121129 89984
rect 120743 89921 120809 89944
rect 120895 89921 120977 89944
rect 121063 89921 121129 89944
rect 120743 89902 121129 89921
rect 135863 90007 136249 90026
rect 135863 89984 135929 90007
rect 136015 89984 136097 90007
rect 136183 89984 136249 90007
rect 135863 89944 135872 89984
rect 135912 89944 135929 89984
rect 136015 89944 136036 89984
rect 136076 89944 136097 89984
rect 136183 89944 136200 89984
rect 136240 89944 136249 89984
rect 135863 89921 135929 89944
rect 136015 89921 136097 89944
rect 136183 89921 136249 89944
rect 135863 89902 136249 89921
rect 150983 90007 151369 90026
rect 150983 89984 151049 90007
rect 151135 89984 151217 90007
rect 151303 89984 151369 90007
rect 150983 89944 150992 89984
rect 151032 89944 151049 89984
rect 151135 89944 151156 89984
rect 151196 89944 151217 89984
rect 151303 89944 151320 89984
rect 151360 89944 151369 89984
rect 150983 89921 151049 89944
rect 151135 89921 151217 89944
rect 151303 89921 151369 89944
rect 150983 89902 151369 89921
rect 74143 89251 74529 89270
rect 74143 89228 74209 89251
rect 74295 89228 74377 89251
rect 74463 89228 74529 89251
rect 74143 89188 74152 89228
rect 74192 89188 74209 89228
rect 74295 89188 74316 89228
rect 74356 89188 74377 89228
rect 74463 89188 74480 89228
rect 74520 89188 74529 89228
rect 74143 89165 74209 89188
rect 74295 89165 74377 89188
rect 74463 89165 74529 89188
rect 74143 89146 74529 89165
rect 89263 89251 89649 89270
rect 89263 89228 89329 89251
rect 89415 89228 89497 89251
rect 89583 89228 89649 89251
rect 89263 89188 89272 89228
rect 89312 89188 89329 89228
rect 89415 89188 89436 89228
rect 89476 89188 89497 89228
rect 89583 89188 89600 89228
rect 89640 89188 89649 89228
rect 89263 89165 89329 89188
rect 89415 89165 89497 89188
rect 89583 89165 89649 89188
rect 89263 89146 89649 89165
rect 104383 89251 104769 89270
rect 104383 89228 104449 89251
rect 104535 89228 104617 89251
rect 104703 89228 104769 89251
rect 104383 89188 104392 89228
rect 104432 89188 104449 89228
rect 104535 89188 104556 89228
rect 104596 89188 104617 89228
rect 104703 89188 104720 89228
rect 104760 89188 104769 89228
rect 104383 89165 104449 89188
rect 104535 89165 104617 89188
rect 104703 89165 104769 89188
rect 104383 89146 104769 89165
rect 119503 89251 119889 89270
rect 119503 89228 119569 89251
rect 119655 89228 119737 89251
rect 119823 89228 119889 89251
rect 119503 89188 119512 89228
rect 119552 89188 119569 89228
rect 119655 89188 119676 89228
rect 119716 89188 119737 89228
rect 119823 89188 119840 89228
rect 119880 89188 119889 89228
rect 119503 89165 119569 89188
rect 119655 89165 119737 89188
rect 119823 89165 119889 89188
rect 119503 89146 119889 89165
rect 134623 89251 135009 89270
rect 134623 89228 134689 89251
rect 134775 89228 134857 89251
rect 134943 89228 135009 89251
rect 134623 89188 134632 89228
rect 134672 89188 134689 89228
rect 134775 89188 134796 89228
rect 134836 89188 134857 89228
rect 134943 89188 134960 89228
rect 135000 89188 135009 89228
rect 134623 89165 134689 89188
rect 134775 89165 134857 89188
rect 134943 89165 135009 89188
rect 134623 89146 135009 89165
rect 149743 89251 150129 89270
rect 149743 89228 149809 89251
rect 149895 89228 149977 89251
rect 150063 89228 150129 89251
rect 149743 89188 149752 89228
rect 149792 89188 149809 89228
rect 149895 89188 149916 89228
rect 149956 89188 149977 89228
rect 150063 89188 150080 89228
rect 150120 89188 150129 89228
rect 149743 89165 149809 89188
rect 149895 89165 149977 89188
rect 150063 89165 150129 89188
rect 149743 89146 150129 89165
rect 75383 88495 75769 88514
rect 75383 88472 75449 88495
rect 75535 88472 75617 88495
rect 75703 88472 75769 88495
rect 75383 88432 75392 88472
rect 75432 88432 75449 88472
rect 75535 88432 75556 88472
rect 75596 88432 75617 88472
rect 75703 88432 75720 88472
rect 75760 88432 75769 88472
rect 75383 88409 75449 88432
rect 75535 88409 75617 88432
rect 75703 88409 75769 88432
rect 75383 88390 75769 88409
rect 90503 88495 90889 88514
rect 90503 88472 90569 88495
rect 90655 88472 90737 88495
rect 90823 88472 90889 88495
rect 90503 88432 90512 88472
rect 90552 88432 90569 88472
rect 90655 88432 90676 88472
rect 90716 88432 90737 88472
rect 90823 88432 90840 88472
rect 90880 88432 90889 88472
rect 90503 88409 90569 88432
rect 90655 88409 90737 88432
rect 90823 88409 90889 88432
rect 90503 88390 90889 88409
rect 105623 88495 106009 88514
rect 105623 88472 105689 88495
rect 105775 88472 105857 88495
rect 105943 88472 106009 88495
rect 105623 88432 105632 88472
rect 105672 88432 105689 88472
rect 105775 88432 105796 88472
rect 105836 88432 105857 88472
rect 105943 88432 105960 88472
rect 106000 88432 106009 88472
rect 105623 88409 105689 88432
rect 105775 88409 105857 88432
rect 105943 88409 106009 88432
rect 105623 88390 106009 88409
rect 120743 88495 121129 88514
rect 120743 88472 120809 88495
rect 120895 88472 120977 88495
rect 121063 88472 121129 88495
rect 120743 88432 120752 88472
rect 120792 88432 120809 88472
rect 120895 88432 120916 88472
rect 120956 88432 120977 88472
rect 121063 88432 121080 88472
rect 121120 88432 121129 88472
rect 120743 88409 120809 88432
rect 120895 88409 120977 88432
rect 121063 88409 121129 88432
rect 120743 88390 121129 88409
rect 135863 88495 136249 88514
rect 135863 88472 135929 88495
rect 136015 88472 136097 88495
rect 136183 88472 136249 88495
rect 135863 88432 135872 88472
rect 135912 88432 135929 88472
rect 136015 88432 136036 88472
rect 136076 88432 136097 88472
rect 136183 88432 136200 88472
rect 136240 88432 136249 88472
rect 135863 88409 135929 88432
rect 136015 88409 136097 88432
rect 136183 88409 136249 88432
rect 135863 88390 136249 88409
rect 150983 88495 151369 88514
rect 150983 88472 151049 88495
rect 151135 88472 151217 88495
rect 151303 88472 151369 88495
rect 150983 88432 150992 88472
rect 151032 88432 151049 88472
rect 151135 88432 151156 88472
rect 151196 88432 151217 88472
rect 151303 88432 151320 88472
rect 151360 88432 151369 88472
rect 150983 88409 151049 88432
rect 151135 88409 151217 88432
rect 151303 88409 151369 88432
rect 150983 88390 151369 88409
rect 74143 87739 74529 87758
rect 74143 87716 74209 87739
rect 74295 87716 74377 87739
rect 74463 87716 74529 87739
rect 74143 87676 74152 87716
rect 74192 87676 74209 87716
rect 74295 87676 74316 87716
rect 74356 87676 74377 87716
rect 74463 87676 74480 87716
rect 74520 87676 74529 87716
rect 74143 87653 74209 87676
rect 74295 87653 74377 87676
rect 74463 87653 74529 87676
rect 74143 87634 74529 87653
rect 89263 87739 89649 87758
rect 89263 87716 89329 87739
rect 89415 87716 89497 87739
rect 89583 87716 89649 87739
rect 89263 87676 89272 87716
rect 89312 87676 89329 87716
rect 89415 87676 89436 87716
rect 89476 87676 89497 87716
rect 89583 87676 89600 87716
rect 89640 87676 89649 87716
rect 89263 87653 89329 87676
rect 89415 87653 89497 87676
rect 89583 87653 89649 87676
rect 89263 87634 89649 87653
rect 104383 87739 104769 87758
rect 104383 87716 104449 87739
rect 104535 87716 104617 87739
rect 104703 87716 104769 87739
rect 104383 87676 104392 87716
rect 104432 87676 104449 87716
rect 104535 87676 104556 87716
rect 104596 87676 104617 87716
rect 104703 87676 104720 87716
rect 104760 87676 104769 87716
rect 104383 87653 104449 87676
rect 104535 87653 104617 87676
rect 104703 87653 104769 87676
rect 104383 87634 104769 87653
rect 119503 87739 119889 87758
rect 119503 87716 119569 87739
rect 119655 87716 119737 87739
rect 119823 87716 119889 87739
rect 119503 87676 119512 87716
rect 119552 87676 119569 87716
rect 119655 87676 119676 87716
rect 119716 87676 119737 87716
rect 119823 87676 119840 87716
rect 119880 87676 119889 87716
rect 119503 87653 119569 87676
rect 119655 87653 119737 87676
rect 119823 87653 119889 87676
rect 119503 87634 119889 87653
rect 134623 87739 135009 87758
rect 134623 87716 134689 87739
rect 134775 87716 134857 87739
rect 134943 87716 135009 87739
rect 134623 87676 134632 87716
rect 134672 87676 134689 87716
rect 134775 87676 134796 87716
rect 134836 87676 134857 87716
rect 134943 87676 134960 87716
rect 135000 87676 135009 87716
rect 134623 87653 134689 87676
rect 134775 87653 134857 87676
rect 134943 87653 135009 87676
rect 134623 87634 135009 87653
rect 149743 87739 150129 87758
rect 149743 87716 149809 87739
rect 149895 87716 149977 87739
rect 150063 87716 150129 87739
rect 149743 87676 149752 87716
rect 149792 87676 149809 87716
rect 149895 87676 149916 87716
rect 149956 87676 149977 87716
rect 150063 87676 150080 87716
rect 150120 87676 150129 87716
rect 149743 87653 149809 87676
rect 149895 87653 149977 87676
rect 150063 87653 150129 87676
rect 149743 87634 150129 87653
rect 75383 86983 75769 87002
rect 75383 86960 75449 86983
rect 75535 86960 75617 86983
rect 75703 86960 75769 86983
rect 75383 86920 75392 86960
rect 75432 86920 75449 86960
rect 75535 86920 75556 86960
rect 75596 86920 75617 86960
rect 75703 86920 75720 86960
rect 75760 86920 75769 86960
rect 75383 86897 75449 86920
rect 75535 86897 75617 86920
rect 75703 86897 75769 86920
rect 75383 86878 75769 86897
rect 90503 86983 90889 87002
rect 90503 86960 90569 86983
rect 90655 86960 90737 86983
rect 90823 86960 90889 86983
rect 90503 86920 90512 86960
rect 90552 86920 90569 86960
rect 90655 86920 90676 86960
rect 90716 86920 90737 86960
rect 90823 86920 90840 86960
rect 90880 86920 90889 86960
rect 90503 86897 90569 86920
rect 90655 86897 90737 86920
rect 90823 86897 90889 86920
rect 90503 86878 90889 86897
rect 105623 86983 106009 87002
rect 105623 86960 105689 86983
rect 105775 86960 105857 86983
rect 105943 86960 106009 86983
rect 105623 86920 105632 86960
rect 105672 86920 105689 86960
rect 105775 86920 105796 86960
rect 105836 86920 105857 86960
rect 105943 86920 105960 86960
rect 106000 86920 106009 86960
rect 105623 86897 105689 86920
rect 105775 86897 105857 86920
rect 105943 86897 106009 86920
rect 105623 86878 106009 86897
rect 120743 86983 121129 87002
rect 120743 86960 120809 86983
rect 120895 86960 120977 86983
rect 121063 86960 121129 86983
rect 120743 86920 120752 86960
rect 120792 86920 120809 86960
rect 120895 86920 120916 86960
rect 120956 86920 120977 86960
rect 121063 86920 121080 86960
rect 121120 86920 121129 86960
rect 120743 86897 120809 86920
rect 120895 86897 120977 86920
rect 121063 86897 121129 86920
rect 120743 86878 121129 86897
rect 135863 86983 136249 87002
rect 135863 86960 135929 86983
rect 136015 86960 136097 86983
rect 136183 86960 136249 86983
rect 135863 86920 135872 86960
rect 135912 86920 135929 86960
rect 136015 86920 136036 86960
rect 136076 86920 136097 86960
rect 136183 86920 136200 86960
rect 136240 86920 136249 86960
rect 135863 86897 135929 86920
rect 136015 86897 136097 86920
rect 136183 86897 136249 86920
rect 135863 86878 136249 86897
rect 150983 86983 151369 87002
rect 150983 86960 151049 86983
rect 151135 86960 151217 86983
rect 151303 86960 151369 86983
rect 150983 86920 150992 86960
rect 151032 86920 151049 86960
rect 151135 86920 151156 86960
rect 151196 86920 151217 86960
rect 151303 86920 151320 86960
rect 151360 86920 151369 86960
rect 150983 86897 151049 86920
rect 151135 86897 151217 86920
rect 151303 86897 151369 86920
rect 150983 86878 151369 86897
rect 74143 86227 74529 86246
rect 74143 86204 74209 86227
rect 74295 86204 74377 86227
rect 74463 86204 74529 86227
rect 74143 86164 74152 86204
rect 74192 86164 74209 86204
rect 74295 86164 74316 86204
rect 74356 86164 74377 86204
rect 74463 86164 74480 86204
rect 74520 86164 74529 86204
rect 74143 86141 74209 86164
rect 74295 86141 74377 86164
rect 74463 86141 74529 86164
rect 74143 86122 74529 86141
rect 89263 86227 89649 86246
rect 89263 86204 89329 86227
rect 89415 86204 89497 86227
rect 89583 86204 89649 86227
rect 89263 86164 89272 86204
rect 89312 86164 89329 86204
rect 89415 86164 89436 86204
rect 89476 86164 89497 86204
rect 89583 86164 89600 86204
rect 89640 86164 89649 86204
rect 89263 86141 89329 86164
rect 89415 86141 89497 86164
rect 89583 86141 89649 86164
rect 89263 86122 89649 86141
rect 104383 86227 104769 86246
rect 104383 86204 104449 86227
rect 104535 86204 104617 86227
rect 104703 86204 104769 86227
rect 104383 86164 104392 86204
rect 104432 86164 104449 86204
rect 104535 86164 104556 86204
rect 104596 86164 104617 86204
rect 104703 86164 104720 86204
rect 104760 86164 104769 86204
rect 104383 86141 104449 86164
rect 104535 86141 104617 86164
rect 104703 86141 104769 86164
rect 104383 86122 104769 86141
rect 119503 86227 119889 86246
rect 119503 86204 119569 86227
rect 119655 86204 119737 86227
rect 119823 86204 119889 86227
rect 119503 86164 119512 86204
rect 119552 86164 119569 86204
rect 119655 86164 119676 86204
rect 119716 86164 119737 86204
rect 119823 86164 119840 86204
rect 119880 86164 119889 86204
rect 119503 86141 119569 86164
rect 119655 86141 119737 86164
rect 119823 86141 119889 86164
rect 119503 86122 119889 86141
rect 134623 86227 135009 86246
rect 134623 86204 134689 86227
rect 134775 86204 134857 86227
rect 134943 86204 135009 86227
rect 134623 86164 134632 86204
rect 134672 86164 134689 86204
rect 134775 86164 134796 86204
rect 134836 86164 134857 86204
rect 134943 86164 134960 86204
rect 135000 86164 135009 86204
rect 134623 86141 134689 86164
rect 134775 86141 134857 86164
rect 134943 86141 135009 86164
rect 134623 86122 135009 86141
rect 149743 86227 150129 86246
rect 149743 86204 149809 86227
rect 149895 86204 149977 86227
rect 150063 86204 150129 86227
rect 149743 86164 149752 86204
rect 149792 86164 149809 86204
rect 149895 86164 149916 86204
rect 149956 86164 149977 86204
rect 150063 86164 150080 86204
rect 150120 86164 150129 86204
rect 149743 86141 149809 86164
rect 149895 86141 149977 86164
rect 150063 86141 150129 86164
rect 149743 86122 150129 86141
rect 75383 85471 75769 85490
rect 75383 85448 75449 85471
rect 75535 85448 75617 85471
rect 75703 85448 75769 85471
rect 75383 85408 75392 85448
rect 75432 85408 75449 85448
rect 75535 85408 75556 85448
rect 75596 85408 75617 85448
rect 75703 85408 75720 85448
rect 75760 85408 75769 85448
rect 75383 85385 75449 85408
rect 75535 85385 75617 85408
rect 75703 85385 75769 85408
rect 75383 85366 75769 85385
rect 90503 85471 90889 85490
rect 90503 85448 90569 85471
rect 90655 85448 90737 85471
rect 90823 85448 90889 85471
rect 90503 85408 90512 85448
rect 90552 85408 90569 85448
rect 90655 85408 90676 85448
rect 90716 85408 90737 85448
rect 90823 85408 90840 85448
rect 90880 85408 90889 85448
rect 90503 85385 90569 85408
rect 90655 85385 90737 85408
rect 90823 85385 90889 85408
rect 90503 85366 90889 85385
rect 105623 85471 106009 85490
rect 105623 85448 105689 85471
rect 105775 85448 105857 85471
rect 105943 85448 106009 85471
rect 105623 85408 105632 85448
rect 105672 85408 105689 85448
rect 105775 85408 105796 85448
rect 105836 85408 105857 85448
rect 105943 85408 105960 85448
rect 106000 85408 106009 85448
rect 105623 85385 105689 85408
rect 105775 85385 105857 85408
rect 105943 85385 106009 85408
rect 105623 85366 106009 85385
rect 120743 85471 121129 85490
rect 120743 85448 120809 85471
rect 120895 85448 120977 85471
rect 121063 85448 121129 85471
rect 120743 85408 120752 85448
rect 120792 85408 120809 85448
rect 120895 85408 120916 85448
rect 120956 85408 120977 85448
rect 121063 85408 121080 85448
rect 121120 85408 121129 85448
rect 120743 85385 120809 85408
rect 120895 85385 120977 85408
rect 121063 85385 121129 85408
rect 120743 85366 121129 85385
rect 135863 85471 136249 85490
rect 135863 85448 135929 85471
rect 136015 85448 136097 85471
rect 136183 85448 136249 85471
rect 135863 85408 135872 85448
rect 135912 85408 135929 85448
rect 136015 85408 136036 85448
rect 136076 85408 136097 85448
rect 136183 85408 136200 85448
rect 136240 85408 136249 85448
rect 135863 85385 135929 85408
rect 136015 85385 136097 85408
rect 136183 85385 136249 85408
rect 135863 85366 136249 85385
rect 150983 85471 151369 85490
rect 150983 85448 151049 85471
rect 151135 85448 151217 85471
rect 151303 85448 151369 85471
rect 150983 85408 150992 85448
rect 151032 85408 151049 85448
rect 151135 85408 151156 85448
rect 151196 85408 151217 85448
rect 151303 85408 151320 85448
rect 151360 85408 151369 85448
rect 150983 85385 151049 85408
rect 151135 85385 151217 85408
rect 151303 85385 151369 85408
rect 150983 85366 151369 85385
rect 74143 84715 74529 84734
rect 74143 84692 74209 84715
rect 74295 84692 74377 84715
rect 74463 84692 74529 84715
rect 74143 84652 74152 84692
rect 74192 84652 74209 84692
rect 74295 84652 74316 84692
rect 74356 84652 74377 84692
rect 74463 84652 74480 84692
rect 74520 84652 74529 84692
rect 74143 84629 74209 84652
rect 74295 84629 74377 84652
rect 74463 84629 74529 84652
rect 74143 84610 74529 84629
rect 89263 84715 89649 84734
rect 89263 84692 89329 84715
rect 89415 84692 89497 84715
rect 89583 84692 89649 84715
rect 89263 84652 89272 84692
rect 89312 84652 89329 84692
rect 89415 84652 89436 84692
rect 89476 84652 89497 84692
rect 89583 84652 89600 84692
rect 89640 84652 89649 84692
rect 89263 84629 89329 84652
rect 89415 84629 89497 84652
rect 89583 84629 89649 84652
rect 89263 84610 89649 84629
rect 104383 84715 104769 84734
rect 104383 84692 104449 84715
rect 104535 84692 104617 84715
rect 104703 84692 104769 84715
rect 104383 84652 104392 84692
rect 104432 84652 104449 84692
rect 104535 84652 104556 84692
rect 104596 84652 104617 84692
rect 104703 84652 104720 84692
rect 104760 84652 104769 84692
rect 104383 84629 104449 84652
rect 104535 84629 104617 84652
rect 104703 84629 104769 84652
rect 104383 84610 104769 84629
rect 119503 84715 119889 84734
rect 119503 84692 119569 84715
rect 119655 84692 119737 84715
rect 119823 84692 119889 84715
rect 119503 84652 119512 84692
rect 119552 84652 119569 84692
rect 119655 84652 119676 84692
rect 119716 84652 119737 84692
rect 119823 84652 119840 84692
rect 119880 84652 119889 84692
rect 119503 84629 119569 84652
rect 119655 84629 119737 84652
rect 119823 84629 119889 84652
rect 119503 84610 119889 84629
rect 134623 84715 135009 84734
rect 134623 84692 134689 84715
rect 134775 84692 134857 84715
rect 134943 84692 135009 84715
rect 134623 84652 134632 84692
rect 134672 84652 134689 84692
rect 134775 84652 134796 84692
rect 134836 84652 134857 84692
rect 134943 84652 134960 84692
rect 135000 84652 135009 84692
rect 134623 84629 134689 84652
rect 134775 84629 134857 84652
rect 134943 84629 135009 84652
rect 134623 84610 135009 84629
rect 149743 84715 150129 84734
rect 149743 84692 149809 84715
rect 149895 84692 149977 84715
rect 150063 84692 150129 84715
rect 149743 84652 149752 84692
rect 149792 84652 149809 84692
rect 149895 84652 149916 84692
rect 149956 84652 149977 84692
rect 150063 84652 150080 84692
rect 150120 84652 150129 84692
rect 149743 84629 149809 84652
rect 149895 84629 149977 84652
rect 150063 84629 150129 84652
rect 149743 84610 150129 84629
rect 75383 83959 75769 83978
rect 75383 83936 75449 83959
rect 75535 83936 75617 83959
rect 75703 83936 75769 83959
rect 75383 83896 75392 83936
rect 75432 83896 75449 83936
rect 75535 83896 75556 83936
rect 75596 83896 75617 83936
rect 75703 83896 75720 83936
rect 75760 83896 75769 83936
rect 75383 83873 75449 83896
rect 75535 83873 75617 83896
rect 75703 83873 75769 83896
rect 75383 83854 75769 83873
rect 90503 83959 90889 83978
rect 90503 83936 90569 83959
rect 90655 83936 90737 83959
rect 90823 83936 90889 83959
rect 90503 83896 90512 83936
rect 90552 83896 90569 83936
rect 90655 83896 90676 83936
rect 90716 83896 90737 83936
rect 90823 83896 90840 83936
rect 90880 83896 90889 83936
rect 90503 83873 90569 83896
rect 90655 83873 90737 83896
rect 90823 83873 90889 83896
rect 90503 83854 90889 83873
rect 105623 83959 106009 83978
rect 105623 83936 105689 83959
rect 105775 83936 105857 83959
rect 105943 83936 106009 83959
rect 105623 83896 105632 83936
rect 105672 83896 105689 83936
rect 105775 83896 105796 83936
rect 105836 83896 105857 83936
rect 105943 83896 105960 83936
rect 106000 83896 106009 83936
rect 105623 83873 105689 83896
rect 105775 83873 105857 83896
rect 105943 83873 106009 83896
rect 105623 83854 106009 83873
rect 120743 83959 121129 83978
rect 120743 83936 120809 83959
rect 120895 83936 120977 83959
rect 121063 83936 121129 83959
rect 120743 83896 120752 83936
rect 120792 83896 120809 83936
rect 120895 83896 120916 83936
rect 120956 83896 120977 83936
rect 121063 83896 121080 83936
rect 121120 83896 121129 83936
rect 120743 83873 120809 83896
rect 120895 83873 120977 83896
rect 121063 83873 121129 83896
rect 120743 83854 121129 83873
rect 135863 83959 136249 83978
rect 135863 83936 135929 83959
rect 136015 83936 136097 83959
rect 136183 83936 136249 83959
rect 135863 83896 135872 83936
rect 135912 83896 135929 83936
rect 136015 83896 136036 83936
rect 136076 83896 136097 83936
rect 136183 83896 136200 83936
rect 136240 83896 136249 83936
rect 135863 83873 135929 83896
rect 136015 83873 136097 83896
rect 136183 83873 136249 83896
rect 135863 83854 136249 83873
rect 150983 83959 151369 83978
rect 150983 83936 151049 83959
rect 151135 83936 151217 83959
rect 151303 83936 151369 83959
rect 150983 83896 150992 83936
rect 151032 83896 151049 83936
rect 151135 83896 151156 83936
rect 151196 83896 151217 83936
rect 151303 83896 151320 83936
rect 151360 83896 151369 83936
rect 150983 83873 151049 83896
rect 151135 83873 151217 83896
rect 151303 83873 151369 83896
rect 150983 83854 151369 83873
rect 74143 83203 74529 83222
rect 74143 83180 74209 83203
rect 74295 83180 74377 83203
rect 74463 83180 74529 83203
rect 74143 83140 74152 83180
rect 74192 83140 74209 83180
rect 74295 83140 74316 83180
rect 74356 83140 74377 83180
rect 74463 83140 74480 83180
rect 74520 83140 74529 83180
rect 74143 83117 74209 83140
rect 74295 83117 74377 83140
rect 74463 83117 74529 83140
rect 74143 83098 74529 83117
rect 89263 83203 89649 83222
rect 89263 83180 89329 83203
rect 89415 83180 89497 83203
rect 89583 83180 89649 83203
rect 89263 83140 89272 83180
rect 89312 83140 89329 83180
rect 89415 83140 89436 83180
rect 89476 83140 89497 83180
rect 89583 83140 89600 83180
rect 89640 83140 89649 83180
rect 89263 83117 89329 83140
rect 89415 83117 89497 83140
rect 89583 83117 89649 83140
rect 89263 83098 89649 83117
rect 104383 83203 104769 83222
rect 104383 83180 104449 83203
rect 104535 83180 104617 83203
rect 104703 83180 104769 83203
rect 104383 83140 104392 83180
rect 104432 83140 104449 83180
rect 104535 83140 104556 83180
rect 104596 83140 104617 83180
rect 104703 83140 104720 83180
rect 104760 83140 104769 83180
rect 104383 83117 104449 83140
rect 104535 83117 104617 83140
rect 104703 83117 104769 83140
rect 104383 83098 104769 83117
rect 119503 83203 119889 83222
rect 119503 83180 119569 83203
rect 119655 83180 119737 83203
rect 119823 83180 119889 83203
rect 119503 83140 119512 83180
rect 119552 83140 119569 83180
rect 119655 83140 119676 83180
rect 119716 83140 119737 83180
rect 119823 83140 119840 83180
rect 119880 83140 119889 83180
rect 119503 83117 119569 83140
rect 119655 83117 119737 83140
rect 119823 83117 119889 83140
rect 119503 83098 119889 83117
rect 134623 83203 135009 83222
rect 134623 83180 134689 83203
rect 134775 83180 134857 83203
rect 134943 83180 135009 83203
rect 134623 83140 134632 83180
rect 134672 83140 134689 83180
rect 134775 83140 134796 83180
rect 134836 83140 134857 83180
rect 134943 83140 134960 83180
rect 135000 83140 135009 83180
rect 134623 83117 134689 83140
rect 134775 83117 134857 83140
rect 134943 83117 135009 83140
rect 134623 83098 135009 83117
rect 149743 83203 150129 83222
rect 149743 83180 149809 83203
rect 149895 83180 149977 83203
rect 150063 83180 150129 83203
rect 149743 83140 149752 83180
rect 149792 83140 149809 83180
rect 149895 83140 149916 83180
rect 149956 83140 149977 83180
rect 150063 83140 150080 83180
rect 150120 83140 150129 83180
rect 149743 83117 149809 83140
rect 149895 83117 149977 83140
rect 150063 83117 150129 83140
rect 149743 83098 150129 83117
rect 75383 82447 75769 82466
rect 75383 82424 75449 82447
rect 75535 82424 75617 82447
rect 75703 82424 75769 82447
rect 75383 82384 75392 82424
rect 75432 82384 75449 82424
rect 75535 82384 75556 82424
rect 75596 82384 75617 82424
rect 75703 82384 75720 82424
rect 75760 82384 75769 82424
rect 75383 82361 75449 82384
rect 75535 82361 75617 82384
rect 75703 82361 75769 82384
rect 75383 82342 75769 82361
rect 90503 82447 90889 82466
rect 90503 82424 90569 82447
rect 90655 82424 90737 82447
rect 90823 82424 90889 82447
rect 90503 82384 90512 82424
rect 90552 82384 90569 82424
rect 90655 82384 90676 82424
rect 90716 82384 90737 82424
rect 90823 82384 90840 82424
rect 90880 82384 90889 82424
rect 90503 82361 90569 82384
rect 90655 82361 90737 82384
rect 90823 82361 90889 82384
rect 90503 82342 90889 82361
rect 105623 82447 106009 82466
rect 105623 82424 105689 82447
rect 105775 82424 105857 82447
rect 105943 82424 106009 82447
rect 105623 82384 105632 82424
rect 105672 82384 105689 82424
rect 105775 82384 105796 82424
rect 105836 82384 105857 82424
rect 105943 82384 105960 82424
rect 106000 82384 106009 82424
rect 105623 82361 105689 82384
rect 105775 82361 105857 82384
rect 105943 82361 106009 82384
rect 105623 82342 106009 82361
rect 120743 82447 121129 82466
rect 120743 82424 120809 82447
rect 120895 82424 120977 82447
rect 121063 82424 121129 82447
rect 120743 82384 120752 82424
rect 120792 82384 120809 82424
rect 120895 82384 120916 82424
rect 120956 82384 120977 82424
rect 121063 82384 121080 82424
rect 121120 82384 121129 82424
rect 120743 82361 120809 82384
rect 120895 82361 120977 82384
rect 121063 82361 121129 82384
rect 120743 82342 121129 82361
rect 135863 82447 136249 82466
rect 135863 82424 135929 82447
rect 136015 82424 136097 82447
rect 136183 82424 136249 82447
rect 135863 82384 135872 82424
rect 135912 82384 135929 82424
rect 136015 82384 136036 82424
rect 136076 82384 136097 82424
rect 136183 82384 136200 82424
rect 136240 82384 136249 82424
rect 135863 82361 135929 82384
rect 136015 82361 136097 82384
rect 136183 82361 136249 82384
rect 135863 82342 136249 82361
rect 150983 82447 151369 82466
rect 150983 82424 151049 82447
rect 151135 82424 151217 82447
rect 151303 82424 151369 82447
rect 150983 82384 150992 82424
rect 151032 82384 151049 82424
rect 151135 82384 151156 82424
rect 151196 82384 151217 82424
rect 151303 82384 151320 82424
rect 151360 82384 151369 82424
rect 150983 82361 151049 82384
rect 151135 82361 151217 82384
rect 151303 82361 151369 82384
rect 150983 82342 151369 82361
rect 74143 81691 74529 81710
rect 74143 81668 74209 81691
rect 74295 81668 74377 81691
rect 74463 81668 74529 81691
rect 74143 81628 74152 81668
rect 74192 81628 74209 81668
rect 74295 81628 74316 81668
rect 74356 81628 74377 81668
rect 74463 81628 74480 81668
rect 74520 81628 74529 81668
rect 74143 81605 74209 81628
rect 74295 81605 74377 81628
rect 74463 81605 74529 81628
rect 74143 81586 74529 81605
rect 89263 81691 89649 81710
rect 89263 81668 89329 81691
rect 89415 81668 89497 81691
rect 89583 81668 89649 81691
rect 89263 81628 89272 81668
rect 89312 81628 89329 81668
rect 89415 81628 89436 81668
rect 89476 81628 89497 81668
rect 89583 81628 89600 81668
rect 89640 81628 89649 81668
rect 89263 81605 89329 81628
rect 89415 81605 89497 81628
rect 89583 81605 89649 81628
rect 89263 81586 89649 81605
rect 104383 81691 104769 81710
rect 104383 81668 104449 81691
rect 104535 81668 104617 81691
rect 104703 81668 104769 81691
rect 104383 81628 104392 81668
rect 104432 81628 104449 81668
rect 104535 81628 104556 81668
rect 104596 81628 104617 81668
rect 104703 81628 104720 81668
rect 104760 81628 104769 81668
rect 104383 81605 104449 81628
rect 104535 81605 104617 81628
rect 104703 81605 104769 81628
rect 104383 81586 104769 81605
rect 119503 81691 119889 81710
rect 119503 81668 119569 81691
rect 119655 81668 119737 81691
rect 119823 81668 119889 81691
rect 119503 81628 119512 81668
rect 119552 81628 119569 81668
rect 119655 81628 119676 81668
rect 119716 81628 119737 81668
rect 119823 81628 119840 81668
rect 119880 81628 119889 81668
rect 119503 81605 119569 81628
rect 119655 81605 119737 81628
rect 119823 81605 119889 81628
rect 119503 81586 119889 81605
rect 134623 81691 135009 81710
rect 134623 81668 134689 81691
rect 134775 81668 134857 81691
rect 134943 81668 135009 81691
rect 134623 81628 134632 81668
rect 134672 81628 134689 81668
rect 134775 81628 134796 81668
rect 134836 81628 134857 81668
rect 134943 81628 134960 81668
rect 135000 81628 135009 81668
rect 134623 81605 134689 81628
rect 134775 81605 134857 81628
rect 134943 81605 135009 81628
rect 134623 81586 135009 81605
rect 149743 81691 150129 81710
rect 149743 81668 149809 81691
rect 149895 81668 149977 81691
rect 150063 81668 150129 81691
rect 149743 81628 149752 81668
rect 149792 81628 149809 81668
rect 149895 81628 149916 81668
rect 149956 81628 149977 81668
rect 150063 81628 150080 81668
rect 150120 81628 150129 81668
rect 149743 81605 149809 81628
rect 149895 81605 149977 81628
rect 150063 81605 150129 81628
rect 149743 81586 150129 81605
rect 75383 80935 75769 80954
rect 75383 80912 75449 80935
rect 75535 80912 75617 80935
rect 75703 80912 75769 80935
rect 75383 80872 75392 80912
rect 75432 80872 75449 80912
rect 75535 80872 75556 80912
rect 75596 80872 75617 80912
rect 75703 80872 75720 80912
rect 75760 80872 75769 80912
rect 75383 80849 75449 80872
rect 75535 80849 75617 80872
rect 75703 80849 75769 80872
rect 75383 80830 75769 80849
rect 90503 80935 90889 80954
rect 90503 80912 90569 80935
rect 90655 80912 90737 80935
rect 90823 80912 90889 80935
rect 90503 80872 90512 80912
rect 90552 80872 90569 80912
rect 90655 80872 90676 80912
rect 90716 80872 90737 80912
rect 90823 80872 90840 80912
rect 90880 80872 90889 80912
rect 90503 80849 90569 80872
rect 90655 80849 90737 80872
rect 90823 80849 90889 80872
rect 90503 80830 90889 80849
rect 105623 80935 106009 80954
rect 105623 80912 105689 80935
rect 105775 80912 105857 80935
rect 105943 80912 106009 80935
rect 105623 80872 105632 80912
rect 105672 80872 105689 80912
rect 105775 80872 105796 80912
rect 105836 80872 105857 80912
rect 105943 80872 105960 80912
rect 106000 80872 106009 80912
rect 105623 80849 105689 80872
rect 105775 80849 105857 80872
rect 105943 80849 106009 80872
rect 105623 80830 106009 80849
rect 120743 80935 121129 80954
rect 120743 80912 120809 80935
rect 120895 80912 120977 80935
rect 121063 80912 121129 80935
rect 120743 80872 120752 80912
rect 120792 80872 120809 80912
rect 120895 80872 120916 80912
rect 120956 80872 120977 80912
rect 121063 80872 121080 80912
rect 121120 80872 121129 80912
rect 120743 80849 120809 80872
rect 120895 80849 120977 80872
rect 121063 80849 121129 80872
rect 120743 80830 121129 80849
rect 135863 80935 136249 80954
rect 135863 80912 135929 80935
rect 136015 80912 136097 80935
rect 136183 80912 136249 80935
rect 135863 80872 135872 80912
rect 135912 80872 135929 80912
rect 136015 80872 136036 80912
rect 136076 80872 136097 80912
rect 136183 80872 136200 80912
rect 136240 80872 136249 80912
rect 135863 80849 135929 80872
rect 136015 80849 136097 80872
rect 136183 80849 136249 80872
rect 135863 80830 136249 80849
rect 150983 80935 151369 80954
rect 150983 80912 151049 80935
rect 151135 80912 151217 80935
rect 151303 80912 151369 80935
rect 150983 80872 150992 80912
rect 151032 80872 151049 80912
rect 151135 80872 151156 80912
rect 151196 80872 151217 80912
rect 151303 80872 151320 80912
rect 151360 80872 151369 80912
rect 150983 80849 151049 80872
rect 151135 80849 151217 80872
rect 151303 80849 151369 80872
rect 150983 80830 151369 80849
rect 74143 80179 74529 80198
rect 74143 80156 74209 80179
rect 74295 80156 74377 80179
rect 74463 80156 74529 80179
rect 74143 80116 74152 80156
rect 74192 80116 74209 80156
rect 74295 80116 74316 80156
rect 74356 80116 74377 80156
rect 74463 80116 74480 80156
rect 74520 80116 74529 80156
rect 74143 80093 74209 80116
rect 74295 80093 74377 80116
rect 74463 80093 74529 80116
rect 74143 80074 74529 80093
rect 89263 80179 89649 80198
rect 89263 80156 89329 80179
rect 89415 80156 89497 80179
rect 89583 80156 89649 80179
rect 89263 80116 89272 80156
rect 89312 80116 89329 80156
rect 89415 80116 89436 80156
rect 89476 80116 89497 80156
rect 89583 80116 89600 80156
rect 89640 80116 89649 80156
rect 89263 80093 89329 80116
rect 89415 80093 89497 80116
rect 89583 80093 89649 80116
rect 89263 80074 89649 80093
rect 104383 80179 104769 80198
rect 104383 80156 104449 80179
rect 104535 80156 104617 80179
rect 104703 80156 104769 80179
rect 104383 80116 104392 80156
rect 104432 80116 104449 80156
rect 104535 80116 104556 80156
rect 104596 80116 104617 80156
rect 104703 80116 104720 80156
rect 104760 80116 104769 80156
rect 104383 80093 104449 80116
rect 104535 80093 104617 80116
rect 104703 80093 104769 80116
rect 104383 80074 104769 80093
rect 119503 80179 119889 80198
rect 119503 80156 119569 80179
rect 119655 80156 119737 80179
rect 119823 80156 119889 80179
rect 119503 80116 119512 80156
rect 119552 80116 119569 80156
rect 119655 80116 119676 80156
rect 119716 80116 119737 80156
rect 119823 80116 119840 80156
rect 119880 80116 119889 80156
rect 119503 80093 119569 80116
rect 119655 80093 119737 80116
rect 119823 80093 119889 80116
rect 119503 80074 119889 80093
rect 134623 80179 135009 80198
rect 134623 80156 134689 80179
rect 134775 80156 134857 80179
rect 134943 80156 135009 80179
rect 134623 80116 134632 80156
rect 134672 80116 134689 80156
rect 134775 80116 134796 80156
rect 134836 80116 134857 80156
rect 134943 80116 134960 80156
rect 135000 80116 135009 80156
rect 134623 80093 134689 80116
rect 134775 80093 134857 80116
rect 134943 80093 135009 80116
rect 134623 80074 135009 80093
rect 149743 80179 150129 80198
rect 149743 80156 149809 80179
rect 149895 80156 149977 80179
rect 150063 80156 150129 80179
rect 149743 80116 149752 80156
rect 149792 80116 149809 80156
rect 149895 80116 149916 80156
rect 149956 80116 149977 80156
rect 150063 80116 150080 80156
rect 150120 80116 150129 80156
rect 149743 80093 149809 80116
rect 149895 80093 149977 80116
rect 150063 80093 150129 80116
rect 149743 80074 150129 80093
rect 75383 79423 75769 79442
rect 75383 79400 75449 79423
rect 75535 79400 75617 79423
rect 75703 79400 75769 79423
rect 75383 79360 75392 79400
rect 75432 79360 75449 79400
rect 75535 79360 75556 79400
rect 75596 79360 75617 79400
rect 75703 79360 75720 79400
rect 75760 79360 75769 79400
rect 75383 79337 75449 79360
rect 75535 79337 75617 79360
rect 75703 79337 75769 79360
rect 75383 79318 75769 79337
rect 90503 79423 90889 79442
rect 90503 79400 90569 79423
rect 90655 79400 90737 79423
rect 90823 79400 90889 79423
rect 90503 79360 90512 79400
rect 90552 79360 90569 79400
rect 90655 79360 90676 79400
rect 90716 79360 90737 79400
rect 90823 79360 90840 79400
rect 90880 79360 90889 79400
rect 90503 79337 90569 79360
rect 90655 79337 90737 79360
rect 90823 79337 90889 79360
rect 90503 79318 90889 79337
rect 105623 79423 106009 79442
rect 105623 79400 105689 79423
rect 105775 79400 105857 79423
rect 105943 79400 106009 79423
rect 105623 79360 105632 79400
rect 105672 79360 105689 79400
rect 105775 79360 105796 79400
rect 105836 79360 105857 79400
rect 105943 79360 105960 79400
rect 106000 79360 106009 79400
rect 105623 79337 105689 79360
rect 105775 79337 105857 79360
rect 105943 79337 106009 79360
rect 105623 79318 106009 79337
rect 120743 79423 121129 79442
rect 120743 79400 120809 79423
rect 120895 79400 120977 79423
rect 121063 79400 121129 79423
rect 120743 79360 120752 79400
rect 120792 79360 120809 79400
rect 120895 79360 120916 79400
rect 120956 79360 120977 79400
rect 121063 79360 121080 79400
rect 121120 79360 121129 79400
rect 120743 79337 120809 79360
rect 120895 79337 120977 79360
rect 121063 79337 121129 79360
rect 120743 79318 121129 79337
rect 135863 79423 136249 79442
rect 135863 79400 135929 79423
rect 136015 79400 136097 79423
rect 136183 79400 136249 79423
rect 135863 79360 135872 79400
rect 135912 79360 135929 79400
rect 136015 79360 136036 79400
rect 136076 79360 136097 79400
rect 136183 79360 136200 79400
rect 136240 79360 136249 79400
rect 135863 79337 135929 79360
rect 136015 79337 136097 79360
rect 136183 79337 136249 79360
rect 135863 79318 136249 79337
rect 150983 79423 151369 79442
rect 150983 79400 151049 79423
rect 151135 79400 151217 79423
rect 151303 79400 151369 79423
rect 150983 79360 150992 79400
rect 151032 79360 151049 79400
rect 151135 79360 151156 79400
rect 151196 79360 151217 79400
rect 151303 79360 151320 79400
rect 151360 79360 151369 79400
rect 150983 79337 151049 79360
rect 151135 79337 151217 79360
rect 151303 79337 151369 79360
rect 150983 79318 151369 79337
rect 74143 78667 74529 78686
rect 74143 78644 74209 78667
rect 74295 78644 74377 78667
rect 74463 78644 74529 78667
rect 74143 78604 74152 78644
rect 74192 78604 74209 78644
rect 74295 78604 74316 78644
rect 74356 78604 74377 78644
rect 74463 78604 74480 78644
rect 74520 78604 74529 78644
rect 74143 78581 74209 78604
rect 74295 78581 74377 78604
rect 74463 78581 74529 78604
rect 74143 78562 74529 78581
rect 89263 78667 89649 78686
rect 89263 78644 89329 78667
rect 89415 78644 89497 78667
rect 89583 78644 89649 78667
rect 89263 78604 89272 78644
rect 89312 78604 89329 78644
rect 89415 78604 89436 78644
rect 89476 78604 89497 78644
rect 89583 78604 89600 78644
rect 89640 78604 89649 78644
rect 89263 78581 89329 78604
rect 89415 78581 89497 78604
rect 89583 78581 89649 78604
rect 89263 78562 89649 78581
rect 104383 78667 104769 78686
rect 104383 78644 104449 78667
rect 104535 78644 104617 78667
rect 104703 78644 104769 78667
rect 104383 78604 104392 78644
rect 104432 78604 104449 78644
rect 104535 78604 104556 78644
rect 104596 78604 104617 78644
rect 104703 78604 104720 78644
rect 104760 78604 104769 78644
rect 104383 78581 104449 78604
rect 104535 78581 104617 78604
rect 104703 78581 104769 78604
rect 104383 78562 104769 78581
rect 119503 78667 119889 78686
rect 119503 78644 119569 78667
rect 119655 78644 119737 78667
rect 119823 78644 119889 78667
rect 119503 78604 119512 78644
rect 119552 78604 119569 78644
rect 119655 78604 119676 78644
rect 119716 78604 119737 78644
rect 119823 78604 119840 78644
rect 119880 78604 119889 78644
rect 119503 78581 119569 78604
rect 119655 78581 119737 78604
rect 119823 78581 119889 78604
rect 119503 78562 119889 78581
rect 134623 78667 135009 78686
rect 134623 78644 134689 78667
rect 134775 78644 134857 78667
rect 134943 78644 135009 78667
rect 134623 78604 134632 78644
rect 134672 78604 134689 78644
rect 134775 78604 134796 78644
rect 134836 78604 134857 78644
rect 134943 78604 134960 78644
rect 135000 78604 135009 78644
rect 134623 78581 134689 78604
rect 134775 78581 134857 78604
rect 134943 78581 135009 78604
rect 134623 78562 135009 78581
rect 149743 78667 150129 78686
rect 149743 78644 149809 78667
rect 149895 78644 149977 78667
rect 150063 78644 150129 78667
rect 149743 78604 149752 78644
rect 149792 78604 149809 78644
rect 149895 78604 149916 78644
rect 149956 78604 149977 78644
rect 150063 78604 150080 78644
rect 150120 78604 150129 78644
rect 149743 78581 149809 78604
rect 149895 78581 149977 78604
rect 150063 78581 150129 78604
rect 149743 78562 150129 78581
rect 75383 77911 75769 77930
rect 75383 77888 75449 77911
rect 75535 77888 75617 77911
rect 75703 77888 75769 77911
rect 75383 77848 75392 77888
rect 75432 77848 75449 77888
rect 75535 77848 75556 77888
rect 75596 77848 75617 77888
rect 75703 77848 75720 77888
rect 75760 77848 75769 77888
rect 75383 77825 75449 77848
rect 75535 77825 75617 77848
rect 75703 77825 75769 77848
rect 75383 77806 75769 77825
rect 90503 77911 90889 77930
rect 90503 77888 90569 77911
rect 90655 77888 90737 77911
rect 90823 77888 90889 77911
rect 90503 77848 90512 77888
rect 90552 77848 90569 77888
rect 90655 77848 90676 77888
rect 90716 77848 90737 77888
rect 90823 77848 90840 77888
rect 90880 77848 90889 77888
rect 90503 77825 90569 77848
rect 90655 77825 90737 77848
rect 90823 77825 90889 77848
rect 90503 77806 90889 77825
rect 105623 77911 106009 77930
rect 105623 77888 105689 77911
rect 105775 77888 105857 77911
rect 105943 77888 106009 77911
rect 105623 77848 105632 77888
rect 105672 77848 105689 77888
rect 105775 77848 105796 77888
rect 105836 77848 105857 77888
rect 105943 77848 105960 77888
rect 106000 77848 106009 77888
rect 105623 77825 105689 77848
rect 105775 77825 105857 77848
rect 105943 77825 106009 77848
rect 105623 77806 106009 77825
rect 120743 77911 121129 77930
rect 120743 77888 120809 77911
rect 120895 77888 120977 77911
rect 121063 77888 121129 77911
rect 120743 77848 120752 77888
rect 120792 77848 120809 77888
rect 120895 77848 120916 77888
rect 120956 77848 120977 77888
rect 121063 77848 121080 77888
rect 121120 77848 121129 77888
rect 120743 77825 120809 77848
rect 120895 77825 120977 77848
rect 121063 77825 121129 77848
rect 120743 77806 121129 77825
rect 135863 77911 136249 77930
rect 135863 77888 135929 77911
rect 136015 77888 136097 77911
rect 136183 77888 136249 77911
rect 135863 77848 135872 77888
rect 135912 77848 135929 77888
rect 136015 77848 136036 77888
rect 136076 77848 136097 77888
rect 136183 77848 136200 77888
rect 136240 77848 136249 77888
rect 135863 77825 135929 77848
rect 136015 77825 136097 77848
rect 136183 77825 136249 77848
rect 135863 77806 136249 77825
rect 150983 77911 151369 77930
rect 150983 77888 151049 77911
rect 151135 77888 151217 77911
rect 151303 77888 151369 77911
rect 150983 77848 150992 77888
rect 151032 77848 151049 77888
rect 151135 77848 151156 77888
rect 151196 77848 151217 77888
rect 151303 77848 151320 77888
rect 151360 77848 151369 77888
rect 150983 77825 151049 77848
rect 151135 77825 151217 77848
rect 151303 77825 151369 77848
rect 150983 77806 151369 77825
rect 74143 77155 74529 77174
rect 74143 77132 74209 77155
rect 74295 77132 74377 77155
rect 74463 77132 74529 77155
rect 74143 77092 74152 77132
rect 74192 77092 74209 77132
rect 74295 77092 74316 77132
rect 74356 77092 74377 77132
rect 74463 77092 74480 77132
rect 74520 77092 74529 77132
rect 74143 77069 74209 77092
rect 74295 77069 74377 77092
rect 74463 77069 74529 77092
rect 74143 77050 74529 77069
rect 89263 77155 89649 77174
rect 89263 77132 89329 77155
rect 89415 77132 89497 77155
rect 89583 77132 89649 77155
rect 89263 77092 89272 77132
rect 89312 77092 89329 77132
rect 89415 77092 89436 77132
rect 89476 77092 89497 77132
rect 89583 77092 89600 77132
rect 89640 77092 89649 77132
rect 89263 77069 89329 77092
rect 89415 77069 89497 77092
rect 89583 77069 89649 77092
rect 89263 77050 89649 77069
rect 104383 77155 104769 77174
rect 104383 77132 104449 77155
rect 104535 77132 104617 77155
rect 104703 77132 104769 77155
rect 104383 77092 104392 77132
rect 104432 77092 104449 77132
rect 104535 77092 104556 77132
rect 104596 77092 104617 77132
rect 104703 77092 104720 77132
rect 104760 77092 104769 77132
rect 104383 77069 104449 77092
rect 104535 77069 104617 77092
rect 104703 77069 104769 77092
rect 104383 77050 104769 77069
rect 119503 77155 119889 77174
rect 119503 77132 119569 77155
rect 119655 77132 119737 77155
rect 119823 77132 119889 77155
rect 119503 77092 119512 77132
rect 119552 77092 119569 77132
rect 119655 77092 119676 77132
rect 119716 77092 119737 77132
rect 119823 77092 119840 77132
rect 119880 77092 119889 77132
rect 119503 77069 119569 77092
rect 119655 77069 119737 77092
rect 119823 77069 119889 77092
rect 119503 77050 119889 77069
rect 134623 77155 135009 77174
rect 134623 77132 134689 77155
rect 134775 77132 134857 77155
rect 134943 77132 135009 77155
rect 134623 77092 134632 77132
rect 134672 77092 134689 77132
rect 134775 77092 134796 77132
rect 134836 77092 134857 77132
rect 134943 77092 134960 77132
rect 135000 77092 135009 77132
rect 134623 77069 134689 77092
rect 134775 77069 134857 77092
rect 134943 77069 135009 77092
rect 134623 77050 135009 77069
rect 149743 77155 150129 77174
rect 149743 77132 149809 77155
rect 149895 77132 149977 77155
rect 150063 77132 150129 77155
rect 149743 77092 149752 77132
rect 149792 77092 149809 77132
rect 149895 77092 149916 77132
rect 149956 77092 149977 77132
rect 150063 77092 150080 77132
rect 150120 77092 150129 77132
rect 149743 77069 149809 77092
rect 149895 77069 149977 77092
rect 150063 77069 150129 77092
rect 149743 77050 150129 77069
rect 75383 76399 75769 76418
rect 75383 76376 75449 76399
rect 75535 76376 75617 76399
rect 75703 76376 75769 76399
rect 75383 76336 75392 76376
rect 75432 76336 75449 76376
rect 75535 76336 75556 76376
rect 75596 76336 75617 76376
rect 75703 76336 75720 76376
rect 75760 76336 75769 76376
rect 75383 76313 75449 76336
rect 75535 76313 75617 76336
rect 75703 76313 75769 76336
rect 75383 76294 75769 76313
rect 90503 76399 90889 76418
rect 90503 76376 90569 76399
rect 90655 76376 90737 76399
rect 90823 76376 90889 76399
rect 90503 76336 90512 76376
rect 90552 76336 90569 76376
rect 90655 76336 90676 76376
rect 90716 76336 90737 76376
rect 90823 76336 90840 76376
rect 90880 76336 90889 76376
rect 90503 76313 90569 76336
rect 90655 76313 90737 76336
rect 90823 76313 90889 76336
rect 90503 76294 90889 76313
rect 105623 76399 106009 76418
rect 105623 76376 105689 76399
rect 105775 76376 105857 76399
rect 105943 76376 106009 76399
rect 105623 76336 105632 76376
rect 105672 76336 105689 76376
rect 105775 76336 105796 76376
rect 105836 76336 105857 76376
rect 105943 76336 105960 76376
rect 106000 76336 106009 76376
rect 105623 76313 105689 76336
rect 105775 76313 105857 76336
rect 105943 76313 106009 76336
rect 105623 76294 106009 76313
rect 120743 76399 121129 76418
rect 120743 76376 120809 76399
rect 120895 76376 120977 76399
rect 121063 76376 121129 76399
rect 120743 76336 120752 76376
rect 120792 76336 120809 76376
rect 120895 76336 120916 76376
rect 120956 76336 120977 76376
rect 121063 76336 121080 76376
rect 121120 76336 121129 76376
rect 120743 76313 120809 76336
rect 120895 76313 120977 76336
rect 121063 76313 121129 76336
rect 120743 76294 121129 76313
rect 135863 76399 136249 76418
rect 135863 76376 135929 76399
rect 136015 76376 136097 76399
rect 136183 76376 136249 76399
rect 135863 76336 135872 76376
rect 135912 76336 135929 76376
rect 136015 76336 136036 76376
rect 136076 76336 136097 76376
rect 136183 76336 136200 76376
rect 136240 76336 136249 76376
rect 135863 76313 135929 76336
rect 136015 76313 136097 76336
rect 136183 76313 136249 76336
rect 135863 76294 136249 76313
rect 150983 76399 151369 76418
rect 150983 76376 151049 76399
rect 151135 76376 151217 76399
rect 151303 76376 151369 76399
rect 150983 76336 150992 76376
rect 151032 76336 151049 76376
rect 151135 76336 151156 76376
rect 151196 76336 151217 76376
rect 151303 76336 151320 76376
rect 151360 76336 151369 76376
rect 150983 76313 151049 76336
rect 151135 76313 151217 76336
rect 151303 76313 151369 76336
rect 150983 76294 151369 76313
rect 74143 75643 74529 75662
rect 74143 75620 74209 75643
rect 74295 75620 74377 75643
rect 74463 75620 74529 75643
rect 74143 75580 74152 75620
rect 74192 75580 74209 75620
rect 74295 75580 74316 75620
rect 74356 75580 74377 75620
rect 74463 75580 74480 75620
rect 74520 75580 74529 75620
rect 74143 75557 74209 75580
rect 74295 75557 74377 75580
rect 74463 75557 74529 75580
rect 74143 75538 74529 75557
rect 89263 75643 89649 75662
rect 89263 75620 89329 75643
rect 89415 75620 89497 75643
rect 89583 75620 89649 75643
rect 89263 75580 89272 75620
rect 89312 75580 89329 75620
rect 89415 75580 89436 75620
rect 89476 75580 89497 75620
rect 89583 75580 89600 75620
rect 89640 75580 89649 75620
rect 89263 75557 89329 75580
rect 89415 75557 89497 75580
rect 89583 75557 89649 75580
rect 89263 75538 89649 75557
rect 104383 75643 104769 75662
rect 104383 75620 104449 75643
rect 104535 75620 104617 75643
rect 104703 75620 104769 75643
rect 104383 75580 104392 75620
rect 104432 75580 104449 75620
rect 104535 75580 104556 75620
rect 104596 75580 104617 75620
rect 104703 75580 104720 75620
rect 104760 75580 104769 75620
rect 104383 75557 104449 75580
rect 104535 75557 104617 75580
rect 104703 75557 104769 75580
rect 104383 75538 104769 75557
rect 119503 75643 119889 75662
rect 119503 75620 119569 75643
rect 119655 75620 119737 75643
rect 119823 75620 119889 75643
rect 119503 75580 119512 75620
rect 119552 75580 119569 75620
rect 119655 75580 119676 75620
rect 119716 75580 119737 75620
rect 119823 75580 119840 75620
rect 119880 75580 119889 75620
rect 119503 75557 119569 75580
rect 119655 75557 119737 75580
rect 119823 75557 119889 75580
rect 119503 75538 119889 75557
rect 134623 75643 135009 75662
rect 134623 75620 134689 75643
rect 134775 75620 134857 75643
rect 134943 75620 135009 75643
rect 134623 75580 134632 75620
rect 134672 75580 134689 75620
rect 134775 75580 134796 75620
rect 134836 75580 134857 75620
rect 134943 75580 134960 75620
rect 135000 75580 135009 75620
rect 134623 75557 134689 75580
rect 134775 75557 134857 75580
rect 134943 75557 135009 75580
rect 134623 75538 135009 75557
rect 149743 75643 150129 75662
rect 149743 75620 149809 75643
rect 149895 75620 149977 75643
rect 150063 75620 150129 75643
rect 149743 75580 149752 75620
rect 149792 75580 149809 75620
rect 149895 75580 149916 75620
rect 149956 75580 149977 75620
rect 150063 75580 150080 75620
rect 150120 75580 150129 75620
rect 149743 75557 149809 75580
rect 149895 75557 149977 75580
rect 150063 75557 150129 75580
rect 149743 75538 150129 75557
rect 75383 74887 75769 74906
rect 75383 74864 75449 74887
rect 75535 74864 75617 74887
rect 75703 74864 75769 74887
rect 75383 74824 75392 74864
rect 75432 74824 75449 74864
rect 75535 74824 75556 74864
rect 75596 74824 75617 74864
rect 75703 74824 75720 74864
rect 75760 74824 75769 74864
rect 75383 74801 75449 74824
rect 75535 74801 75617 74824
rect 75703 74801 75769 74824
rect 75383 74782 75769 74801
rect 90503 74887 90889 74906
rect 90503 74864 90569 74887
rect 90655 74864 90737 74887
rect 90823 74864 90889 74887
rect 90503 74824 90512 74864
rect 90552 74824 90569 74864
rect 90655 74824 90676 74864
rect 90716 74824 90737 74864
rect 90823 74824 90840 74864
rect 90880 74824 90889 74864
rect 90503 74801 90569 74824
rect 90655 74801 90737 74824
rect 90823 74801 90889 74824
rect 90503 74782 90889 74801
rect 105623 74887 106009 74906
rect 105623 74864 105689 74887
rect 105775 74864 105857 74887
rect 105943 74864 106009 74887
rect 105623 74824 105632 74864
rect 105672 74824 105689 74864
rect 105775 74824 105796 74864
rect 105836 74824 105857 74864
rect 105943 74824 105960 74864
rect 106000 74824 106009 74864
rect 105623 74801 105689 74824
rect 105775 74801 105857 74824
rect 105943 74801 106009 74824
rect 105623 74782 106009 74801
rect 120743 74887 121129 74906
rect 120743 74864 120809 74887
rect 120895 74864 120977 74887
rect 121063 74864 121129 74887
rect 120743 74824 120752 74864
rect 120792 74824 120809 74864
rect 120895 74824 120916 74864
rect 120956 74824 120977 74864
rect 121063 74824 121080 74864
rect 121120 74824 121129 74864
rect 120743 74801 120809 74824
rect 120895 74801 120977 74824
rect 121063 74801 121129 74824
rect 120743 74782 121129 74801
rect 135863 74887 136249 74906
rect 135863 74864 135929 74887
rect 136015 74864 136097 74887
rect 136183 74864 136249 74887
rect 135863 74824 135872 74864
rect 135912 74824 135929 74864
rect 136015 74824 136036 74864
rect 136076 74824 136097 74864
rect 136183 74824 136200 74864
rect 136240 74824 136249 74864
rect 135863 74801 135929 74824
rect 136015 74801 136097 74824
rect 136183 74801 136249 74824
rect 135863 74782 136249 74801
rect 150983 74887 151369 74906
rect 150983 74864 151049 74887
rect 151135 74864 151217 74887
rect 151303 74864 151369 74887
rect 150983 74824 150992 74864
rect 151032 74824 151049 74864
rect 151135 74824 151156 74864
rect 151196 74824 151217 74864
rect 151303 74824 151320 74864
rect 151360 74824 151369 74864
rect 150983 74801 151049 74824
rect 151135 74801 151217 74824
rect 151303 74801 151369 74824
rect 150983 74782 151369 74801
rect 74143 74131 74529 74150
rect 74143 74108 74209 74131
rect 74295 74108 74377 74131
rect 74463 74108 74529 74131
rect 74143 74068 74152 74108
rect 74192 74068 74209 74108
rect 74295 74068 74316 74108
rect 74356 74068 74377 74108
rect 74463 74068 74480 74108
rect 74520 74068 74529 74108
rect 74143 74045 74209 74068
rect 74295 74045 74377 74068
rect 74463 74045 74529 74068
rect 74143 74026 74529 74045
rect 89263 74131 89649 74150
rect 89263 74108 89329 74131
rect 89415 74108 89497 74131
rect 89583 74108 89649 74131
rect 89263 74068 89272 74108
rect 89312 74068 89329 74108
rect 89415 74068 89436 74108
rect 89476 74068 89497 74108
rect 89583 74068 89600 74108
rect 89640 74068 89649 74108
rect 89263 74045 89329 74068
rect 89415 74045 89497 74068
rect 89583 74045 89649 74068
rect 89263 74026 89649 74045
rect 104383 74131 104769 74150
rect 104383 74108 104449 74131
rect 104535 74108 104617 74131
rect 104703 74108 104769 74131
rect 104383 74068 104392 74108
rect 104432 74068 104449 74108
rect 104535 74068 104556 74108
rect 104596 74068 104617 74108
rect 104703 74068 104720 74108
rect 104760 74068 104769 74108
rect 104383 74045 104449 74068
rect 104535 74045 104617 74068
rect 104703 74045 104769 74068
rect 104383 74026 104769 74045
rect 119503 74131 119889 74150
rect 119503 74108 119569 74131
rect 119655 74108 119737 74131
rect 119823 74108 119889 74131
rect 119503 74068 119512 74108
rect 119552 74068 119569 74108
rect 119655 74068 119676 74108
rect 119716 74068 119737 74108
rect 119823 74068 119840 74108
rect 119880 74068 119889 74108
rect 119503 74045 119569 74068
rect 119655 74045 119737 74068
rect 119823 74045 119889 74068
rect 119503 74026 119889 74045
rect 134623 74131 135009 74150
rect 134623 74108 134689 74131
rect 134775 74108 134857 74131
rect 134943 74108 135009 74131
rect 134623 74068 134632 74108
rect 134672 74068 134689 74108
rect 134775 74068 134796 74108
rect 134836 74068 134857 74108
rect 134943 74068 134960 74108
rect 135000 74068 135009 74108
rect 134623 74045 134689 74068
rect 134775 74045 134857 74068
rect 134943 74045 135009 74068
rect 134623 74026 135009 74045
rect 149743 74131 150129 74150
rect 149743 74108 149809 74131
rect 149895 74108 149977 74131
rect 150063 74108 150129 74131
rect 149743 74068 149752 74108
rect 149792 74068 149809 74108
rect 149895 74068 149916 74108
rect 149956 74068 149977 74108
rect 150063 74068 150080 74108
rect 150120 74068 150129 74108
rect 149743 74045 149809 74068
rect 149895 74045 149977 74068
rect 150063 74045 150129 74068
rect 149743 74026 150129 74045
rect 75383 73375 75769 73394
rect 75383 73352 75449 73375
rect 75535 73352 75617 73375
rect 75703 73352 75769 73375
rect 75383 73312 75392 73352
rect 75432 73312 75449 73352
rect 75535 73312 75556 73352
rect 75596 73312 75617 73352
rect 75703 73312 75720 73352
rect 75760 73312 75769 73352
rect 75383 73289 75449 73312
rect 75535 73289 75617 73312
rect 75703 73289 75769 73312
rect 75383 73270 75769 73289
rect 90503 73375 90889 73394
rect 90503 73352 90569 73375
rect 90655 73352 90737 73375
rect 90823 73352 90889 73375
rect 90503 73312 90512 73352
rect 90552 73312 90569 73352
rect 90655 73312 90676 73352
rect 90716 73312 90737 73352
rect 90823 73312 90840 73352
rect 90880 73312 90889 73352
rect 90503 73289 90569 73312
rect 90655 73289 90737 73312
rect 90823 73289 90889 73312
rect 90503 73270 90889 73289
rect 105623 73375 106009 73394
rect 105623 73352 105689 73375
rect 105775 73352 105857 73375
rect 105943 73352 106009 73375
rect 105623 73312 105632 73352
rect 105672 73312 105689 73352
rect 105775 73312 105796 73352
rect 105836 73312 105857 73352
rect 105943 73312 105960 73352
rect 106000 73312 106009 73352
rect 105623 73289 105689 73312
rect 105775 73289 105857 73312
rect 105943 73289 106009 73312
rect 105623 73270 106009 73289
rect 120743 73375 121129 73394
rect 120743 73352 120809 73375
rect 120895 73352 120977 73375
rect 121063 73352 121129 73375
rect 120743 73312 120752 73352
rect 120792 73312 120809 73352
rect 120895 73312 120916 73352
rect 120956 73312 120977 73352
rect 121063 73312 121080 73352
rect 121120 73312 121129 73352
rect 120743 73289 120809 73312
rect 120895 73289 120977 73312
rect 121063 73289 121129 73312
rect 120743 73270 121129 73289
rect 135863 73375 136249 73394
rect 135863 73352 135929 73375
rect 136015 73352 136097 73375
rect 136183 73352 136249 73375
rect 135863 73312 135872 73352
rect 135912 73312 135929 73352
rect 136015 73312 136036 73352
rect 136076 73312 136097 73352
rect 136183 73312 136200 73352
rect 136240 73312 136249 73352
rect 135863 73289 135929 73312
rect 136015 73289 136097 73312
rect 136183 73289 136249 73312
rect 135863 73270 136249 73289
rect 150983 73375 151369 73394
rect 150983 73352 151049 73375
rect 151135 73352 151217 73375
rect 151303 73352 151369 73375
rect 150983 73312 150992 73352
rect 151032 73312 151049 73352
rect 151135 73312 151156 73352
rect 151196 73312 151217 73352
rect 151303 73312 151320 73352
rect 151360 73312 151369 73352
rect 150983 73289 151049 73312
rect 151135 73289 151217 73312
rect 151303 73289 151369 73312
rect 150983 73270 151369 73289
rect 74143 72619 74529 72638
rect 74143 72596 74209 72619
rect 74295 72596 74377 72619
rect 74463 72596 74529 72619
rect 74143 72556 74152 72596
rect 74192 72556 74209 72596
rect 74295 72556 74316 72596
rect 74356 72556 74377 72596
rect 74463 72556 74480 72596
rect 74520 72556 74529 72596
rect 74143 72533 74209 72556
rect 74295 72533 74377 72556
rect 74463 72533 74529 72556
rect 74143 72514 74529 72533
rect 89263 72619 89649 72638
rect 89263 72596 89329 72619
rect 89415 72596 89497 72619
rect 89583 72596 89649 72619
rect 89263 72556 89272 72596
rect 89312 72556 89329 72596
rect 89415 72556 89436 72596
rect 89476 72556 89497 72596
rect 89583 72556 89600 72596
rect 89640 72556 89649 72596
rect 89263 72533 89329 72556
rect 89415 72533 89497 72556
rect 89583 72533 89649 72556
rect 89263 72514 89649 72533
rect 104383 72619 104769 72638
rect 104383 72596 104449 72619
rect 104535 72596 104617 72619
rect 104703 72596 104769 72619
rect 104383 72556 104392 72596
rect 104432 72556 104449 72596
rect 104535 72556 104556 72596
rect 104596 72556 104617 72596
rect 104703 72556 104720 72596
rect 104760 72556 104769 72596
rect 104383 72533 104449 72556
rect 104535 72533 104617 72556
rect 104703 72533 104769 72556
rect 104383 72514 104769 72533
rect 119503 72619 119889 72638
rect 119503 72596 119569 72619
rect 119655 72596 119737 72619
rect 119823 72596 119889 72619
rect 119503 72556 119512 72596
rect 119552 72556 119569 72596
rect 119655 72556 119676 72596
rect 119716 72556 119737 72596
rect 119823 72556 119840 72596
rect 119880 72556 119889 72596
rect 119503 72533 119569 72556
rect 119655 72533 119737 72556
rect 119823 72533 119889 72556
rect 119503 72514 119889 72533
rect 134623 72619 135009 72638
rect 134623 72596 134689 72619
rect 134775 72596 134857 72619
rect 134943 72596 135009 72619
rect 134623 72556 134632 72596
rect 134672 72556 134689 72596
rect 134775 72556 134796 72596
rect 134836 72556 134857 72596
rect 134943 72556 134960 72596
rect 135000 72556 135009 72596
rect 134623 72533 134689 72556
rect 134775 72533 134857 72556
rect 134943 72533 135009 72556
rect 134623 72514 135009 72533
rect 149743 72619 150129 72638
rect 149743 72596 149809 72619
rect 149895 72596 149977 72619
rect 150063 72596 150129 72619
rect 149743 72556 149752 72596
rect 149792 72556 149809 72596
rect 149895 72556 149916 72596
rect 149956 72556 149977 72596
rect 150063 72556 150080 72596
rect 150120 72556 150129 72596
rect 149743 72533 149809 72556
rect 149895 72533 149977 72556
rect 150063 72533 150129 72556
rect 149743 72514 150129 72533
rect 75383 71863 75769 71882
rect 75383 71840 75449 71863
rect 75535 71840 75617 71863
rect 75703 71840 75769 71863
rect 75383 71800 75392 71840
rect 75432 71800 75449 71840
rect 75535 71800 75556 71840
rect 75596 71800 75617 71840
rect 75703 71800 75720 71840
rect 75760 71800 75769 71840
rect 75383 71777 75449 71800
rect 75535 71777 75617 71800
rect 75703 71777 75769 71800
rect 75383 71758 75769 71777
rect 90503 71863 90889 71882
rect 90503 71840 90569 71863
rect 90655 71840 90737 71863
rect 90823 71840 90889 71863
rect 90503 71800 90512 71840
rect 90552 71800 90569 71840
rect 90655 71800 90676 71840
rect 90716 71800 90737 71840
rect 90823 71800 90840 71840
rect 90880 71800 90889 71840
rect 90503 71777 90569 71800
rect 90655 71777 90737 71800
rect 90823 71777 90889 71800
rect 90503 71758 90889 71777
rect 105623 71863 106009 71882
rect 105623 71840 105689 71863
rect 105775 71840 105857 71863
rect 105943 71840 106009 71863
rect 105623 71800 105632 71840
rect 105672 71800 105689 71840
rect 105775 71800 105796 71840
rect 105836 71800 105857 71840
rect 105943 71800 105960 71840
rect 106000 71800 106009 71840
rect 105623 71777 105689 71800
rect 105775 71777 105857 71800
rect 105943 71777 106009 71800
rect 105623 71758 106009 71777
rect 120743 71863 121129 71882
rect 120743 71840 120809 71863
rect 120895 71840 120977 71863
rect 121063 71840 121129 71863
rect 120743 71800 120752 71840
rect 120792 71800 120809 71840
rect 120895 71800 120916 71840
rect 120956 71800 120977 71840
rect 121063 71800 121080 71840
rect 121120 71800 121129 71840
rect 120743 71777 120809 71800
rect 120895 71777 120977 71800
rect 121063 71777 121129 71800
rect 120743 71758 121129 71777
rect 135863 71863 136249 71882
rect 135863 71840 135929 71863
rect 136015 71840 136097 71863
rect 136183 71840 136249 71863
rect 135863 71800 135872 71840
rect 135912 71800 135929 71840
rect 136015 71800 136036 71840
rect 136076 71800 136097 71840
rect 136183 71800 136200 71840
rect 136240 71800 136249 71840
rect 135863 71777 135929 71800
rect 136015 71777 136097 71800
rect 136183 71777 136249 71800
rect 135863 71758 136249 71777
rect 150983 71863 151369 71882
rect 150983 71840 151049 71863
rect 151135 71840 151217 71863
rect 151303 71840 151369 71863
rect 150983 71800 150992 71840
rect 151032 71800 151049 71840
rect 151135 71800 151156 71840
rect 151196 71800 151217 71840
rect 151303 71800 151320 71840
rect 151360 71800 151369 71840
rect 150983 71777 151049 71800
rect 151135 71777 151217 71800
rect 151303 71777 151369 71800
rect 150983 71758 151369 71777
<< via5 >>
rect 75449 151976 75535 151999
rect 75617 151976 75703 151999
rect 75449 151936 75474 151976
rect 75474 151936 75514 151976
rect 75514 151936 75535 151976
rect 75617 151936 75638 151976
rect 75638 151936 75678 151976
rect 75678 151936 75703 151976
rect 75449 151913 75535 151936
rect 75617 151913 75703 151936
rect 90569 151976 90655 151999
rect 90737 151976 90823 151999
rect 90569 151936 90594 151976
rect 90594 151936 90634 151976
rect 90634 151936 90655 151976
rect 90737 151936 90758 151976
rect 90758 151936 90798 151976
rect 90798 151936 90823 151976
rect 90569 151913 90655 151936
rect 90737 151913 90823 151936
rect 105689 151976 105775 151999
rect 105857 151976 105943 151999
rect 105689 151936 105714 151976
rect 105714 151936 105754 151976
rect 105754 151936 105775 151976
rect 105857 151936 105878 151976
rect 105878 151936 105918 151976
rect 105918 151936 105943 151976
rect 105689 151913 105775 151936
rect 105857 151913 105943 151936
rect 120809 151976 120895 151999
rect 120977 151976 121063 151999
rect 120809 151936 120834 151976
rect 120834 151936 120874 151976
rect 120874 151936 120895 151976
rect 120977 151936 120998 151976
rect 120998 151936 121038 151976
rect 121038 151936 121063 151976
rect 120809 151913 120895 151936
rect 120977 151913 121063 151936
rect 135929 151976 136015 151999
rect 136097 151976 136183 151999
rect 135929 151936 135954 151976
rect 135954 151936 135994 151976
rect 135994 151936 136015 151976
rect 136097 151936 136118 151976
rect 136118 151936 136158 151976
rect 136158 151936 136183 151976
rect 135929 151913 136015 151936
rect 136097 151913 136183 151936
rect 151049 151976 151135 151999
rect 151217 151976 151303 151999
rect 151049 151936 151074 151976
rect 151074 151936 151114 151976
rect 151114 151936 151135 151976
rect 151217 151936 151238 151976
rect 151238 151936 151278 151976
rect 151278 151936 151303 151976
rect 151049 151913 151135 151936
rect 151217 151913 151303 151936
rect 74209 151220 74295 151243
rect 74377 151220 74463 151243
rect 74209 151180 74234 151220
rect 74234 151180 74274 151220
rect 74274 151180 74295 151220
rect 74377 151180 74398 151220
rect 74398 151180 74438 151220
rect 74438 151180 74463 151220
rect 74209 151157 74295 151180
rect 74377 151157 74463 151180
rect 89329 151220 89415 151243
rect 89497 151220 89583 151243
rect 89329 151180 89354 151220
rect 89354 151180 89394 151220
rect 89394 151180 89415 151220
rect 89497 151180 89518 151220
rect 89518 151180 89558 151220
rect 89558 151180 89583 151220
rect 89329 151157 89415 151180
rect 89497 151157 89583 151180
rect 104449 151220 104535 151243
rect 104617 151220 104703 151243
rect 104449 151180 104474 151220
rect 104474 151180 104514 151220
rect 104514 151180 104535 151220
rect 104617 151180 104638 151220
rect 104638 151180 104678 151220
rect 104678 151180 104703 151220
rect 104449 151157 104535 151180
rect 104617 151157 104703 151180
rect 119569 151220 119655 151243
rect 119737 151220 119823 151243
rect 119569 151180 119594 151220
rect 119594 151180 119634 151220
rect 119634 151180 119655 151220
rect 119737 151180 119758 151220
rect 119758 151180 119798 151220
rect 119798 151180 119823 151220
rect 119569 151157 119655 151180
rect 119737 151157 119823 151180
rect 134689 151220 134775 151243
rect 134857 151220 134943 151243
rect 134689 151180 134714 151220
rect 134714 151180 134754 151220
rect 134754 151180 134775 151220
rect 134857 151180 134878 151220
rect 134878 151180 134918 151220
rect 134918 151180 134943 151220
rect 134689 151157 134775 151180
rect 134857 151157 134943 151180
rect 149809 151220 149895 151243
rect 149977 151220 150063 151243
rect 149809 151180 149834 151220
rect 149834 151180 149874 151220
rect 149874 151180 149895 151220
rect 149977 151180 149998 151220
rect 149998 151180 150038 151220
rect 150038 151180 150063 151220
rect 149809 151157 149895 151180
rect 149977 151157 150063 151180
rect 75449 150464 75535 150487
rect 75617 150464 75703 150487
rect 75449 150424 75474 150464
rect 75474 150424 75514 150464
rect 75514 150424 75535 150464
rect 75617 150424 75638 150464
rect 75638 150424 75678 150464
rect 75678 150424 75703 150464
rect 75449 150401 75535 150424
rect 75617 150401 75703 150424
rect 90569 150464 90655 150487
rect 90737 150464 90823 150487
rect 90569 150424 90594 150464
rect 90594 150424 90634 150464
rect 90634 150424 90655 150464
rect 90737 150424 90758 150464
rect 90758 150424 90798 150464
rect 90798 150424 90823 150464
rect 90569 150401 90655 150424
rect 90737 150401 90823 150424
rect 105689 150464 105775 150487
rect 105857 150464 105943 150487
rect 105689 150424 105714 150464
rect 105714 150424 105754 150464
rect 105754 150424 105775 150464
rect 105857 150424 105878 150464
rect 105878 150424 105918 150464
rect 105918 150424 105943 150464
rect 105689 150401 105775 150424
rect 105857 150401 105943 150424
rect 120809 150464 120895 150487
rect 120977 150464 121063 150487
rect 120809 150424 120834 150464
rect 120834 150424 120874 150464
rect 120874 150424 120895 150464
rect 120977 150424 120998 150464
rect 120998 150424 121038 150464
rect 121038 150424 121063 150464
rect 120809 150401 120895 150424
rect 120977 150401 121063 150424
rect 135929 150464 136015 150487
rect 136097 150464 136183 150487
rect 135929 150424 135954 150464
rect 135954 150424 135994 150464
rect 135994 150424 136015 150464
rect 136097 150424 136118 150464
rect 136118 150424 136158 150464
rect 136158 150424 136183 150464
rect 135929 150401 136015 150424
rect 136097 150401 136183 150424
rect 151049 150464 151135 150487
rect 151217 150464 151303 150487
rect 151049 150424 151074 150464
rect 151074 150424 151114 150464
rect 151114 150424 151135 150464
rect 151217 150424 151238 150464
rect 151238 150424 151278 150464
rect 151278 150424 151303 150464
rect 151049 150401 151135 150424
rect 151217 150401 151303 150424
rect 74209 149708 74295 149731
rect 74377 149708 74463 149731
rect 74209 149668 74234 149708
rect 74234 149668 74274 149708
rect 74274 149668 74295 149708
rect 74377 149668 74398 149708
rect 74398 149668 74438 149708
rect 74438 149668 74463 149708
rect 74209 149645 74295 149668
rect 74377 149645 74463 149668
rect 89329 149708 89415 149731
rect 89497 149708 89583 149731
rect 89329 149668 89354 149708
rect 89354 149668 89394 149708
rect 89394 149668 89415 149708
rect 89497 149668 89518 149708
rect 89518 149668 89558 149708
rect 89558 149668 89583 149708
rect 89329 149645 89415 149668
rect 89497 149645 89583 149668
rect 104449 149708 104535 149731
rect 104617 149708 104703 149731
rect 104449 149668 104474 149708
rect 104474 149668 104514 149708
rect 104514 149668 104535 149708
rect 104617 149668 104638 149708
rect 104638 149668 104678 149708
rect 104678 149668 104703 149708
rect 104449 149645 104535 149668
rect 104617 149645 104703 149668
rect 119569 149708 119655 149731
rect 119737 149708 119823 149731
rect 119569 149668 119594 149708
rect 119594 149668 119634 149708
rect 119634 149668 119655 149708
rect 119737 149668 119758 149708
rect 119758 149668 119798 149708
rect 119798 149668 119823 149708
rect 119569 149645 119655 149668
rect 119737 149645 119823 149668
rect 134689 149708 134775 149731
rect 134857 149708 134943 149731
rect 134689 149668 134714 149708
rect 134714 149668 134754 149708
rect 134754 149668 134775 149708
rect 134857 149668 134878 149708
rect 134878 149668 134918 149708
rect 134918 149668 134943 149708
rect 134689 149645 134775 149668
rect 134857 149645 134943 149668
rect 149809 149708 149895 149731
rect 149977 149708 150063 149731
rect 149809 149668 149834 149708
rect 149834 149668 149874 149708
rect 149874 149668 149895 149708
rect 149977 149668 149998 149708
rect 149998 149668 150038 149708
rect 150038 149668 150063 149708
rect 149809 149645 149895 149668
rect 149977 149645 150063 149668
rect 75449 148952 75535 148975
rect 75617 148952 75703 148975
rect 75449 148912 75474 148952
rect 75474 148912 75514 148952
rect 75514 148912 75535 148952
rect 75617 148912 75638 148952
rect 75638 148912 75678 148952
rect 75678 148912 75703 148952
rect 75449 148889 75535 148912
rect 75617 148889 75703 148912
rect 90569 148952 90655 148975
rect 90737 148952 90823 148975
rect 90569 148912 90594 148952
rect 90594 148912 90634 148952
rect 90634 148912 90655 148952
rect 90737 148912 90758 148952
rect 90758 148912 90798 148952
rect 90798 148912 90823 148952
rect 90569 148889 90655 148912
rect 90737 148889 90823 148912
rect 105689 148952 105775 148975
rect 105857 148952 105943 148975
rect 105689 148912 105714 148952
rect 105714 148912 105754 148952
rect 105754 148912 105775 148952
rect 105857 148912 105878 148952
rect 105878 148912 105918 148952
rect 105918 148912 105943 148952
rect 105689 148889 105775 148912
rect 105857 148889 105943 148912
rect 120809 148952 120895 148975
rect 120977 148952 121063 148975
rect 120809 148912 120834 148952
rect 120834 148912 120874 148952
rect 120874 148912 120895 148952
rect 120977 148912 120998 148952
rect 120998 148912 121038 148952
rect 121038 148912 121063 148952
rect 120809 148889 120895 148912
rect 120977 148889 121063 148912
rect 135929 148952 136015 148975
rect 136097 148952 136183 148975
rect 135929 148912 135954 148952
rect 135954 148912 135994 148952
rect 135994 148912 136015 148952
rect 136097 148912 136118 148952
rect 136118 148912 136158 148952
rect 136158 148912 136183 148952
rect 135929 148889 136015 148912
rect 136097 148889 136183 148912
rect 151049 148952 151135 148975
rect 151217 148952 151303 148975
rect 151049 148912 151074 148952
rect 151074 148912 151114 148952
rect 151114 148912 151135 148952
rect 151217 148912 151238 148952
rect 151238 148912 151278 148952
rect 151278 148912 151303 148952
rect 151049 148889 151135 148912
rect 151217 148889 151303 148912
rect 74209 148196 74295 148219
rect 74377 148196 74463 148219
rect 74209 148156 74234 148196
rect 74234 148156 74274 148196
rect 74274 148156 74295 148196
rect 74377 148156 74398 148196
rect 74398 148156 74438 148196
rect 74438 148156 74463 148196
rect 74209 148133 74295 148156
rect 74377 148133 74463 148156
rect 89329 148196 89415 148219
rect 89497 148196 89583 148219
rect 89329 148156 89354 148196
rect 89354 148156 89394 148196
rect 89394 148156 89415 148196
rect 89497 148156 89518 148196
rect 89518 148156 89558 148196
rect 89558 148156 89583 148196
rect 89329 148133 89415 148156
rect 89497 148133 89583 148156
rect 104449 148196 104535 148219
rect 104617 148196 104703 148219
rect 104449 148156 104474 148196
rect 104474 148156 104514 148196
rect 104514 148156 104535 148196
rect 104617 148156 104638 148196
rect 104638 148156 104678 148196
rect 104678 148156 104703 148196
rect 104449 148133 104535 148156
rect 104617 148133 104703 148156
rect 119569 148196 119655 148219
rect 119737 148196 119823 148219
rect 119569 148156 119594 148196
rect 119594 148156 119634 148196
rect 119634 148156 119655 148196
rect 119737 148156 119758 148196
rect 119758 148156 119798 148196
rect 119798 148156 119823 148196
rect 119569 148133 119655 148156
rect 119737 148133 119823 148156
rect 134689 148196 134775 148219
rect 134857 148196 134943 148219
rect 134689 148156 134714 148196
rect 134714 148156 134754 148196
rect 134754 148156 134775 148196
rect 134857 148156 134878 148196
rect 134878 148156 134918 148196
rect 134918 148156 134943 148196
rect 134689 148133 134775 148156
rect 134857 148133 134943 148156
rect 149809 148196 149895 148219
rect 149977 148196 150063 148219
rect 149809 148156 149834 148196
rect 149834 148156 149874 148196
rect 149874 148156 149895 148196
rect 149977 148156 149998 148196
rect 149998 148156 150038 148196
rect 150038 148156 150063 148196
rect 149809 148133 149895 148156
rect 149977 148133 150063 148156
rect 75449 147440 75535 147463
rect 75617 147440 75703 147463
rect 75449 147400 75474 147440
rect 75474 147400 75514 147440
rect 75514 147400 75535 147440
rect 75617 147400 75638 147440
rect 75638 147400 75678 147440
rect 75678 147400 75703 147440
rect 75449 147377 75535 147400
rect 75617 147377 75703 147400
rect 90569 147440 90655 147463
rect 90737 147440 90823 147463
rect 90569 147400 90594 147440
rect 90594 147400 90634 147440
rect 90634 147400 90655 147440
rect 90737 147400 90758 147440
rect 90758 147400 90798 147440
rect 90798 147400 90823 147440
rect 90569 147377 90655 147400
rect 90737 147377 90823 147400
rect 105689 147440 105775 147463
rect 105857 147440 105943 147463
rect 105689 147400 105714 147440
rect 105714 147400 105754 147440
rect 105754 147400 105775 147440
rect 105857 147400 105878 147440
rect 105878 147400 105918 147440
rect 105918 147400 105943 147440
rect 105689 147377 105775 147400
rect 105857 147377 105943 147400
rect 120809 147440 120895 147463
rect 120977 147440 121063 147463
rect 120809 147400 120834 147440
rect 120834 147400 120874 147440
rect 120874 147400 120895 147440
rect 120977 147400 120998 147440
rect 120998 147400 121038 147440
rect 121038 147400 121063 147440
rect 120809 147377 120895 147400
rect 120977 147377 121063 147400
rect 135929 147440 136015 147463
rect 136097 147440 136183 147463
rect 135929 147400 135954 147440
rect 135954 147400 135994 147440
rect 135994 147400 136015 147440
rect 136097 147400 136118 147440
rect 136118 147400 136158 147440
rect 136158 147400 136183 147440
rect 135929 147377 136015 147400
rect 136097 147377 136183 147400
rect 151049 147440 151135 147463
rect 151217 147440 151303 147463
rect 151049 147400 151074 147440
rect 151074 147400 151114 147440
rect 151114 147400 151135 147440
rect 151217 147400 151238 147440
rect 151238 147400 151278 147440
rect 151278 147400 151303 147440
rect 151049 147377 151135 147400
rect 151217 147377 151303 147400
rect 74209 146684 74295 146707
rect 74377 146684 74463 146707
rect 74209 146644 74234 146684
rect 74234 146644 74274 146684
rect 74274 146644 74295 146684
rect 74377 146644 74398 146684
rect 74398 146644 74438 146684
rect 74438 146644 74463 146684
rect 74209 146621 74295 146644
rect 74377 146621 74463 146644
rect 89329 146684 89415 146707
rect 89497 146684 89583 146707
rect 89329 146644 89354 146684
rect 89354 146644 89394 146684
rect 89394 146644 89415 146684
rect 89497 146644 89518 146684
rect 89518 146644 89558 146684
rect 89558 146644 89583 146684
rect 89329 146621 89415 146644
rect 89497 146621 89583 146644
rect 104449 146684 104535 146707
rect 104617 146684 104703 146707
rect 104449 146644 104474 146684
rect 104474 146644 104514 146684
rect 104514 146644 104535 146684
rect 104617 146644 104638 146684
rect 104638 146644 104678 146684
rect 104678 146644 104703 146684
rect 104449 146621 104535 146644
rect 104617 146621 104703 146644
rect 119569 146684 119655 146707
rect 119737 146684 119823 146707
rect 119569 146644 119594 146684
rect 119594 146644 119634 146684
rect 119634 146644 119655 146684
rect 119737 146644 119758 146684
rect 119758 146644 119798 146684
rect 119798 146644 119823 146684
rect 119569 146621 119655 146644
rect 119737 146621 119823 146644
rect 134689 146684 134775 146707
rect 134857 146684 134943 146707
rect 134689 146644 134714 146684
rect 134714 146644 134754 146684
rect 134754 146644 134775 146684
rect 134857 146644 134878 146684
rect 134878 146644 134918 146684
rect 134918 146644 134943 146684
rect 134689 146621 134775 146644
rect 134857 146621 134943 146644
rect 149809 146684 149895 146707
rect 149977 146684 150063 146707
rect 149809 146644 149834 146684
rect 149834 146644 149874 146684
rect 149874 146644 149895 146684
rect 149977 146644 149998 146684
rect 149998 146644 150038 146684
rect 150038 146644 150063 146684
rect 149809 146621 149895 146644
rect 149977 146621 150063 146644
rect 75449 145928 75535 145951
rect 75617 145928 75703 145951
rect 75449 145888 75474 145928
rect 75474 145888 75514 145928
rect 75514 145888 75535 145928
rect 75617 145888 75638 145928
rect 75638 145888 75678 145928
rect 75678 145888 75703 145928
rect 75449 145865 75535 145888
rect 75617 145865 75703 145888
rect 90569 145928 90655 145951
rect 90737 145928 90823 145951
rect 90569 145888 90594 145928
rect 90594 145888 90634 145928
rect 90634 145888 90655 145928
rect 90737 145888 90758 145928
rect 90758 145888 90798 145928
rect 90798 145888 90823 145928
rect 90569 145865 90655 145888
rect 90737 145865 90823 145888
rect 105689 145928 105775 145951
rect 105857 145928 105943 145951
rect 105689 145888 105714 145928
rect 105714 145888 105754 145928
rect 105754 145888 105775 145928
rect 105857 145888 105878 145928
rect 105878 145888 105918 145928
rect 105918 145888 105943 145928
rect 105689 145865 105775 145888
rect 105857 145865 105943 145888
rect 120809 145928 120895 145951
rect 120977 145928 121063 145951
rect 120809 145888 120834 145928
rect 120834 145888 120874 145928
rect 120874 145888 120895 145928
rect 120977 145888 120998 145928
rect 120998 145888 121038 145928
rect 121038 145888 121063 145928
rect 120809 145865 120895 145888
rect 120977 145865 121063 145888
rect 135929 145928 136015 145951
rect 136097 145928 136183 145951
rect 135929 145888 135954 145928
rect 135954 145888 135994 145928
rect 135994 145888 136015 145928
rect 136097 145888 136118 145928
rect 136118 145888 136158 145928
rect 136158 145888 136183 145928
rect 135929 145865 136015 145888
rect 136097 145865 136183 145888
rect 151049 145928 151135 145951
rect 151217 145928 151303 145951
rect 151049 145888 151074 145928
rect 151074 145888 151114 145928
rect 151114 145888 151135 145928
rect 151217 145888 151238 145928
rect 151238 145888 151278 145928
rect 151278 145888 151303 145928
rect 151049 145865 151135 145888
rect 151217 145865 151303 145888
rect 74209 145172 74295 145195
rect 74377 145172 74463 145195
rect 74209 145132 74234 145172
rect 74234 145132 74274 145172
rect 74274 145132 74295 145172
rect 74377 145132 74398 145172
rect 74398 145132 74438 145172
rect 74438 145132 74463 145172
rect 74209 145109 74295 145132
rect 74377 145109 74463 145132
rect 89329 145172 89415 145195
rect 89497 145172 89583 145195
rect 89329 145132 89354 145172
rect 89354 145132 89394 145172
rect 89394 145132 89415 145172
rect 89497 145132 89518 145172
rect 89518 145132 89558 145172
rect 89558 145132 89583 145172
rect 89329 145109 89415 145132
rect 89497 145109 89583 145132
rect 104449 145172 104535 145195
rect 104617 145172 104703 145195
rect 104449 145132 104474 145172
rect 104474 145132 104514 145172
rect 104514 145132 104535 145172
rect 104617 145132 104638 145172
rect 104638 145132 104678 145172
rect 104678 145132 104703 145172
rect 104449 145109 104535 145132
rect 104617 145109 104703 145132
rect 119569 145172 119655 145195
rect 119737 145172 119823 145195
rect 119569 145132 119594 145172
rect 119594 145132 119634 145172
rect 119634 145132 119655 145172
rect 119737 145132 119758 145172
rect 119758 145132 119798 145172
rect 119798 145132 119823 145172
rect 119569 145109 119655 145132
rect 119737 145109 119823 145132
rect 134689 145172 134775 145195
rect 134857 145172 134943 145195
rect 134689 145132 134714 145172
rect 134714 145132 134754 145172
rect 134754 145132 134775 145172
rect 134857 145132 134878 145172
rect 134878 145132 134918 145172
rect 134918 145132 134943 145172
rect 134689 145109 134775 145132
rect 134857 145109 134943 145132
rect 149809 145172 149895 145195
rect 149977 145172 150063 145195
rect 149809 145132 149834 145172
rect 149834 145132 149874 145172
rect 149874 145132 149895 145172
rect 149977 145132 149998 145172
rect 149998 145132 150038 145172
rect 150038 145132 150063 145172
rect 149809 145109 149895 145132
rect 149977 145109 150063 145132
rect 75449 144416 75535 144439
rect 75617 144416 75703 144439
rect 75449 144376 75474 144416
rect 75474 144376 75514 144416
rect 75514 144376 75535 144416
rect 75617 144376 75638 144416
rect 75638 144376 75678 144416
rect 75678 144376 75703 144416
rect 75449 144353 75535 144376
rect 75617 144353 75703 144376
rect 90569 144416 90655 144439
rect 90737 144416 90823 144439
rect 90569 144376 90594 144416
rect 90594 144376 90634 144416
rect 90634 144376 90655 144416
rect 90737 144376 90758 144416
rect 90758 144376 90798 144416
rect 90798 144376 90823 144416
rect 90569 144353 90655 144376
rect 90737 144353 90823 144376
rect 105689 144416 105775 144439
rect 105857 144416 105943 144439
rect 105689 144376 105714 144416
rect 105714 144376 105754 144416
rect 105754 144376 105775 144416
rect 105857 144376 105878 144416
rect 105878 144376 105918 144416
rect 105918 144376 105943 144416
rect 105689 144353 105775 144376
rect 105857 144353 105943 144376
rect 120809 144416 120895 144439
rect 120977 144416 121063 144439
rect 120809 144376 120834 144416
rect 120834 144376 120874 144416
rect 120874 144376 120895 144416
rect 120977 144376 120998 144416
rect 120998 144376 121038 144416
rect 121038 144376 121063 144416
rect 120809 144353 120895 144376
rect 120977 144353 121063 144376
rect 135929 144416 136015 144439
rect 136097 144416 136183 144439
rect 135929 144376 135954 144416
rect 135954 144376 135994 144416
rect 135994 144376 136015 144416
rect 136097 144376 136118 144416
rect 136118 144376 136158 144416
rect 136158 144376 136183 144416
rect 135929 144353 136015 144376
rect 136097 144353 136183 144376
rect 151049 144416 151135 144439
rect 151217 144416 151303 144439
rect 151049 144376 151074 144416
rect 151074 144376 151114 144416
rect 151114 144376 151135 144416
rect 151217 144376 151238 144416
rect 151238 144376 151278 144416
rect 151278 144376 151303 144416
rect 151049 144353 151135 144376
rect 151217 144353 151303 144376
rect 74209 143660 74295 143683
rect 74377 143660 74463 143683
rect 74209 143620 74234 143660
rect 74234 143620 74274 143660
rect 74274 143620 74295 143660
rect 74377 143620 74398 143660
rect 74398 143620 74438 143660
rect 74438 143620 74463 143660
rect 74209 143597 74295 143620
rect 74377 143597 74463 143620
rect 89329 143660 89415 143683
rect 89497 143660 89583 143683
rect 89329 143620 89354 143660
rect 89354 143620 89394 143660
rect 89394 143620 89415 143660
rect 89497 143620 89518 143660
rect 89518 143620 89558 143660
rect 89558 143620 89583 143660
rect 89329 143597 89415 143620
rect 89497 143597 89583 143620
rect 104449 143660 104535 143683
rect 104617 143660 104703 143683
rect 104449 143620 104474 143660
rect 104474 143620 104514 143660
rect 104514 143620 104535 143660
rect 104617 143620 104638 143660
rect 104638 143620 104678 143660
rect 104678 143620 104703 143660
rect 104449 143597 104535 143620
rect 104617 143597 104703 143620
rect 119569 143660 119655 143683
rect 119737 143660 119823 143683
rect 119569 143620 119594 143660
rect 119594 143620 119634 143660
rect 119634 143620 119655 143660
rect 119737 143620 119758 143660
rect 119758 143620 119798 143660
rect 119798 143620 119823 143660
rect 119569 143597 119655 143620
rect 119737 143597 119823 143620
rect 134689 143660 134775 143683
rect 134857 143660 134943 143683
rect 134689 143620 134714 143660
rect 134714 143620 134754 143660
rect 134754 143620 134775 143660
rect 134857 143620 134878 143660
rect 134878 143620 134918 143660
rect 134918 143620 134943 143660
rect 134689 143597 134775 143620
rect 134857 143597 134943 143620
rect 149809 143660 149895 143683
rect 149977 143660 150063 143683
rect 149809 143620 149834 143660
rect 149834 143620 149874 143660
rect 149874 143620 149895 143660
rect 149977 143620 149998 143660
rect 149998 143620 150038 143660
rect 150038 143620 150063 143660
rect 149809 143597 149895 143620
rect 149977 143597 150063 143620
rect 75449 142904 75535 142927
rect 75617 142904 75703 142927
rect 75449 142864 75474 142904
rect 75474 142864 75514 142904
rect 75514 142864 75535 142904
rect 75617 142864 75638 142904
rect 75638 142864 75678 142904
rect 75678 142864 75703 142904
rect 75449 142841 75535 142864
rect 75617 142841 75703 142864
rect 90569 142904 90655 142927
rect 90737 142904 90823 142927
rect 90569 142864 90594 142904
rect 90594 142864 90634 142904
rect 90634 142864 90655 142904
rect 90737 142864 90758 142904
rect 90758 142864 90798 142904
rect 90798 142864 90823 142904
rect 90569 142841 90655 142864
rect 90737 142841 90823 142864
rect 105689 142904 105775 142927
rect 105857 142904 105943 142927
rect 105689 142864 105714 142904
rect 105714 142864 105754 142904
rect 105754 142864 105775 142904
rect 105857 142864 105878 142904
rect 105878 142864 105918 142904
rect 105918 142864 105943 142904
rect 105689 142841 105775 142864
rect 105857 142841 105943 142864
rect 120809 142904 120895 142927
rect 120977 142904 121063 142927
rect 120809 142864 120834 142904
rect 120834 142864 120874 142904
rect 120874 142864 120895 142904
rect 120977 142864 120998 142904
rect 120998 142864 121038 142904
rect 121038 142864 121063 142904
rect 120809 142841 120895 142864
rect 120977 142841 121063 142864
rect 135929 142904 136015 142927
rect 136097 142904 136183 142927
rect 135929 142864 135954 142904
rect 135954 142864 135994 142904
rect 135994 142864 136015 142904
rect 136097 142864 136118 142904
rect 136118 142864 136158 142904
rect 136158 142864 136183 142904
rect 135929 142841 136015 142864
rect 136097 142841 136183 142864
rect 151049 142904 151135 142927
rect 151217 142904 151303 142927
rect 151049 142864 151074 142904
rect 151074 142864 151114 142904
rect 151114 142864 151135 142904
rect 151217 142864 151238 142904
rect 151238 142864 151278 142904
rect 151278 142864 151303 142904
rect 151049 142841 151135 142864
rect 151217 142841 151303 142864
rect 74209 142148 74295 142171
rect 74377 142148 74463 142171
rect 74209 142108 74234 142148
rect 74234 142108 74274 142148
rect 74274 142108 74295 142148
rect 74377 142108 74398 142148
rect 74398 142108 74438 142148
rect 74438 142108 74463 142148
rect 74209 142085 74295 142108
rect 74377 142085 74463 142108
rect 89329 142148 89415 142171
rect 89497 142148 89583 142171
rect 89329 142108 89354 142148
rect 89354 142108 89394 142148
rect 89394 142108 89415 142148
rect 89497 142108 89518 142148
rect 89518 142108 89558 142148
rect 89558 142108 89583 142148
rect 89329 142085 89415 142108
rect 89497 142085 89583 142108
rect 104449 142148 104535 142171
rect 104617 142148 104703 142171
rect 104449 142108 104474 142148
rect 104474 142108 104514 142148
rect 104514 142108 104535 142148
rect 104617 142108 104638 142148
rect 104638 142108 104678 142148
rect 104678 142108 104703 142148
rect 104449 142085 104535 142108
rect 104617 142085 104703 142108
rect 119569 142148 119655 142171
rect 119737 142148 119823 142171
rect 119569 142108 119594 142148
rect 119594 142108 119634 142148
rect 119634 142108 119655 142148
rect 119737 142108 119758 142148
rect 119758 142108 119798 142148
rect 119798 142108 119823 142148
rect 119569 142085 119655 142108
rect 119737 142085 119823 142108
rect 134689 142148 134775 142171
rect 134857 142148 134943 142171
rect 134689 142108 134714 142148
rect 134714 142108 134754 142148
rect 134754 142108 134775 142148
rect 134857 142108 134878 142148
rect 134878 142108 134918 142148
rect 134918 142108 134943 142148
rect 134689 142085 134775 142108
rect 134857 142085 134943 142108
rect 149809 142148 149895 142171
rect 149977 142148 150063 142171
rect 149809 142108 149834 142148
rect 149834 142108 149874 142148
rect 149874 142108 149895 142148
rect 149977 142108 149998 142148
rect 149998 142108 150038 142148
rect 150038 142108 150063 142148
rect 149809 142085 149895 142108
rect 149977 142085 150063 142108
rect 75449 141392 75535 141415
rect 75617 141392 75703 141415
rect 75449 141352 75474 141392
rect 75474 141352 75514 141392
rect 75514 141352 75535 141392
rect 75617 141352 75638 141392
rect 75638 141352 75678 141392
rect 75678 141352 75703 141392
rect 75449 141329 75535 141352
rect 75617 141329 75703 141352
rect 90569 141392 90655 141415
rect 90737 141392 90823 141415
rect 90569 141352 90594 141392
rect 90594 141352 90634 141392
rect 90634 141352 90655 141392
rect 90737 141352 90758 141392
rect 90758 141352 90798 141392
rect 90798 141352 90823 141392
rect 90569 141329 90655 141352
rect 90737 141329 90823 141352
rect 105689 141392 105775 141415
rect 105857 141392 105943 141415
rect 105689 141352 105714 141392
rect 105714 141352 105754 141392
rect 105754 141352 105775 141392
rect 105857 141352 105878 141392
rect 105878 141352 105918 141392
rect 105918 141352 105943 141392
rect 105689 141329 105775 141352
rect 105857 141329 105943 141352
rect 120809 141392 120895 141415
rect 120977 141392 121063 141415
rect 120809 141352 120834 141392
rect 120834 141352 120874 141392
rect 120874 141352 120895 141392
rect 120977 141352 120998 141392
rect 120998 141352 121038 141392
rect 121038 141352 121063 141392
rect 120809 141329 120895 141352
rect 120977 141329 121063 141352
rect 135929 141392 136015 141415
rect 136097 141392 136183 141415
rect 135929 141352 135954 141392
rect 135954 141352 135994 141392
rect 135994 141352 136015 141392
rect 136097 141352 136118 141392
rect 136118 141352 136158 141392
rect 136158 141352 136183 141392
rect 135929 141329 136015 141352
rect 136097 141329 136183 141352
rect 151049 141392 151135 141415
rect 151217 141392 151303 141415
rect 151049 141352 151074 141392
rect 151074 141352 151114 141392
rect 151114 141352 151135 141392
rect 151217 141352 151238 141392
rect 151238 141352 151278 141392
rect 151278 141352 151303 141392
rect 151049 141329 151135 141352
rect 151217 141329 151303 141352
rect 74209 140636 74295 140659
rect 74377 140636 74463 140659
rect 74209 140596 74234 140636
rect 74234 140596 74274 140636
rect 74274 140596 74295 140636
rect 74377 140596 74398 140636
rect 74398 140596 74438 140636
rect 74438 140596 74463 140636
rect 74209 140573 74295 140596
rect 74377 140573 74463 140596
rect 89329 140636 89415 140659
rect 89497 140636 89583 140659
rect 89329 140596 89354 140636
rect 89354 140596 89394 140636
rect 89394 140596 89415 140636
rect 89497 140596 89518 140636
rect 89518 140596 89558 140636
rect 89558 140596 89583 140636
rect 89329 140573 89415 140596
rect 89497 140573 89583 140596
rect 104449 140636 104535 140659
rect 104617 140636 104703 140659
rect 104449 140596 104474 140636
rect 104474 140596 104514 140636
rect 104514 140596 104535 140636
rect 104617 140596 104638 140636
rect 104638 140596 104678 140636
rect 104678 140596 104703 140636
rect 104449 140573 104535 140596
rect 104617 140573 104703 140596
rect 119569 140636 119655 140659
rect 119737 140636 119823 140659
rect 119569 140596 119594 140636
rect 119594 140596 119634 140636
rect 119634 140596 119655 140636
rect 119737 140596 119758 140636
rect 119758 140596 119798 140636
rect 119798 140596 119823 140636
rect 119569 140573 119655 140596
rect 119737 140573 119823 140596
rect 134689 140636 134775 140659
rect 134857 140636 134943 140659
rect 134689 140596 134714 140636
rect 134714 140596 134754 140636
rect 134754 140596 134775 140636
rect 134857 140596 134878 140636
rect 134878 140596 134918 140636
rect 134918 140596 134943 140636
rect 134689 140573 134775 140596
rect 134857 140573 134943 140596
rect 149809 140636 149895 140659
rect 149977 140636 150063 140659
rect 149809 140596 149834 140636
rect 149834 140596 149874 140636
rect 149874 140596 149895 140636
rect 149977 140596 149998 140636
rect 149998 140596 150038 140636
rect 150038 140596 150063 140636
rect 149809 140573 149895 140596
rect 149977 140573 150063 140596
rect 75449 139880 75535 139903
rect 75617 139880 75703 139903
rect 75449 139840 75474 139880
rect 75474 139840 75514 139880
rect 75514 139840 75535 139880
rect 75617 139840 75638 139880
rect 75638 139840 75678 139880
rect 75678 139840 75703 139880
rect 75449 139817 75535 139840
rect 75617 139817 75703 139840
rect 90569 139880 90655 139903
rect 90737 139880 90823 139903
rect 90569 139840 90594 139880
rect 90594 139840 90634 139880
rect 90634 139840 90655 139880
rect 90737 139840 90758 139880
rect 90758 139840 90798 139880
rect 90798 139840 90823 139880
rect 90569 139817 90655 139840
rect 90737 139817 90823 139840
rect 105689 139880 105775 139903
rect 105857 139880 105943 139903
rect 105689 139840 105714 139880
rect 105714 139840 105754 139880
rect 105754 139840 105775 139880
rect 105857 139840 105878 139880
rect 105878 139840 105918 139880
rect 105918 139840 105943 139880
rect 105689 139817 105775 139840
rect 105857 139817 105943 139840
rect 120809 139880 120895 139903
rect 120977 139880 121063 139903
rect 120809 139840 120834 139880
rect 120834 139840 120874 139880
rect 120874 139840 120895 139880
rect 120977 139840 120998 139880
rect 120998 139840 121038 139880
rect 121038 139840 121063 139880
rect 120809 139817 120895 139840
rect 120977 139817 121063 139840
rect 135929 139880 136015 139903
rect 136097 139880 136183 139903
rect 135929 139840 135954 139880
rect 135954 139840 135994 139880
rect 135994 139840 136015 139880
rect 136097 139840 136118 139880
rect 136118 139840 136158 139880
rect 136158 139840 136183 139880
rect 135929 139817 136015 139840
rect 136097 139817 136183 139840
rect 151049 139880 151135 139903
rect 151217 139880 151303 139903
rect 151049 139840 151074 139880
rect 151074 139840 151114 139880
rect 151114 139840 151135 139880
rect 151217 139840 151238 139880
rect 151238 139840 151278 139880
rect 151278 139840 151303 139880
rect 151049 139817 151135 139840
rect 151217 139817 151303 139840
rect 74209 139124 74295 139147
rect 74377 139124 74463 139147
rect 74209 139084 74234 139124
rect 74234 139084 74274 139124
rect 74274 139084 74295 139124
rect 74377 139084 74398 139124
rect 74398 139084 74438 139124
rect 74438 139084 74463 139124
rect 74209 139061 74295 139084
rect 74377 139061 74463 139084
rect 89329 139124 89415 139147
rect 89497 139124 89583 139147
rect 89329 139084 89354 139124
rect 89354 139084 89394 139124
rect 89394 139084 89415 139124
rect 89497 139084 89518 139124
rect 89518 139084 89558 139124
rect 89558 139084 89583 139124
rect 89329 139061 89415 139084
rect 89497 139061 89583 139084
rect 104449 139124 104535 139147
rect 104617 139124 104703 139147
rect 104449 139084 104474 139124
rect 104474 139084 104514 139124
rect 104514 139084 104535 139124
rect 104617 139084 104638 139124
rect 104638 139084 104678 139124
rect 104678 139084 104703 139124
rect 104449 139061 104535 139084
rect 104617 139061 104703 139084
rect 119569 139124 119655 139147
rect 119737 139124 119823 139147
rect 119569 139084 119594 139124
rect 119594 139084 119634 139124
rect 119634 139084 119655 139124
rect 119737 139084 119758 139124
rect 119758 139084 119798 139124
rect 119798 139084 119823 139124
rect 119569 139061 119655 139084
rect 119737 139061 119823 139084
rect 134689 139124 134775 139147
rect 134857 139124 134943 139147
rect 134689 139084 134714 139124
rect 134714 139084 134754 139124
rect 134754 139084 134775 139124
rect 134857 139084 134878 139124
rect 134878 139084 134918 139124
rect 134918 139084 134943 139124
rect 134689 139061 134775 139084
rect 134857 139061 134943 139084
rect 149809 139124 149895 139147
rect 149977 139124 150063 139147
rect 149809 139084 149834 139124
rect 149834 139084 149874 139124
rect 149874 139084 149895 139124
rect 149977 139084 149998 139124
rect 149998 139084 150038 139124
rect 150038 139084 150063 139124
rect 149809 139061 149895 139084
rect 149977 139061 150063 139084
rect 75449 138368 75535 138391
rect 75617 138368 75703 138391
rect 75449 138328 75474 138368
rect 75474 138328 75514 138368
rect 75514 138328 75535 138368
rect 75617 138328 75638 138368
rect 75638 138328 75678 138368
rect 75678 138328 75703 138368
rect 75449 138305 75535 138328
rect 75617 138305 75703 138328
rect 90569 138368 90655 138391
rect 90737 138368 90823 138391
rect 90569 138328 90594 138368
rect 90594 138328 90634 138368
rect 90634 138328 90655 138368
rect 90737 138328 90758 138368
rect 90758 138328 90798 138368
rect 90798 138328 90823 138368
rect 90569 138305 90655 138328
rect 90737 138305 90823 138328
rect 105689 138368 105775 138391
rect 105857 138368 105943 138391
rect 105689 138328 105714 138368
rect 105714 138328 105754 138368
rect 105754 138328 105775 138368
rect 105857 138328 105878 138368
rect 105878 138328 105918 138368
rect 105918 138328 105943 138368
rect 105689 138305 105775 138328
rect 105857 138305 105943 138328
rect 120809 138368 120895 138391
rect 120977 138368 121063 138391
rect 120809 138328 120834 138368
rect 120834 138328 120874 138368
rect 120874 138328 120895 138368
rect 120977 138328 120998 138368
rect 120998 138328 121038 138368
rect 121038 138328 121063 138368
rect 120809 138305 120895 138328
rect 120977 138305 121063 138328
rect 135929 138368 136015 138391
rect 136097 138368 136183 138391
rect 135929 138328 135954 138368
rect 135954 138328 135994 138368
rect 135994 138328 136015 138368
rect 136097 138328 136118 138368
rect 136118 138328 136158 138368
rect 136158 138328 136183 138368
rect 135929 138305 136015 138328
rect 136097 138305 136183 138328
rect 151049 138368 151135 138391
rect 151217 138368 151303 138391
rect 151049 138328 151074 138368
rect 151074 138328 151114 138368
rect 151114 138328 151135 138368
rect 151217 138328 151238 138368
rect 151238 138328 151278 138368
rect 151278 138328 151303 138368
rect 151049 138305 151135 138328
rect 151217 138305 151303 138328
rect 74209 137612 74295 137635
rect 74377 137612 74463 137635
rect 74209 137572 74234 137612
rect 74234 137572 74274 137612
rect 74274 137572 74295 137612
rect 74377 137572 74398 137612
rect 74398 137572 74438 137612
rect 74438 137572 74463 137612
rect 74209 137549 74295 137572
rect 74377 137549 74463 137572
rect 89329 137612 89415 137635
rect 89497 137612 89583 137635
rect 89329 137572 89354 137612
rect 89354 137572 89394 137612
rect 89394 137572 89415 137612
rect 89497 137572 89518 137612
rect 89518 137572 89558 137612
rect 89558 137572 89583 137612
rect 89329 137549 89415 137572
rect 89497 137549 89583 137572
rect 104449 137612 104535 137635
rect 104617 137612 104703 137635
rect 104449 137572 104474 137612
rect 104474 137572 104514 137612
rect 104514 137572 104535 137612
rect 104617 137572 104638 137612
rect 104638 137572 104678 137612
rect 104678 137572 104703 137612
rect 104449 137549 104535 137572
rect 104617 137549 104703 137572
rect 119569 137612 119655 137635
rect 119737 137612 119823 137635
rect 119569 137572 119594 137612
rect 119594 137572 119634 137612
rect 119634 137572 119655 137612
rect 119737 137572 119758 137612
rect 119758 137572 119798 137612
rect 119798 137572 119823 137612
rect 119569 137549 119655 137572
rect 119737 137549 119823 137572
rect 134689 137612 134775 137635
rect 134857 137612 134943 137635
rect 134689 137572 134714 137612
rect 134714 137572 134754 137612
rect 134754 137572 134775 137612
rect 134857 137572 134878 137612
rect 134878 137572 134918 137612
rect 134918 137572 134943 137612
rect 134689 137549 134775 137572
rect 134857 137549 134943 137572
rect 149809 137612 149895 137635
rect 149977 137612 150063 137635
rect 149809 137572 149834 137612
rect 149834 137572 149874 137612
rect 149874 137572 149895 137612
rect 149977 137572 149998 137612
rect 149998 137572 150038 137612
rect 150038 137572 150063 137612
rect 149809 137549 149895 137572
rect 149977 137549 150063 137572
rect 75449 136856 75535 136879
rect 75617 136856 75703 136879
rect 75449 136816 75474 136856
rect 75474 136816 75514 136856
rect 75514 136816 75535 136856
rect 75617 136816 75638 136856
rect 75638 136816 75678 136856
rect 75678 136816 75703 136856
rect 75449 136793 75535 136816
rect 75617 136793 75703 136816
rect 90569 136856 90655 136879
rect 90737 136856 90823 136879
rect 90569 136816 90594 136856
rect 90594 136816 90634 136856
rect 90634 136816 90655 136856
rect 90737 136816 90758 136856
rect 90758 136816 90798 136856
rect 90798 136816 90823 136856
rect 90569 136793 90655 136816
rect 90737 136793 90823 136816
rect 105689 136856 105775 136879
rect 105857 136856 105943 136879
rect 105689 136816 105714 136856
rect 105714 136816 105754 136856
rect 105754 136816 105775 136856
rect 105857 136816 105878 136856
rect 105878 136816 105918 136856
rect 105918 136816 105943 136856
rect 105689 136793 105775 136816
rect 105857 136793 105943 136816
rect 120809 136856 120895 136879
rect 120977 136856 121063 136879
rect 120809 136816 120834 136856
rect 120834 136816 120874 136856
rect 120874 136816 120895 136856
rect 120977 136816 120998 136856
rect 120998 136816 121038 136856
rect 121038 136816 121063 136856
rect 120809 136793 120895 136816
rect 120977 136793 121063 136816
rect 135929 136856 136015 136879
rect 136097 136856 136183 136879
rect 135929 136816 135954 136856
rect 135954 136816 135994 136856
rect 135994 136816 136015 136856
rect 136097 136816 136118 136856
rect 136118 136816 136158 136856
rect 136158 136816 136183 136856
rect 135929 136793 136015 136816
rect 136097 136793 136183 136816
rect 151049 136856 151135 136879
rect 151217 136856 151303 136879
rect 151049 136816 151074 136856
rect 151074 136816 151114 136856
rect 151114 136816 151135 136856
rect 151217 136816 151238 136856
rect 151238 136816 151278 136856
rect 151278 136816 151303 136856
rect 151049 136793 151135 136816
rect 151217 136793 151303 136816
rect 74209 136100 74295 136123
rect 74377 136100 74463 136123
rect 74209 136060 74234 136100
rect 74234 136060 74274 136100
rect 74274 136060 74295 136100
rect 74377 136060 74398 136100
rect 74398 136060 74438 136100
rect 74438 136060 74463 136100
rect 74209 136037 74295 136060
rect 74377 136037 74463 136060
rect 89329 136100 89415 136123
rect 89497 136100 89583 136123
rect 89329 136060 89354 136100
rect 89354 136060 89394 136100
rect 89394 136060 89415 136100
rect 89497 136060 89518 136100
rect 89518 136060 89558 136100
rect 89558 136060 89583 136100
rect 89329 136037 89415 136060
rect 89497 136037 89583 136060
rect 104449 136100 104535 136123
rect 104617 136100 104703 136123
rect 104449 136060 104474 136100
rect 104474 136060 104514 136100
rect 104514 136060 104535 136100
rect 104617 136060 104638 136100
rect 104638 136060 104678 136100
rect 104678 136060 104703 136100
rect 104449 136037 104535 136060
rect 104617 136037 104703 136060
rect 119569 136100 119655 136123
rect 119737 136100 119823 136123
rect 119569 136060 119594 136100
rect 119594 136060 119634 136100
rect 119634 136060 119655 136100
rect 119737 136060 119758 136100
rect 119758 136060 119798 136100
rect 119798 136060 119823 136100
rect 119569 136037 119655 136060
rect 119737 136037 119823 136060
rect 134689 136100 134775 136123
rect 134857 136100 134943 136123
rect 134689 136060 134714 136100
rect 134714 136060 134754 136100
rect 134754 136060 134775 136100
rect 134857 136060 134878 136100
rect 134878 136060 134918 136100
rect 134918 136060 134943 136100
rect 134689 136037 134775 136060
rect 134857 136037 134943 136060
rect 149809 136100 149895 136123
rect 149977 136100 150063 136123
rect 149809 136060 149834 136100
rect 149834 136060 149874 136100
rect 149874 136060 149895 136100
rect 149977 136060 149998 136100
rect 149998 136060 150038 136100
rect 150038 136060 150063 136100
rect 149809 136037 149895 136060
rect 149977 136037 150063 136060
rect 75449 135344 75535 135367
rect 75617 135344 75703 135367
rect 75449 135304 75474 135344
rect 75474 135304 75514 135344
rect 75514 135304 75535 135344
rect 75617 135304 75638 135344
rect 75638 135304 75678 135344
rect 75678 135304 75703 135344
rect 75449 135281 75535 135304
rect 75617 135281 75703 135304
rect 90569 135344 90655 135367
rect 90737 135344 90823 135367
rect 90569 135304 90594 135344
rect 90594 135304 90634 135344
rect 90634 135304 90655 135344
rect 90737 135304 90758 135344
rect 90758 135304 90798 135344
rect 90798 135304 90823 135344
rect 90569 135281 90655 135304
rect 90737 135281 90823 135304
rect 105689 135344 105775 135367
rect 105857 135344 105943 135367
rect 105689 135304 105714 135344
rect 105714 135304 105754 135344
rect 105754 135304 105775 135344
rect 105857 135304 105878 135344
rect 105878 135304 105918 135344
rect 105918 135304 105943 135344
rect 105689 135281 105775 135304
rect 105857 135281 105943 135304
rect 120809 135344 120895 135367
rect 120977 135344 121063 135367
rect 120809 135304 120834 135344
rect 120834 135304 120874 135344
rect 120874 135304 120895 135344
rect 120977 135304 120998 135344
rect 120998 135304 121038 135344
rect 121038 135304 121063 135344
rect 120809 135281 120895 135304
rect 120977 135281 121063 135304
rect 135929 135344 136015 135367
rect 136097 135344 136183 135367
rect 135929 135304 135954 135344
rect 135954 135304 135994 135344
rect 135994 135304 136015 135344
rect 136097 135304 136118 135344
rect 136118 135304 136158 135344
rect 136158 135304 136183 135344
rect 135929 135281 136015 135304
rect 136097 135281 136183 135304
rect 151049 135344 151135 135367
rect 151217 135344 151303 135367
rect 151049 135304 151074 135344
rect 151074 135304 151114 135344
rect 151114 135304 151135 135344
rect 151217 135304 151238 135344
rect 151238 135304 151278 135344
rect 151278 135304 151303 135344
rect 151049 135281 151135 135304
rect 151217 135281 151303 135304
rect 74209 134588 74295 134611
rect 74377 134588 74463 134611
rect 74209 134548 74234 134588
rect 74234 134548 74274 134588
rect 74274 134548 74295 134588
rect 74377 134548 74398 134588
rect 74398 134548 74438 134588
rect 74438 134548 74463 134588
rect 74209 134525 74295 134548
rect 74377 134525 74463 134548
rect 89329 134588 89415 134611
rect 89497 134588 89583 134611
rect 89329 134548 89354 134588
rect 89354 134548 89394 134588
rect 89394 134548 89415 134588
rect 89497 134548 89518 134588
rect 89518 134548 89558 134588
rect 89558 134548 89583 134588
rect 89329 134525 89415 134548
rect 89497 134525 89583 134548
rect 104449 134588 104535 134611
rect 104617 134588 104703 134611
rect 104449 134548 104474 134588
rect 104474 134548 104514 134588
rect 104514 134548 104535 134588
rect 104617 134548 104638 134588
rect 104638 134548 104678 134588
rect 104678 134548 104703 134588
rect 104449 134525 104535 134548
rect 104617 134525 104703 134548
rect 119569 134588 119655 134611
rect 119737 134588 119823 134611
rect 119569 134548 119594 134588
rect 119594 134548 119634 134588
rect 119634 134548 119655 134588
rect 119737 134548 119758 134588
rect 119758 134548 119798 134588
rect 119798 134548 119823 134588
rect 119569 134525 119655 134548
rect 119737 134525 119823 134548
rect 134689 134588 134775 134611
rect 134857 134588 134943 134611
rect 134689 134548 134714 134588
rect 134714 134548 134754 134588
rect 134754 134548 134775 134588
rect 134857 134548 134878 134588
rect 134878 134548 134918 134588
rect 134918 134548 134943 134588
rect 134689 134525 134775 134548
rect 134857 134525 134943 134548
rect 149809 134588 149895 134611
rect 149977 134588 150063 134611
rect 149809 134548 149834 134588
rect 149834 134548 149874 134588
rect 149874 134548 149895 134588
rect 149977 134548 149998 134588
rect 149998 134548 150038 134588
rect 150038 134548 150063 134588
rect 149809 134525 149895 134548
rect 149977 134525 150063 134548
rect 75449 133832 75535 133855
rect 75617 133832 75703 133855
rect 75449 133792 75474 133832
rect 75474 133792 75514 133832
rect 75514 133792 75535 133832
rect 75617 133792 75638 133832
rect 75638 133792 75678 133832
rect 75678 133792 75703 133832
rect 75449 133769 75535 133792
rect 75617 133769 75703 133792
rect 90569 133832 90655 133855
rect 90737 133832 90823 133855
rect 90569 133792 90594 133832
rect 90594 133792 90634 133832
rect 90634 133792 90655 133832
rect 90737 133792 90758 133832
rect 90758 133792 90798 133832
rect 90798 133792 90823 133832
rect 90569 133769 90655 133792
rect 90737 133769 90823 133792
rect 105689 133832 105775 133855
rect 105857 133832 105943 133855
rect 105689 133792 105714 133832
rect 105714 133792 105754 133832
rect 105754 133792 105775 133832
rect 105857 133792 105878 133832
rect 105878 133792 105918 133832
rect 105918 133792 105943 133832
rect 105689 133769 105775 133792
rect 105857 133769 105943 133792
rect 120809 133832 120895 133855
rect 120977 133832 121063 133855
rect 120809 133792 120834 133832
rect 120834 133792 120874 133832
rect 120874 133792 120895 133832
rect 120977 133792 120998 133832
rect 120998 133792 121038 133832
rect 121038 133792 121063 133832
rect 120809 133769 120895 133792
rect 120977 133769 121063 133792
rect 135929 133832 136015 133855
rect 136097 133832 136183 133855
rect 135929 133792 135954 133832
rect 135954 133792 135994 133832
rect 135994 133792 136015 133832
rect 136097 133792 136118 133832
rect 136118 133792 136158 133832
rect 136158 133792 136183 133832
rect 135929 133769 136015 133792
rect 136097 133769 136183 133792
rect 151049 133832 151135 133855
rect 151217 133832 151303 133855
rect 151049 133792 151074 133832
rect 151074 133792 151114 133832
rect 151114 133792 151135 133832
rect 151217 133792 151238 133832
rect 151238 133792 151278 133832
rect 151278 133792 151303 133832
rect 151049 133769 151135 133792
rect 151217 133769 151303 133792
rect 74209 133076 74295 133099
rect 74377 133076 74463 133099
rect 74209 133036 74234 133076
rect 74234 133036 74274 133076
rect 74274 133036 74295 133076
rect 74377 133036 74398 133076
rect 74398 133036 74438 133076
rect 74438 133036 74463 133076
rect 74209 133013 74295 133036
rect 74377 133013 74463 133036
rect 89329 133076 89415 133099
rect 89497 133076 89583 133099
rect 89329 133036 89354 133076
rect 89354 133036 89394 133076
rect 89394 133036 89415 133076
rect 89497 133036 89518 133076
rect 89518 133036 89558 133076
rect 89558 133036 89583 133076
rect 89329 133013 89415 133036
rect 89497 133013 89583 133036
rect 104449 133076 104535 133099
rect 104617 133076 104703 133099
rect 104449 133036 104474 133076
rect 104474 133036 104514 133076
rect 104514 133036 104535 133076
rect 104617 133036 104638 133076
rect 104638 133036 104678 133076
rect 104678 133036 104703 133076
rect 104449 133013 104535 133036
rect 104617 133013 104703 133036
rect 119569 133076 119655 133099
rect 119737 133076 119823 133099
rect 119569 133036 119594 133076
rect 119594 133036 119634 133076
rect 119634 133036 119655 133076
rect 119737 133036 119758 133076
rect 119758 133036 119798 133076
rect 119798 133036 119823 133076
rect 119569 133013 119655 133036
rect 119737 133013 119823 133036
rect 134689 133076 134775 133099
rect 134857 133076 134943 133099
rect 134689 133036 134714 133076
rect 134714 133036 134754 133076
rect 134754 133036 134775 133076
rect 134857 133036 134878 133076
rect 134878 133036 134918 133076
rect 134918 133036 134943 133076
rect 134689 133013 134775 133036
rect 134857 133013 134943 133036
rect 149809 133076 149895 133099
rect 149977 133076 150063 133099
rect 149809 133036 149834 133076
rect 149834 133036 149874 133076
rect 149874 133036 149895 133076
rect 149977 133036 149998 133076
rect 149998 133036 150038 133076
rect 150038 133036 150063 133076
rect 149809 133013 149895 133036
rect 149977 133013 150063 133036
rect 75449 132320 75535 132343
rect 75617 132320 75703 132343
rect 75449 132280 75474 132320
rect 75474 132280 75514 132320
rect 75514 132280 75535 132320
rect 75617 132280 75638 132320
rect 75638 132280 75678 132320
rect 75678 132280 75703 132320
rect 75449 132257 75535 132280
rect 75617 132257 75703 132280
rect 90569 132320 90655 132343
rect 90737 132320 90823 132343
rect 90569 132280 90594 132320
rect 90594 132280 90634 132320
rect 90634 132280 90655 132320
rect 90737 132280 90758 132320
rect 90758 132280 90798 132320
rect 90798 132280 90823 132320
rect 90569 132257 90655 132280
rect 90737 132257 90823 132280
rect 105689 132320 105775 132343
rect 105857 132320 105943 132343
rect 105689 132280 105714 132320
rect 105714 132280 105754 132320
rect 105754 132280 105775 132320
rect 105857 132280 105878 132320
rect 105878 132280 105918 132320
rect 105918 132280 105943 132320
rect 105689 132257 105775 132280
rect 105857 132257 105943 132280
rect 120809 132320 120895 132343
rect 120977 132320 121063 132343
rect 120809 132280 120834 132320
rect 120834 132280 120874 132320
rect 120874 132280 120895 132320
rect 120977 132280 120998 132320
rect 120998 132280 121038 132320
rect 121038 132280 121063 132320
rect 120809 132257 120895 132280
rect 120977 132257 121063 132280
rect 135929 132320 136015 132343
rect 136097 132320 136183 132343
rect 135929 132280 135954 132320
rect 135954 132280 135994 132320
rect 135994 132280 136015 132320
rect 136097 132280 136118 132320
rect 136118 132280 136158 132320
rect 136158 132280 136183 132320
rect 135929 132257 136015 132280
rect 136097 132257 136183 132280
rect 151049 132320 151135 132343
rect 151217 132320 151303 132343
rect 151049 132280 151074 132320
rect 151074 132280 151114 132320
rect 151114 132280 151135 132320
rect 151217 132280 151238 132320
rect 151238 132280 151278 132320
rect 151278 132280 151303 132320
rect 151049 132257 151135 132280
rect 151217 132257 151303 132280
rect 74209 131564 74295 131587
rect 74377 131564 74463 131587
rect 74209 131524 74234 131564
rect 74234 131524 74274 131564
rect 74274 131524 74295 131564
rect 74377 131524 74398 131564
rect 74398 131524 74438 131564
rect 74438 131524 74463 131564
rect 74209 131501 74295 131524
rect 74377 131501 74463 131524
rect 89329 131564 89415 131587
rect 89497 131564 89583 131587
rect 89329 131524 89354 131564
rect 89354 131524 89394 131564
rect 89394 131524 89415 131564
rect 89497 131524 89518 131564
rect 89518 131524 89558 131564
rect 89558 131524 89583 131564
rect 89329 131501 89415 131524
rect 89497 131501 89583 131524
rect 104449 131564 104535 131587
rect 104617 131564 104703 131587
rect 104449 131524 104474 131564
rect 104474 131524 104514 131564
rect 104514 131524 104535 131564
rect 104617 131524 104638 131564
rect 104638 131524 104678 131564
rect 104678 131524 104703 131564
rect 104449 131501 104535 131524
rect 104617 131501 104703 131524
rect 119569 131564 119655 131587
rect 119737 131564 119823 131587
rect 119569 131524 119594 131564
rect 119594 131524 119634 131564
rect 119634 131524 119655 131564
rect 119737 131524 119758 131564
rect 119758 131524 119798 131564
rect 119798 131524 119823 131564
rect 119569 131501 119655 131524
rect 119737 131501 119823 131524
rect 134689 131564 134775 131587
rect 134857 131564 134943 131587
rect 134689 131524 134714 131564
rect 134714 131524 134754 131564
rect 134754 131524 134775 131564
rect 134857 131524 134878 131564
rect 134878 131524 134918 131564
rect 134918 131524 134943 131564
rect 134689 131501 134775 131524
rect 134857 131501 134943 131524
rect 149809 131564 149895 131587
rect 149977 131564 150063 131587
rect 149809 131524 149834 131564
rect 149834 131524 149874 131564
rect 149874 131524 149895 131564
rect 149977 131524 149998 131564
rect 149998 131524 150038 131564
rect 150038 131524 150063 131564
rect 149809 131501 149895 131524
rect 149977 131501 150063 131524
rect 75449 130808 75535 130831
rect 75617 130808 75703 130831
rect 75449 130768 75474 130808
rect 75474 130768 75514 130808
rect 75514 130768 75535 130808
rect 75617 130768 75638 130808
rect 75638 130768 75678 130808
rect 75678 130768 75703 130808
rect 75449 130745 75535 130768
rect 75617 130745 75703 130768
rect 90569 130808 90655 130831
rect 90737 130808 90823 130831
rect 90569 130768 90594 130808
rect 90594 130768 90634 130808
rect 90634 130768 90655 130808
rect 90737 130768 90758 130808
rect 90758 130768 90798 130808
rect 90798 130768 90823 130808
rect 90569 130745 90655 130768
rect 90737 130745 90823 130768
rect 105689 130808 105775 130831
rect 105857 130808 105943 130831
rect 105689 130768 105714 130808
rect 105714 130768 105754 130808
rect 105754 130768 105775 130808
rect 105857 130768 105878 130808
rect 105878 130768 105918 130808
rect 105918 130768 105943 130808
rect 105689 130745 105775 130768
rect 105857 130745 105943 130768
rect 120809 130808 120895 130831
rect 120977 130808 121063 130831
rect 120809 130768 120834 130808
rect 120834 130768 120874 130808
rect 120874 130768 120895 130808
rect 120977 130768 120998 130808
rect 120998 130768 121038 130808
rect 121038 130768 121063 130808
rect 120809 130745 120895 130768
rect 120977 130745 121063 130768
rect 135929 130808 136015 130831
rect 136097 130808 136183 130831
rect 135929 130768 135954 130808
rect 135954 130768 135994 130808
rect 135994 130768 136015 130808
rect 136097 130768 136118 130808
rect 136118 130768 136158 130808
rect 136158 130768 136183 130808
rect 135929 130745 136015 130768
rect 136097 130745 136183 130768
rect 151049 130808 151135 130831
rect 151217 130808 151303 130831
rect 151049 130768 151074 130808
rect 151074 130768 151114 130808
rect 151114 130768 151135 130808
rect 151217 130768 151238 130808
rect 151238 130768 151278 130808
rect 151278 130768 151303 130808
rect 151049 130745 151135 130768
rect 151217 130745 151303 130768
rect 74209 130052 74295 130075
rect 74377 130052 74463 130075
rect 74209 130012 74234 130052
rect 74234 130012 74274 130052
rect 74274 130012 74295 130052
rect 74377 130012 74398 130052
rect 74398 130012 74438 130052
rect 74438 130012 74463 130052
rect 74209 129989 74295 130012
rect 74377 129989 74463 130012
rect 89329 130052 89415 130075
rect 89497 130052 89583 130075
rect 89329 130012 89354 130052
rect 89354 130012 89394 130052
rect 89394 130012 89415 130052
rect 89497 130012 89518 130052
rect 89518 130012 89558 130052
rect 89558 130012 89583 130052
rect 89329 129989 89415 130012
rect 89497 129989 89583 130012
rect 104449 130052 104535 130075
rect 104617 130052 104703 130075
rect 104449 130012 104474 130052
rect 104474 130012 104514 130052
rect 104514 130012 104535 130052
rect 104617 130012 104638 130052
rect 104638 130012 104678 130052
rect 104678 130012 104703 130052
rect 104449 129989 104535 130012
rect 104617 129989 104703 130012
rect 119569 130052 119655 130075
rect 119737 130052 119823 130075
rect 119569 130012 119594 130052
rect 119594 130012 119634 130052
rect 119634 130012 119655 130052
rect 119737 130012 119758 130052
rect 119758 130012 119798 130052
rect 119798 130012 119823 130052
rect 119569 129989 119655 130012
rect 119737 129989 119823 130012
rect 134689 130052 134775 130075
rect 134857 130052 134943 130075
rect 134689 130012 134714 130052
rect 134714 130012 134754 130052
rect 134754 130012 134775 130052
rect 134857 130012 134878 130052
rect 134878 130012 134918 130052
rect 134918 130012 134943 130052
rect 134689 129989 134775 130012
rect 134857 129989 134943 130012
rect 149809 130052 149895 130075
rect 149977 130052 150063 130075
rect 149809 130012 149834 130052
rect 149834 130012 149874 130052
rect 149874 130012 149895 130052
rect 149977 130012 149998 130052
rect 149998 130012 150038 130052
rect 150038 130012 150063 130052
rect 149809 129989 149895 130012
rect 149977 129989 150063 130012
rect 75449 129296 75535 129319
rect 75617 129296 75703 129319
rect 75449 129256 75474 129296
rect 75474 129256 75514 129296
rect 75514 129256 75535 129296
rect 75617 129256 75638 129296
rect 75638 129256 75678 129296
rect 75678 129256 75703 129296
rect 75449 129233 75535 129256
rect 75617 129233 75703 129256
rect 90569 129296 90655 129319
rect 90737 129296 90823 129319
rect 90569 129256 90594 129296
rect 90594 129256 90634 129296
rect 90634 129256 90655 129296
rect 90737 129256 90758 129296
rect 90758 129256 90798 129296
rect 90798 129256 90823 129296
rect 90569 129233 90655 129256
rect 90737 129233 90823 129256
rect 105689 129296 105775 129319
rect 105857 129296 105943 129319
rect 105689 129256 105714 129296
rect 105714 129256 105754 129296
rect 105754 129256 105775 129296
rect 105857 129256 105878 129296
rect 105878 129256 105918 129296
rect 105918 129256 105943 129296
rect 105689 129233 105775 129256
rect 105857 129233 105943 129256
rect 120809 129296 120895 129319
rect 120977 129296 121063 129319
rect 120809 129256 120834 129296
rect 120834 129256 120874 129296
rect 120874 129256 120895 129296
rect 120977 129256 120998 129296
rect 120998 129256 121038 129296
rect 121038 129256 121063 129296
rect 120809 129233 120895 129256
rect 120977 129233 121063 129256
rect 135929 129296 136015 129319
rect 136097 129296 136183 129319
rect 135929 129256 135954 129296
rect 135954 129256 135994 129296
rect 135994 129256 136015 129296
rect 136097 129256 136118 129296
rect 136118 129256 136158 129296
rect 136158 129256 136183 129296
rect 135929 129233 136015 129256
rect 136097 129233 136183 129256
rect 151049 129296 151135 129319
rect 151217 129296 151303 129319
rect 151049 129256 151074 129296
rect 151074 129256 151114 129296
rect 151114 129256 151135 129296
rect 151217 129256 151238 129296
rect 151238 129256 151278 129296
rect 151278 129256 151303 129296
rect 151049 129233 151135 129256
rect 151217 129233 151303 129256
rect 74209 128540 74295 128563
rect 74377 128540 74463 128563
rect 74209 128500 74234 128540
rect 74234 128500 74274 128540
rect 74274 128500 74295 128540
rect 74377 128500 74398 128540
rect 74398 128500 74438 128540
rect 74438 128500 74463 128540
rect 74209 128477 74295 128500
rect 74377 128477 74463 128500
rect 89329 128540 89415 128563
rect 89497 128540 89583 128563
rect 89329 128500 89354 128540
rect 89354 128500 89394 128540
rect 89394 128500 89415 128540
rect 89497 128500 89518 128540
rect 89518 128500 89558 128540
rect 89558 128500 89583 128540
rect 89329 128477 89415 128500
rect 89497 128477 89583 128500
rect 104449 128540 104535 128563
rect 104617 128540 104703 128563
rect 104449 128500 104474 128540
rect 104474 128500 104514 128540
rect 104514 128500 104535 128540
rect 104617 128500 104638 128540
rect 104638 128500 104678 128540
rect 104678 128500 104703 128540
rect 104449 128477 104535 128500
rect 104617 128477 104703 128500
rect 119569 128540 119655 128563
rect 119737 128540 119823 128563
rect 119569 128500 119594 128540
rect 119594 128500 119634 128540
rect 119634 128500 119655 128540
rect 119737 128500 119758 128540
rect 119758 128500 119798 128540
rect 119798 128500 119823 128540
rect 119569 128477 119655 128500
rect 119737 128477 119823 128500
rect 134689 128540 134775 128563
rect 134857 128540 134943 128563
rect 134689 128500 134714 128540
rect 134714 128500 134754 128540
rect 134754 128500 134775 128540
rect 134857 128500 134878 128540
rect 134878 128500 134918 128540
rect 134918 128500 134943 128540
rect 134689 128477 134775 128500
rect 134857 128477 134943 128500
rect 149809 128540 149895 128563
rect 149977 128540 150063 128563
rect 149809 128500 149834 128540
rect 149834 128500 149874 128540
rect 149874 128500 149895 128540
rect 149977 128500 149998 128540
rect 149998 128500 150038 128540
rect 150038 128500 150063 128540
rect 149809 128477 149895 128500
rect 149977 128477 150063 128500
rect 75449 127784 75535 127807
rect 75617 127784 75703 127807
rect 75449 127744 75474 127784
rect 75474 127744 75514 127784
rect 75514 127744 75535 127784
rect 75617 127744 75638 127784
rect 75638 127744 75678 127784
rect 75678 127744 75703 127784
rect 75449 127721 75535 127744
rect 75617 127721 75703 127744
rect 90569 127784 90655 127807
rect 90737 127784 90823 127807
rect 90569 127744 90594 127784
rect 90594 127744 90634 127784
rect 90634 127744 90655 127784
rect 90737 127744 90758 127784
rect 90758 127744 90798 127784
rect 90798 127744 90823 127784
rect 90569 127721 90655 127744
rect 90737 127721 90823 127744
rect 105689 127784 105775 127807
rect 105857 127784 105943 127807
rect 105689 127744 105714 127784
rect 105714 127744 105754 127784
rect 105754 127744 105775 127784
rect 105857 127744 105878 127784
rect 105878 127744 105918 127784
rect 105918 127744 105943 127784
rect 105689 127721 105775 127744
rect 105857 127721 105943 127744
rect 120809 127784 120895 127807
rect 120977 127784 121063 127807
rect 120809 127744 120834 127784
rect 120834 127744 120874 127784
rect 120874 127744 120895 127784
rect 120977 127744 120998 127784
rect 120998 127744 121038 127784
rect 121038 127744 121063 127784
rect 120809 127721 120895 127744
rect 120977 127721 121063 127744
rect 135929 127784 136015 127807
rect 136097 127784 136183 127807
rect 135929 127744 135954 127784
rect 135954 127744 135994 127784
rect 135994 127744 136015 127784
rect 136097 127744 136118 127784
rect 136118 127744 136158 127784
rect 136158 127744 136183 127784
rect 135929 127721 136015 127744
rect 136097 127721 136183 127744
rect 151049 127784 151135 127807
rect 151217 127784 151303 127807
rect 151049 127744 151074 127784
rect 151074 127744 151114 127784
rect 151114 127744 151135 127784
rect 151217 127744 151238 127784
rect 151238 127744 151278 127784
rect 151278 127744 151303 127784
rect 151049 127721 151135 127744
rect 151217 127721 151303 127744
rect 74209 127028 74295 127051
rect 74377 127028 74463 127051
rect 74209 126988 74234 127028
rect 74234 126988 74274 127028
rect 74274 126988 74295 127028
rect 74377 126988 74398 127028
rect 74398 126988 74438 127028
rect 74438 126988 74463 127028
rect 74209 126965 74295 126988
rect 74377 126965 74463 126988
rect 89329 127028 89415 127051
rect 89497 127028 89583 127051
rect 89329 126988 89354 127028
rect 89354 126988 89394 127028
rect 89394 126988 89415 127028
rect 89497 126988 89518 127028
rect 89518 126988 89558 127028
rect 89558 126988 89583 127028
rect 89329 126965 89415 126988
rect 89497 126965 89583 126988
rect 104449 127028 104535 127051
rect 104617 127028 104703 127051
rect 104449 126988 104474 127028
rect 104474 126988 104514 127028
rect 104514 126988 104535 127028
rect 104617 126988 104638 127028
rect 104638 126988 104678 127028
rect 104678 126988 104703 127028
rect 104449 126965 104535 126988
rect 104617 126965 104703 126988
rect 119569 127028 119655 127051
rect 119737 127028 119823 127051
rect 119569 126988 119594 127028
rect 119594 126988 119634 127028
rect 119634 126988 119655 127028
rect 119737 126988 119758 127028
rect 119758 126988 119798 127028
rect 119798 126988 119823 127028
rect 119569 126965 119655 126988
rect 119737 126965 119823 126988
rect 134689 127028 134775 127051
rect 134857 127028 134943 127051
rect 134689 126988 134714 127028
rect 134714 126988 134754 127028
rect 134754 126988 134775 127028
rect 134857 126988 134878 127028
rect 134878 126988 134918 127028
rect 134918 126988 134943 127028
rect 134689 126965 134775 126988
rect 134857 126965 134943 126988
rect 149809 127028 149895 127051
rect 149977 127028 150063 127051
rect 149809 126988 149834 127028
rect 149834 126988 149874 127028
rect 149874 126988 149895 127028
rect 149977 126988 149998 127028
rect 149998 126988 150038 127028
rect 150038 126988 150063 127028
rect 149809 126965 149895 126988
rect 149977 126965 150063 126988
rect 75449 126272 75535 126295
rect 75617 126272 75703 126295
rect 75449 126232 75474 126272
rect 75474 126232 75514 126272
rect 75514 126232 75535 126272
rect 75617 126232 75638 126272
rect 75638 126232 75678 126272
rect 75678 126232 75703 126272
rect 75449 126209 75535 126232
rect 75617 126209 75703 126232
rect 90569 126272 90655 126295
rect 90737 126272 90823 126295
rect 90569 126232 90594 126272
rect 90594 126232 90634 126272
rect 90634 126232 90655 126272
rect 90737 126232 90758 126272
rect 90758 126232 90798 126272
rect 90798 126232 90823 126272
rect 90569 126209 90655 126232
rect 90737 126209 90823 126232
rect 105689 126272 105775 126295
rect 105857 126272 105943 126295
rect 105689 126232 105714 126272
rect 105714 126232 105754 126272
rect 105754 126232 105775 126272
rect 105857 126232 105878 126272
rect 105878 126232 105918 126272
rect 105918 126232 105943 126272
rect 105689 126209 105775 126232
rect 105857 126209 105943 126232
rect 120809 126272 120895 126295
rect 120977 126272 121063 126295
rect 120809 126232 120834 126272
rect 120834 126232 120874 126272
rect 120874 126232 120895 126272
rect 120977 126232 120998 126272
rect 120998 126232 121038 126272
rect 121038 126232 121063 126272
rect 120809 126209 120895 126232
rect 120977 126209 121063 126232
rect 135929 126272 136015 126295
rect 136097 126272 136183 126295
rect 135929 126232 135954 126272
rect 135954 126232 135994 126272
rect 135994 126232 136015 126272
rect 136097 126232 136118 126272
rect 136118 126232 136158 126272
rect 136158 126232 136183 126272
rect 135929 126209 136015 126232
rect 136097 126209 136183 126232
rect 151049 126272 151135 126295
rect 151217 126272 151303 126295
rect 151049 126232 151074 126272
rect 151074 126232 151114 126272
rect 151114 126232 151135 126272
rect 151217 126232 151238 126272
rect 151238 126232 151278 126272
rect 151278 126232 151303 126272
rect 151049 126209 151135 126232
rect 151217 126209 151303 126232
rect 74209 125516 74295 125539
rect 74377 125516 74463 125539
rect 74209 125476 74234 125516
rect 74234 125476 74274 125516
rect 74274 125476 74295 125516
rect 74377 125476 74398 125516
rect 74398 125476 74438 125516
rect 74438 125476 74463 125516
rect 74209 125453 74295 125476
rect 74377 125453 74463 125476
rect 89329 125516 89415 125539
rect 89497 125516 89583 125539
rect 89329 125476 89354 125516
rect 89354 125476 89394 125516
rect 89394 125476 89415 125516
rect 89497 125476 89518 125516
rect 89518 125476 89558 125516
rect 89558 125476 89583 125516
rect 89329 125453 89415 125476
rect 89497 125453 89583 125476
rect 104449 125516 104535 125539
rect 104617 125516 104703 125539
rect 104449 125476 104474 125516
rect 104474 125476 104514 125516
rect 104514 125476 104535 125516
rect 104617 125476 104638 125516
rect 104638 125476 104678 125516
rect 104678 125476 104703 125516
rect 104449 125453 104535 125476
rect 104617 125453 104703 125476
rect 119569 125516 119655 125539
rect 119737 125516 119823 125539
rect 119569 125476 119594 125516
rect 119594 125476 119634 125516
rect 119634 125476 119655 125516
rect 119737 125476 119758 125516
rect 119758 125476 119798 125516
rect 119798 125476 119823 125516
rect 119569 125453 119655 125476
rect 119737 125453 119823 125476
rect 134689 125516 134775 125539
rect 134857 125516 134943 125539
rect 134689 125476 134714 125516
rect 134714 125476 134754 125516
rect 134754 125476 134775 125516
rect 134857 125476 134878 125516
rect 134878 125476 134918 125516
rect 134918 125476 134943 125516
rect 134689 125453 134775 125476
rect 134857 125453 134943 125476
rect 149809 125516 149895 125539
rect 149977 125516 150063 125539
rect 149809 125476 149834 125516
rect 149834 125476 149874 125516
rect 149874 125476 149895 125516
rect 149977 125476 149998 125516
rect 149998 125476 150038 125516
rect 150038 125476 150063 125516
rect 149809 125453 149895 125476
rect 149977 125453 150063 125476
rect 75449 124760 75535 124783
rect 75617 124760 75703 124783
rect 75449 124720 75474 124760
rect 75474 124720 75514 124760
rect 75514 124720 75535 124760
rect 75617 124720 75638 124760
rect 75638 124720 75678 124760
rect 75678 124720 75703 124760
rect 75449 124697 75535 124720
rect 75617 124697 75703 124720
rect 90569 124760 90655 124783
rect 90737 124760 90823 124783
rect 90569 124720 90594 124760
rect 90594 124720 90634 124760
rect 90634 124720 90655 124760
rect 90737 124720 90758 124760
rect 90758 124720 90798 124760
rect 90798 124720 90823 124760
rect 90569 124697 90655 124720
rect 90737 124697 90823 124720
rect 105689 124760 105775 124783
rect 105857 124760 105943 124783
rect 105689 124720 105714 124760
rect 105714 124720 105754 124760
rect 105754 124720 105775 124760
rect 105857 124720 105878 124760
rect 105878 124720 105918 124760
rect 105918 124720 105943 124760
rect 105689 124697 105775 124720
rect 105857 124697 105943 124720
rect 120809 124760 120895 124783
rect 120977 124760 121063 124783
rect 120809 124720 120834 124760
rect 120834 124720 120874 124760
rect 120874 124720 120895 124760
rect 120977 124720 120998 124760
rect 120998 124720 121038 124760
rect 121038 124720 121063 124760
rect 120809 124697 120895 124720
rect 120977 124697 121063 124720
rect 135929 124760 136015 124783
rect 136097 124760 136183 124783
rect 135929 124720 135954 124760
rect 135954 124720 135994 124760
rect 135994 124720 136015 124760
rect 136097 124720 136118 124760
rect 136118 124720 136158 124760
rect 136158 124720 136183 124760
rect 135929 124697 136015 124720
rect 136097 124697 136183 124720
rect 151049 124760 151135 124783
rect 151217 124760 151303 124783
rect 151049 124720 151074 124760
rect 151074 124720 151114 124760
rect 151114 124720 151135 124760
rect 151217 124720 151238 124760
rect 151238 124720 151278 124760
rect 151278 124720 151303 124760
rect 151049 124697 151135 124720
rect 151217 124697 151303 124720
rect 74209 124004 74295 124027
rect 74377 124004 74463 124027
rect 74209 123964 74234 124004
rect 74234 123964 74274 124004
rect 74274 123964 74295 124004
rect 74377 123964 74398 124004
rect 74398 123964 74438 124004
rect 74438 123964 74463 124004
rect 74209 123941 74295 123964
rect 74377 123941 74463 123964
rect 89329 124004 89415 124027
rect 89497 124004 89583 124027
rect 89329 123964 89354 124004
rect 89354 123964 89394 124004
rect 89394 123964 89415 124004
rect 89497 123964 89518 124004
rect 89518 123964 89558 124004
rect 89558 123964 89583 124004
rect 89329 123941 89415 123964
rect 89497 123941 89583 123964
rect 104449 124004 104535 124027
rect 104617 124004 104703 124027
rect 104449 123964 104474 124004
rect 104474 123964 104514 124004
rect 104514 123964 104535 124004
rect 104617 123964 104638 124004
rect 104638 123964 104678 124004
rect 104678 123964 104703 124004
rect 104449 123941 104535 123964
rect 104617 123941 104703 123964
rect 119569 124004 119655 124027
rect 119737 124004 119823 124027
rect 119569 123964 119594 124004
rect 119594 123964 119634 124004
rect 119634 123964 119655 124004
rect 119737 123964 119758 124004
rect 119758 123964 119798 124004
rect 119798 123964 119823 124004
rect 119569 123941 119655 123964
rect 119737 123941 119823 123964
rect 134689 124004 134775 124027
rect 134857 124004 134943 124027
rect 134689 123964 134714 124004
rect 134714 123964 134754 124004
rect 134754 123964 134775 124004
rect 134857 123964 134878 124004
rect 134878 123964 134918 124004
rect 134918 123964 134943 124004
rect 134689 123941 134775 123964
rect 134857 123941 134943 123964
rect 149809 124004 149895 124027
rect 149977 124004 150063 124027
rect 149809 123964 149834 124004
rect 149834 123964 149874 124004
rect 149874 123964 149895 124004
rect 149977 123964 149998 124004
rect 149998 123964 150038 124004
rect 150038 123964 150063 124004
rect 149809 123941 149895 123964
rect 149977 123941 150063 123964
rect 75449 123248 75535 123271
rect 75617 123248 75703 123271
rect 75449 123208 75474 123248
rect 75474 123208 75514 123248
rect 75514 123208 75535 123248
rect 75617 123208 75638 123248
rect 75638 123208 75678 123248
rect 75678 123208 75703 123248
rect 75449 123185 75535 123208
rect 75617 123185 75703 123208
rect 90569 123248 90655 123271
rect 90737 123248 90823 123271
rect 90569 123208 90594 123248
rect 90594 123208 90634 123248
rect 90634 123208 90655 123248
rect 90737 123208 90758 123248
rect 90758 123208 90798 123248
rect 90798 123208 90823 123248
rect 90569 123185 90655 123208
rect 90737 123185 90823 123208
rect 105689 123248 105775 123271
rect 105857 123248 105943 123271
rect 105689 123208 105714 123248
rect 105714 123208 105754 123248
rect 105754 123208 105775 123248
rect 105857 123208 105878 123248
rect 105878 123208 105918 123248
rect 105918 123208 105943 123248
rect 105689 123185 105775 123208
rect 105857 123185 105943 123208
rect 120809 123248 120895 123271
rect 120977 123248 121063 123271
rect 120809 123208 120834 123248
rect 120834 123208 120874 123248
rect 120874 123208 120895 123248
rect 120977 123208 120998 123248
rect 120998 123208 121038 123248
rect 121038 123208 121063 123248
rect 120809 123185 120895 123208
rect 120977 123185 121063 123208
rect 135929 123248 136015 123271
rect 136097 123248 136183 123271
rect 135929 123208 135954 123248
rect 135954 123208 135994 123248
rect 135994 123208 136015 123248
rect 136097 123208 136118 123248
rect 136118 123208 136158 123248
rect 136158 123208 136183 123248
rect 135929 123185 136015 123208
rect 136097 123185 136183 123208
rect 151049 123248 151135 123271
rect 151217 123248 151303 123271
rect 151049 123208 151074 123248
rect 151074 123208 151114 123248
rect 151114 123208 151135 123248
rect 151217 123208 151238 123248
rect 151238 123208 151278 123248
rect 151278 123208 151303 123248
rect 151049 123185 151135 123208
rect 151217 123185 151303 123208
rect 74209 122492 74295 122515
rect 74377 122492 74463 122515
rect 74209 122452 74234 122492
rect 74234 122452 74274 122492
rect 74274 122452 74295 122492
rect 74377 122452 74398 122492
rect 74398 122452 74438 122492
rect 74438 122452 74463 122492
rect 74209 122429 74295 122452
rect 74377 122429 74463 122452
rect 89329 122492 89415 122515
rect 89497 122492 89583 122515
rect 89329 122452 89354 122492
rect 89354 122452 89394 122492
rect 89394 122452 89415 122492
rect 89497 122452 89518 122492
rect 89518 122452 89558 122492
rect 89558 122452 89583 122492
rect 89329 122429 89415 122452
rect 89497 122429 89583 122452
rect 104449 122492 104535 122515
rect 104617 122492 104703 122515
rect 104449 122452 104474 122492
rect 104474 122452 104514 122492
rect 104514 122452 104535 122492
rect 104617 122452 104638 122492
rect 104638 122452 104678 122492
rect 104678 122452 104703 122492
rect 104449 122429 104535 122452
rect 104617 122429 104703 122452
rect 119569 122492 119655 122515
rect 119737 122492 119823 122515
rect 119569 122452 119594 122492
rect 119594 122452 119634 122492
rect 119634 122452 119655 122492
rect 119737 122452 119758 122492
rect 119758 122452 119798 122492
rect 119798 122452 119823 122492
rect 119569 122429 119655 122452
rect 119737 122429 119823 122452
rect 134689 122492 134775 122515
rect 134857 122492 134943 122515
rect 134689 122452 134714 122492
rect 134714 122452 134754 122492
rect 134754 122452 134775 122492
rect 134857 122452 134878 122492
rect 134878 122452 134918 122492
rect 134918 122452 134943 122492
rect 134689 122429 134775 122452
rect 134857 122429 134943 122452
rect 149809 122492 149895 122515
rect 149977 122492 150063 122515
rect 149809 122452 149834 122492
rect 149834 122452 149874 122492
rect 149874 122452 149895 122492
rect 149977 122452 149998 122492
rect 149998 122452 150038 122492
rect 150038 122452 150063 122492
rect 149809 122429 149895 122452
rect 149977 122429 150063 122452
rect 75449 121736 75535 121759
rect 75617 121736 75703 121759
rect 75449 121696 75474 121736
rect 75474 121696 75514 121736
rect 75514 121696 75535 121736
rect 75617 121696 75638 121736
rect 75638 121696 75678 121736
rect 75678 121696 75703 121736
rect 75449 121673 75535 121696
rect 75617 121673 75703 121696
rect 90569 121736 90655 121759
rect 90737 121736 90823 121759
rect 90569 121696 90594 121736
rect 90594 121696 90634 121736
rect 90634 121696 90655 121736
rect 90737 121696 90758 121736
rect 90758 121696 90798 121736
rect 90798 121696 90823 121736
rect 90569 121673 90655 121696
rect 90737 121673 90823 121696
rect 105689 121736 105775 121759
rect 105857 121736 105943 121759
rect 105689 121696 105714 121736
rect 105714 121696 105754 121736
rect 105754 121696 105775 121736
rect 105857 121696 105878 121736
rect 105878 121696 105918 121736
rect 105918 121696 105943 121736
rect 105689 121673 105775 121696
rect 105857 121673 105943 121696
rect 120809 121736 120895 121759
rect 120977 121736 121063 121759
rect 120809 121696 120834 121736
rect 120834 121696 120874 121736
rect 120874 121696 120895 121736
rect 120977 121696 120998 121736
rect 120998 121696 121038 121736
rect 121038 121696 121063 121736
rect 120809 121673 120895 121696
rect 120977 121673 121063 121696
rect 135929 121736 136015 121759
rect 136097 121736 136183 121759
rect 135929 121696 135954 121736
rect 135954 121696 135994 121736
rect 135994 121696 136015 121736
rect 136097 121696 136118 121736
rect 136118 121696 136158 121736
rect 136158 121696 136183 121736
rect 135929 121673 136015 121696
rect 136097 121673 136183 121696
rect 151049 121736 151135 121759
rect 151217 121736 151303 121759
rect 151049 121696 151074 121736
rect 151074 121696 151114 121736
rect 151114 121696 151135 121736
rect 151217 121696 151238 121736
rect 151238 121696 151278 121736
rect 151278 121696 151303 121736
rect 151049 121673 151135 121696
rect 151217 121673 151303 121696
rect 74209 120980 74295 121003
rect 74377 120980 74463 121003
rect 74209 120940 74234 120980
rect 74234 120940 74274 120980
rect 74274 120940 74295 120980
rect 74377 120940 74398 120980
rect 74398 120940 74438 120980
rect 74438 120940 74463 120980
rect 74209 120917 74295 120940
rect 74377 120917 74463 120940
rect 89329 120980 89415 121003
rect 89497 120980 89583 121003
rect 89329 120940 89354 120980
rect 89354 120940 89394 120980
rect 89394 120940 89415 120980
rect 89497 120940 89518 120980
rect 89518 120940 89558 120980
rect 89558 120940 89583 120980
rect 89329 120917 89415 120940
rect 89497 120917 89583 120940
rect 104449 120980 104535 121003
rect 104617 120980 104703 121003
rect 104449 120940 104474 120980
rect 104474 120940 104514 120980
rect 104514 120940 104535 120980
rect 104617 120940 104638 120980
rect 104638 120940 104678 120980
rect 104678 120940 104703 120980
rect 104449 120917 104535 120940
rect 104617 120917 104703 120940
rect 119569 120980 119655 121003
rect 119737 120980 119823 121003
rect 119569 120940 119594 120980
rect 119594 120940 119634 120980
rect 119634 120940 119655 120980
rect 119737 120940 119758 120980
rect 119758 120940 119798 120980
rect 119798 120940 119823 120980
rect 119569 120917 119655 120940
rect 119737 120917 119823 120940
rect 134689 120980 134775 121003
rect 134857 120980 134943 121003
rect 134689 120940 134714 120980
rect 134714 120940 134754 120980
rect 134754 120940 134775 120980
rect 134857 120940 134878 120980
rect 134878 120940 134918 120980
rect 134918 120940 134943 120980
rect 134689 120917 134775 120940
rect 134857 120917 134943 120940
rect 149809 120980 149895 121003
rect 149977 120980 150063 121003
rect 149809 120940 149834 120980
rect 149834 120940 149874 120980
rect 149874 120940 149895 120980
rect 149977 120940 149998 120980
rect 149998 120940 150038 120980
rect 150038 120940 150063 120980
rect 149809 120917 149895 120940
rect 149977 120917 150063 120940
rect 75449 120224 75535 120247
rect 75617 120224 75703 120247
rect 75449 120184 75474 120224
rect 75474 120184 75514 120224
rect 75514 120184 75535 120224
rect 75617 120184 75638 120224
rect 75638 120184 75678 120224
rect 75678 120184 75703 120224
rect 75449 120161 75535 120184
rect 75617 120161 75703 120184
rect 90569 120224 90655 120247
rect 90737 120224 90823 120247
rect 90569 120184 90594 120224
rect 90594 120184 90634 120224
rect 90634 120184 90655 120224
rect 90737 120184 90758 120224
rect 90758 120184 90798 120224
rect 90798 120184 90823 120224
rect 90569 120161 90655 120184
rect 90737 120161 90823 120184
rect 105689 120224 105775 120247
rect 105857 120224 105943 120247
rect 105689 120184 105714 120224
rect 105714 120184 105754 120224
rect 105754 120184 105775 120224
rect 105857 120184 105878 120224
rect 105878 120184 105918 120224
rect 105918 120184 105943 120224
rect 105689 120161 105775 120184
rect 105857 120161 105943 120184
rect 120809 120224 120895 120247
rect 120977 120224 121063 120247
rect 120809 120184 120834 120224
rect 120834 120184 120874 120224
rect 120874 120184 120895 120224
rect 120977 120184 120998 120224
rect 120998 120184 121038 120224
rect 121038 120184 121063 120224
rect 120809 120161 120895 120184
rect 120977 120161 121063 120184
rect 135929 120224 136015 120247
rect 136097 120224 136183 120247
rect 135929 120184 135954 120224
rect 135954 120184 135994 120224
rect 135994 120184 136015 120224
rect 136097 120184 136118 120224
rect 136118 120184 136158 120224
rect 136158 120184 136183 120224
rect 135929 120161 136015 120184
rect 136097 120161 136183 120184
rect 151049 120224 151135 120247
rect 151217 120224 151303 120247
rect 151049 120184 151074 120224
rect 151074 120184 151114 120224
rect 151114 120184 151135 120224
rect 151217 120184 151238 120224
rect 151238 120184 151278 120224
rect 151278 120184 151303 120224
rect 151049 120161 151135 120184
rect 151217 120161 151303 120184
rect 74209 119468 74295 119491
rect 74377 119468 74463 119491
rect 74209 119428 74234 119468
rect 74234 119428 74274 119468
rect 74274 119428 74295 119468
rect 74377 119428 74398 119468
rect 74398 119428 74438 119468
rect 74438 119428 74463 119468
rect 74209 119405 74295 119428
rect 74377 119405 74463 119428
rect 89329 119468 89415 119491
rect 89497 119468 89583 119491
rect 89329 119428 89354 119468
rect 89354 119428 89394 119468
rect 89394 119428 89415 119468
rect 89497 119428 89518 119468
rect 89518 119428 89558 119468
rect 89558 119428 89583 119468
rect 89329 119405 89415 119428
rect 89497 119405 89583 119428
rect 104449 119468 104535 119491
rect 104617 119468 104703 119491
rect 104449 119428 104474 119468
rect 104474 119428 104514 119468
rect 104514 119428 104535 119468
rect 104617 119428 104638 119468
rect 104638 119428 104678 119468
rect 104678 119428 104703 119468
rect 104449 119405 104535 119428
rect 104617 119405 104703 119428
rect 119569 119468 119655 119491
rect 119737 119468 119823 119491
rect 119569 119428 119594 119468
rect 119594 119428 119634 119468
rect 119634 119428 119655 119468
rect 119737 119428 119758 119468
rect 119758 119428 119798 119468
rect 119798 119428 119823 119468
rect 119569 119405 119655 119428
rect 119737 119405 119823 119428
rect 134689 119468 134775 119491
rect 134857 119468 134943 119491
rect 134689 119428 134714 119468
rect 134714 119428 134754 119468
rect 134754 119428 134775 119468
rect 134857 119428 134878 119468
rect 134878 119428 134918 119468
rect 134918 119428 134943 119468
rect 134689 119405 134775 119428
rect 134857 119405 134943 119428
rect 149809 119468 149895 119491
rect 149977 119468 150063 119491
rect 149809 119428 149834 119468
rect 149834 119428 149874 119468
rect 149874 119428 149895 119468
rect 149977 119428 149998 119468
rect 149998 119428 150038 119468
rect 150038 119428 150063 119468
rect 149809 119405 149895 119428
rect 149977 119405 150063 119428
rect 75449 118712 75535 118735
rect 75617 118712 75703 118735
rect 75449 118672 75474 118712
rect 75474 118672 75514 118712
rect 75514 118672 75535 118712
rect 75617 118672 75638 118712
rect 75638 118672 75678 118712
rect 75678 118672 75703 118712
rect 75449 118649 75535 118672
rect 75617 118649 75703 118672
rect 90569 118712 90655 118735
rect 90737 118712 90823 118735
rect 90569 118672 90594 118712
rect 90594 118672 90634 118712
rect 90634 118672 90655 118712
rect 90737 118672 90758 118712
rect 90758 118672 90798 118712
rect 90798 118672 90823 118712
rect 90569 118649 90655 118672
rect 90737 118649 90823 118672
rect 105689 118712 105775 118735
rect 105857 118712 105943 118735
rect 105689 118672 105714 118712
rect 105714 118672 105754 118712
rect 105754 118672 105775 118712
rect 105857 118672 105878 118712
rect 105878 118672 105918 118712
rect 105918 118672 105943 118712
rect 105689 118649 105775 118672
rect 105857 118649 105943 118672
rect 120809 118712 120895 118735
rect 120977 118712 121063 118735
rect 120809 118672 120834 118712
rect 120834 118672 120874 118712
rect 120874 118672 120895 118712
rect 120977 118672 120998 118712
rect 120998 118672 121038 118712
rect 121038 118672 121063 118712
rect 120809 118649 120895 118672
rect 120977 118649 121063 118672
rect 135929 118712 136015 118735
rect 136097 118712 136183 118735
rect 135929 118672 135954 118712
rect 135954 118672 135994 118712
rect 135994 118672 136015 118712
rect 136097 118672 136118 118712
rect 136118 118672 136158 118712
rect 136158 118672 136183 118712
rect 135929 118649 136015 118672
rect 136097 118649 136183 118672
rect 151049 118712 151135 118735
rect 151217 118712 151303 118735
rect 151049 118672 151074 118712
rect 151074 118672 151114 118712
rect 151114 118672 151135 118712
rect 151217 118672 151238 118712
rect 151238 118672 151278 118712
rect 151278 118672 151303 118712
rect 151049 118649 151135 118672
rect 151217 118649 151303 118672
rect 74209 117956 74295 117979
rect 74377 117956 74463 117979
rect 74209 117916 74234 117956
rect 74234 117916 74274 117956
rect 74274 117916 74295 117956
rect 74377 117916 74398 117956
rect 74398 117916 74438 117956
rect 74438 117916 74463 117956
rect 74209 117893 74295 117916
rect 74377 117893 74463 117916
rect 89329 117956 89415 117979
rect 89497 117956 89583 117979
rect 89329 117916 89354 117956
rect 89354 117916 89394 117956
rect 89394 117916 89415 117956
rect 89497 117916 89518 117956
rect 89518 117916 89558 117956
rect 89558 117916 89583 117956
rect 89329 117893 89415 117916
rect 89497 117893 89583 117916
rect 104449 117956 104535 117979
rect 104617 117956 104703 117979
rect 104449 117916 104474 117956
rect 104474 117916 104514 117956
rect 104514 117916 104535 117956
rect 104617 117916 104638 117956
rect 104638 117916 104678 117956
rect 104678 117916 104703 117956
rect 104449 117893 104535 117916
rect 104617 117893 104703 117916
rect 119569 117956 119655 117979
rect 119737 117956 119823 117979
rect 119569 117916 119594 117956
rect 119594 117916 119634 117956
rect 119634 117916 119655 117956
rect 119737 117916 119758 117956
rect 119758 117916 119798 117956
rect 119798 117916 119823 117956
rect 119569 117893 119655 117916
rect 119737 117893 119823 117916
rect 134689 117956 134775 117979
rect 134857 117956 134943 117979
rect 134689 117916 134714 117956
rect 134714 117916 134754 117956
rect 134754 117916 134775 117956
rect 134857 117916 134878 117956
rect 134878 117916 134918 117956
rect 134918 117916 134943 117956
rect 134689 117893 134775 117916
rect 134857 117893 134943 117916
rect 149809 117956 149895 117979
rect 149977 117956 150063 117979
rect 149809 117916 149834 117956
rect 149834 117916 149874 117956
rect 149874 117916 149895 117956
rect 149977 117916 149998 117956
rect 149998 117916 150038 117956
rect 150038 117916 150063 117956
rect 149809 117893 149895 117916
rect 149977 117893 150063 117916
rect 75449 117200 75535 117223
rect 75617 117200 75703 117223
rect 75449 117160 75474 117200
rect 75474 117160 75514 117200
rect 75514 117160 75535 117200
rect 75617 117160 75638 117200
rect 75638 117160 75678 117200
rect 75678 117160 75703 117200
rect 75449 117137 75535 117160
rect 75617 117137 75703 117160
rect 90569 117200 90655 117223
rect 90737 117200 90823 117223
rect 90569 117160 90594 117200
rect 90594 117160 90634 117200
rect 90634 117160 90655 117200
rect 90737 117160 90758 117200
rect 90758 117160 90798 117200
rect 90798 117160 90823 117200
rect 90569 117137 90655 117160
rect 90737 117137 90823 117160
rect 105689 117200 105775 117223
rect 105857 117200 105943 117223
rect 105689 117160 105714 117200
rect 105714 117160 105754 117200
rect 105754 117160 105775 117200
rect 105857 117160 105878 117200
rect 105878 117160 105918 117200
rect 105918 117160 105943 117200
rect 105689 117137 105775 117160
rect 105857 117137 105943 117160
rect 120809 117200 120895 117223
rect 120977 117200 121063 117223
rect 120809 117160 120834 117200
rect 120834 117160 120874 117200
rect 120874 117160 120895 117200
rect 120977 117160 120998 117200
rect 120998 117160 121038 117200
rect 121038 117160 121063 117200
rect 120809 117137 120895 117160
rect 120977 117137 121063 117160
rect 135929 117200 136015 117223
rect 136097 117200 136183 117223
rect 135929 117160 135954 117200
rect 135954 117160 135994 117200
rect 135994 117160 136015 117200
rect 136097 117160 136118 117200
rect 136118 117160 136158 117200
rect 136158 117160 136183 117200
rect 135929 117137 136015 117160
rect 136097 117137 136183 117160
rect 151049 117200 151135 117223
rect 151217 117200 151303 117223
rect 151049 117160 151074 117200
rect 151074 117160 151114 117200
rect 151114 117160 151135 117200
rect 151217 117160 151238 117200
rect 151238 117160 151278 117200
rect 151278 117160 151303 117200
rect 151049 117137 151135 117160
rect 151217 117137 151303 117160
rect 74209 116444 74295 116467
rect 74377 116444 74463 116467
rect 74209 116404 74234 116444
rect 74234 116404 74274 116444
rect 74274 116404 74295 116444
rect 74377 116404 74398 116444
rect 74398 116404 74438 116444
rect 74438 116404 74463 116444
rect 74209 116381 74295 116404
rect 74377 116381 74463 116404
rect 89329 116444 89415 116467
rect 89497 116444 89583 116467
rect 89329 116404 89354 116444
rect 89354 116404 89394 116444
rect 89394 116404 89415 116444
rect 89497 116404 89518 116444
rect 89518 116404 89558 116444
rect 89558 116404 89583 116444
rect 89329 116381 89415 116404
rect 89497 116381 89583 116404
rect 104449 116444 104535 116467
rect 104617 116444 104703 116467
rect 104449 116404 104474 116444
rect 104474 116404 104514 116444
rect 104514 116404 104535 116444
rect 104617 116404 104638 116444
rect 104638 116404 104678 116444
rect 104678 116404 104703 116444
rect 104449 116381 104535 116404
rect 104617 116381 104703 116404
rect 119569 116444 119655 116467
rect 119737 116444 119823 116467
rect 119569 116404 119594 116444
rect 119594 116404 119634 116444
rect 119634 116404 119655 116444
rect 119737 116404 119758 116444
rect 119758 116404 119798 116444
rect 119798 116404 119823 116444
rect 119569 116381 119655 116404
rect 119737 116381 119823 116404
rect 134689 116444 134775 116467
rect 134857 116444 134943 116467
rect 134689 116404 134714 116444
rect 134714 116404 134754 116444
rect 134754 116404 134775 116444
rect 134857 116404 134878 116444
rect 134878 116404 134918 116444
rect 134918 116404 134943 116444
rect 134689 116381 134775 116404
rect 134857 116381 134943 116404
rect 149809 116444 149895 116467
rect 149977 116444 150063 116467
rect 149809 116404 149834 116444
rect 149834 116404 149874 116444
rect 149874 116404 149895 116444
rect 149977 116404 149998 116444
rect 149998 116404 150038 116444
rect 150038 116404 150063 116444
rect 149809 116381 149895 116404
rect 149977 116381 150063 116404
rect 75449 115688 75535 115711
rect 75617 115688 75703 115711
rect 75449 115648 75474 115688
rect 75474 115648 75514 115688
rect 75514 115648 75535 115688
rect 75617 115648 75638 115688
rect 75638 115648 75678 115688
rect 75678 115648 75703 115688
rect 75449 115625 75535 115648
rect 75617 115625 75703 115648
rect 90569 115688 90655 115711
rect 90737 115688 90823 115711
rect 90569 115648 90594 115688
rect 90594 115648 90634 115688
rect 90634 115648 90655 115688
rect 90737 115648 90758 115688
rect 90758 115648 90798 115688
rect 90798 115648 90823 115688
rect 90569 115625 90655 115648
rect 90737 115625 90823 115648
rect 105689 115688 105775 115711
rect 105857 115688 105943 115711
rect 105689 115648 105714 115688
rect 105714 115648 105754 115688
rect 105754 115648 105775 115688
rect 105857 115648 105878 115688
rect 105878 115648 105918 115688
rect 105918 115648 105943 115688
rect 105689 115625 105775 115648
rect 105857 115625 105943 115648
rect 120809 115688 120895 115711
rect 120977 115688 121063 115711
rect 120809 115648 120834 115688
rect 120834 115648 120874 115688
rect 120874 115648 120895 115688
rect 120977 115648 120998 115688
rect 120998 115648 121038 115688
rect 121038 115648 121063 115688
rect 120809 115625 120895 115648
rect 120977 115625 121063 115648
rect 135929 115688 136015 115711
rect 136097 115688 136183 115711
rect 135929 115648 135954 115688
rect 135954 115648 135994 115688
rect 135994 115648 136015 115688
rect 136097 115648 136118 115688
rect 136118 115648 136158 115688
rect 136158 115648 136183 115688
rect 135929 115625 136015 115648
rect 136097 115625 136183 115648
rect 151049 115688 151135 115711
rect 151217 115688 151303 115711
rect 151049 115648 151074 115688
rect 151074 115648 151114 115688
rect 151114 115648 151135 115688
rect 151217 115648 151238 115688
rect 151238 115648 151278 115688
rect 151278 115648 151303 115688
rect 151049 115625 151135 115648
rect 151217 115625 151303 115648
rect 74209 114932 74295 114955
rect 74377 114932 74463 114955
rect 74209 114892 74234 114932
rect 74234 114892 74274 114932
rect 74274 114892 74295 114932
rect 74377 114892 74398 114932
rect 74398 114892 74438 114932
rect 74438 114892 74463 114932
rect 74209 114869 74295 114892
rect 74377 114869 74463 114892
rect 89329 114932 89415 114955
rect 89497 114932 89583 114955
rect 89329 114892 89354 114932
rect 89354 114892 89394 114932
rect 89394 114892 89415 114932
rect 89497 114892 89518 114932
rect 89518 114892 89558 114932
rect 89558 114892 89583 114932
rect 89329 114869 89415 114892
rect 89497 114869 89583 114892
rect 104449 114932 104535 114955
rect 104617 114932 104703 114955
rect 104449 114892 104474 114932
rect 104474 114892 104514 114932
rect 104514 114892 104535 114932
rect 104617 114892 104638 114932
rect 104638 114892 104678 114932
rect 104678 114892 104703 114932
rect 104449 114869 104535 114892
rect 104617 114869 104703 114892
rect 119569 114932 119655 114955
rect 119737 114932 119823 114955
rect 119569 114892 119594 114932
rect 119594 114892 119634 114932
rect 119634 114892 119655 114932
rect 119737 114892 119758 114932
rect 119758 114892 119798 114932
rect 119798 114892 119823 114932
rect 119569 114869 119655 114892
rect 119737 114869 119823 114892
rect 134689 114932 134775 114955
rect 134857 114932 134943 114955
rect 134689 114892 134714 114932
rect 134714 114892 134754 114932
rect 134754 114892 134775 114932
rect 134857 114892 134878 114932
rect 134878 114892 134918 114932
rect 134918 114892 134943 114932
rect 134689 114869 134775 114892
rect 134857 114869 134943 114892
rect 149809 114932 149895 114955
rect 149977 114932 150063 114955
rect 149809 114892 149834 114932
rect 149834 114892 149874 114932
rect 149874 114892 149895 114932
rect 149977 114892 149998 114932
rect 149998 114892 150038 114932
rect 150038 114892 150063 114932
rect 149809 114869 149895 114892
rect 149977 114869 150063 114892
rect 75449 114176 75535 114199
rect 75617 114176 75703 114199
rect 75449 114136 75474 114176
rect 75474 114136 75514 114176
rect 75514 114136 75535 114176
rect 75617 114136 75638 114176
rect 75638 114136 75678 114176
rect 75678 114136 75703 114176
rect 75449 114113 75535 114136
rect 75617 114113 75703 114136
rect 90569 114176 90655 114199
rect 90737 114176 90823 114199
rect 90569 114136 90594 114176
rect 90594 114136 90634 114176
rect 90634 114136 90655 114176
rect 90737 114136 90758 114176
rect 90758 114136 90798 114176
rect 90798 114136 90823 114176
rect 90569 114113 90655 114136
rect 90737 114113 90823 114136
rect 105689 114176 105775 114199
rect 105857 114176 105943 114199
rect 105689 114136 105714 114176
rect 105714 114136 105754 114176
rect 105754 114136 105775 114176
rect 105857 114136 105878 114176
rect 105878 114136 105918 114176
rect 105918 114136 105943 114176
rect 105689 114113 105775 114136
rect 105857 114113 105943 114136
rect 120809 114176 120895 114199
rect 120977 114176 121063 114199
rect 120809 114136 120834 114176
rect 120834 114136 120874 114176
rect 120874 114136 120895 114176
rect 120977 114136 120998 114176
rect 120998 114136 121038 114176
rect 121038 114136 121063 114176
rect 120809 114113 120895 114136
rect 120977 114113 121063 114136
rect 135929 114176 136015 114199
rect 136097 114176 136183 114199
rect 135929 114136 135954 114176
rect 135954 114136 135994 114176
rect 135994 114136 136015 114176
rect 136097 114136 136118 114176
rect 136118 114136 136158 114176
rect 136158 114136 136183 114176
rect 135929 114113 136015 114136
rect 136097 114113 136183 114136
rect 151049 114176 151135 114199
rect 151217 114176 151303 114199
rect 151049 114136 151074 114176
rect 151074 114136 151114 114176
rect 151114 114136 151135 114176
rect 151217 114136 151238 114176
rect 151238 114136 151278 114176
rect 151278 114136 151303 114176
rect 151049 114113 151135 114136
rect 151217 114113 151303 114136
rect 74209 113420 74295 113443
rect 74377 113420 74463 113443
rect 74209 113380 74234 113420
rect 74234 113380 74274 113420
rect 74274 113380 74295 113420
rect 74377 113380 74398 113420
rect 74398 113380 74438 113420
rect 74438 113380 74463 113420
rect 74209 113357 74295 113380
rect 74377 113357 74463 113380
rect 89329 113420 89415 113443
rect 89497 113420 89583 113443
rect 89329 113380 89354 113420
rect 89354 113380 89394 113420
rect 89394 113380 89415 113420
rect 89497 113380 89518 113420
rect 89518 113380 89558 113420
rect 89558 113380 89583 113420
rect 89329 113357 89415 113380
rect 89497 113357 89583 113380
rect 104449 113420 104535 113443
rect 104617 113420 104703 113443
rect 104449 113380 104474 113420
rect 104474 113380 104514 113420
rect 104514 113380 104535 113420
rect 104617 113380 104638 113420
rect 104638 113380 104678 113420
rect 104678 113380 104703 113420
rect 104449 113357 104535 113380
rect 104617 113357 104703 113380
rect 119569 113420 119655 113443
rect 119737 113420 119823 113443
rect 119569 113380 119594 113420
rect 119594 113380 119634 113420
rect 119634 113380 119655 113420
rect 119737 113380 119758 113420
rect 119758 113380 119798 113420
rect 119798 113380 119823 113420
rect 119569 113357 119655 113380
rect 119737 113357 119823 113380
rect 134689 113420 134775 113443
rect 134857 113420 134943 113443
rect 134689 113380 134714 113420
rect 134714 113380 134754 113420
rect 134754 113380 134775 113420
rect 134857 113380 134878 113420
rect 134878 113380 134918 113420
rect 134918 113380 134943 113420
rect 134689 113357 134775 113380
rect 134857 113357 134943 113380
rect 149809 113420 149895 113443
rect 149977 113420 150063 113443
rect 149809 113380 149834 113420
rect 149834 113380 149874 113420
rect 149874 113380 149895 113420
rect 149977 113380 149998 113420
rect 149998 113380 150038 113420
rect 150038 113380 150063 113420
rect 149809 113357 149895 113380
rect 149977 113357 150063 113380
rect 75449 112664 75535 112687
rect 75617 112664 75703 112687
rect 75449 112624 75474 112664
rect 75474 112624 75514 112664
rect 75514 112624 75535 112664
rect 75617 112624 75638 112664
rect 75638 112624 75678 112664
rect 75678 112624 75703 112664
rect 75449 112601 75535 112624
rect 75617 112601 75703 112624
rect 90569 112664 90655 112687
rect 90737 112664 90823 112687
rect 90569 112624 90594 112664
rect 90594 112624 90634 112664
rect 90634 112624 90655 112664
rect 90737 112624 90758 112664
rect 90758 112624 90798 112664
rect 90798 112624 90823 112664
rect 90569 112601 90655 112624
rect 90737 112601 90823 112624
rect 105689 112664 105775 112687
rect 105857 112664 105943 112687
rect 105689 112624 105714 112664
rect 105714 112624 105754 112664
rect 105754 112624 105775 112664
rect 105857 112624 105878 112664
rect 105878 112624 105918 112664
rect 105918 112624 105943 112664
rect 105689 112601 105775 112624
rect 105857 112601 105943 112624
rect 120809 112664 120895 112687
rect 120977 112664 121063 112687
rect 120809 112624 120834 112664
rect 120834 112624 120874 112664
rect 120874 112624 120895 112664
rect 120977 112624 120998 112664
rect 120998 112624 121038 112664
rect 121038 112624 121063 112664
rect 120809 112601 120895 112624
rect 120977 112601 121063 112624
rect 135929 112664 136015 112687
rect 136097 112664 136183 112687
rect 135929 112624 135954 112664
rect 135954 112624 135994 112664
rect 135994 112624 136015 112664
rect 136097 112624 136118 112664
rect 136118 112624 136158 112664
rect 136158 112624 136183 112664
rect 135929 112601 136015 112624
rect 136097 112601 136183 112624
rect 151049 112664 151135 112687
rect 151217 112664 151303 112687
rect 151049 112624 151074 112664
rect 151074 112624 151114 112664
rect 151114 112624 151135 112664
rect 151217 112624 151238 112664
rect 151238 112624 151278 112664
rect 151278 112624 151303 112664
rect 151049 112601 151135 112624
rect 151217 112601 151303 112624
rect 74209 111908 74295 111931
rect 74377 111908 74463 111931
rect 74209 111868 74234 111908
rect 74234 111868 74274 111908
rect 74274 111868 74295 111908
rect 74377 111868 74398 111908
rect 74398 111868 74438 111908
rect 74438 111868 74463 111908
rect 74209 111845 74295 111868
rect 74377 111845 74463 111868
rect 89329 111908 89415 111931
rect 89497 111908 89583 111931
rect 89329 111868 89354 111908
rect 89354 111868 89394 111908
rect 89394 111868 89415 111908
rect 89497 111868 89518 111908
rect 89518 111868 89558 111908
rect 89558 111868 89583 111908
rect 89329 111845 89415 111868
rect 89497 111845 89583 111868
rect 104449 111908 104535 111931
rect 104617 111908 104703 111931
rect 104449 111868 104474 111908
rect 104474 111868 104514 111908
rect 104514 111868 104535 111908
rect 104617 111868 104638 111908
rect 104638 111868 104678 111908
rect 104678 111868 104703 111908
rect 104449 111845 104535 111868
rect 104617 111845 104703 111868
rect 119569 111908 119655 111931
rect 119737 111908 119823 111931
rect 119569 111868 119594 111908
rect 119594 111868 119634 111908
rect 119634 111868 119655 111908
rect 119737 111868 119758 111908
rect 119758 111868 119798 111908
rect 119798 111868 119823 111908
rect 119569 111845 119655 111868
rect 119737 111845 119823 111868
rect 134689 111908 134775 111931
rect 134857 111908 134943 111931
rect 134689 111868 134714 111908
rect 134714 111868 134754 111908
rect 134754 111868 134775 111908
rect 134857 111868 134878 111908
rect 134878 111868 134918 111908
rect 134918 111868 134943 111908
rect 134689 111845 134775 111868
rect 134857 111845 134943 111868
rect 149809 111908 149895 111931
rect 149977 111908 150063 111931
rect 149809 111868 149834 111908
rect 149834 111868 149874 111908
rect 149874 111868 149895 111908
rect 149977 111868 149998 111908
rect 149998 111868 150038 111908
rect 150038 111868 150063 111908
rect 149809 111845 149895 111868
rect 149977 111845 150063 111868
rect 75449 111152 75535 111175
rect 75617 111152 75703 111175
rect 75449 111112 75474 111152
rect 75474 111112 75514 111152
rect 75514 111112 75535 111152
rect 75617 111112 75638 111152
rect 75638 111112 75678 111152
rect 75678 111112 75703 111152
rect 75449 111089 75535 111112
rect 75617 111089 75703 111112
rect 90569 111152 90655 111175
rect 90737 111152 90823 111175
rect 90569 111112 90594 111152
rect 90594 111112 90634 111152
rect 90634 111112 90655 111152
rect 90737 111112 90758 111152
rect 90758 111112 90798 111152
rect 90798 111112 90823 111152
rect 90569 111089 90655 111112
rect 90737 111089 90823 111112
rect 105689 111152 105775 111175
rect 105857 111152 105943 111175
rect 105689 111112 105714 111152
rect 105714 111112 105754 111152
rect 105754 111112 105775 111152
rect 105857 111112 105878 111152
rect 105878 111112 105918 111152
rect 105918 111112 105943 111152
rect 105689 111089 105775 111112
rect 105857 111089 105943 111112
rect 120809 111152 120895 111175
rect 120977 111152 121063 111175
rect 120809 111112 120834 111152
rect 120834 111112 120874 111152
rect 120874 111112 120895 111152
rect 120977 111112 120998 111152
rect 120998 111112 121038 111152
rect 121038 111112 121063 111152
rect 120809 111089 120895 111112
rect 120977 111089 121063 111112
rect 135929 111152 136015 111175
rect 136097 111152 136183 111175
rect 135929 111112 135954 111152
rect 135954 111112 135994 111152
rect 135994 111112 136015 111152
rect 136097 111112 136118 111152
rect 136118 111112 136158 111152
rect 136158 111112 136183 111152
rect 135929 111089 136015 111112
rect 136097 111089 136183 111112
rect 151049 111152 151135 111175
rect 151217 111152 151303 111175
rect 151049 111112 151074 111152
rect 151074 111112 151114 111152
rect 151114 111112 151135 111152
rect 151217 111112 151238 111152
rect 151238 111112 151278 111152
rect 151278 111112 151303 111152
rect 151049 111089 151135 111112
rect 151217 111089 151303 111112
rect 74209 110396 74295 110419
rect 74377 110396 74463 110419
rect 74209 110356 74234 110396
rect 74234 110356 74274 110396
rect 74274 110356 74295 110396
rect 74377 110356 74398 110396
rect 74398 110356 74438 110396
rect 74438 110356 74463 110396
rect 74209 110333 74295 110356
rect 74377 110333 74463 110356
rect 89329 110396 89415 110419
rect 89497 110396 89583 110419
rect 89329 110356 89354 110396
rect 89354 110356 89394 110396
rect 89394 110356 89415 110396
rect 89497 110356 89518 110396
rect 89518 110356 89558 110396
rect 89558 110356 89583 110396
rect 89329 110333 89415 110356
rect 89497 110333 89583 110356
rect 104449 110396 104535 110419
rect 104617 110396 104703 110419
rect 104449 110356 104474 110396
rect 104474 110356 104514 110396
rect 104514 110356 104535 110396
rect 104617 110356 104638 110396
rect 104638 110356 104678 110396
rect 104678 110356 104703 110396
rect 104449 110333 104535 110356
rect 104617 110333 104703 110356
rect 119569 110396 119655 110419
rect 119737 110396 119823 110419
rect 119569 110356 119594 110396
rect 119594 110356 119634 110396
rect 119634 110356 119655 110396
rect 119737 110356 119758 110396
rect 119758 110356 119798 110396
rect 119798 110356 119823 110396
rect 119569 110333 119655 110356
rect 119737 110333 119823 110356
rect 134689 110396 134775 110419
rect 134857 110396 134943 110419
rect 134689 110356 134714 110396
rect 134714 110356 134754 110396
rect 134754 110356 134775 110396
rect 134857 110356 134878 110396
rect 134878 110356 134918 110396
rect 134918 110356 134943 110396
rect 134689 110333 134775 110356
rect 134857 110333 134943 110356
rect 149809 110396 149895 110419
rect 149977 110396 150063 110419
rect 149809 110356 149834 110396
rect 149834 110356 149874 110396
rect 149874 110356 149895 110396
rect 149977 110356 149998 110396
rect 149998 110356 150038 110396
rect 150038 110356 150063 110396
rect 149809 110333 149895 110356
rect 149977 110333 150063 110356
rect 75449 109640 75535 109663
rect 75617 109640 75703 109663
rect 75449 109600 75474 109640
rect 75474 109600 75514 109640
rect 75514 109600 75535 109640
rect 75617 109600 75638 109640
rect 75638 109600 75678 109640
rect 75678 109600 75703 109640
rect 75449 109577 75535 109600
rect 75617 109577 75703 109600
rect 90569 109640 90655 109663
rect 90737 109640 90823 109663
rect 90569 109600 90594 109640
rect 90594 109600 90634 109640
rect 90634 109600 90655 109640
rect 90737 109600 90758 109640
rect 90758 109600 90798 109640
rect 90798 109600 90823 109640
rect 90569 109577 90655 109600
rect 90737 109577 90823 109600
rect 105689 109640 105775 109663
rect 105857 109640 105943 109663
rect 105689 109600 105714 109640
rect 105714 109600 105754 109640
rect 105754 109600 105775 109640
rect 105857 109600 105878 109640
rect 105878 109600 105918 109640
rect 105918 109600 105943 109640
rect 105689 109577 105775 109600
rect 105857 109577 105943 109600
rect 120809 109640 120895 109663
rect 120977 109640 121063 109663
rect 120809 109600 120834 109640
rect 120834 109600 120874 109640
rect 120874 109600 120895 109640
rect 120977 109600 120998 109640
rect 120998 109600 121038 109640
rect 121038 109600 121063 109640
rect 120809 109577 120895 109600
rect 120977 109577 121063 109600
rect 135929 109640 136015 109663
rect 136097 109640 136183 109663
rect 135929 109600 135954 109640
rect 135954 109600 135994 109640
rect 135994 109600 136015 109640
rect 136097 109600 136118 109640
rect 136118 109600 136158 109640
rect 136158 109600 136183 109640
rect 135929 109577 136015 109600
rect 136097 109577 136183 109600
rect 151049 109640 151135 109663
rect 151217 109640 151303 109663
rect 151049 109600 151074 109640
rect 151074 109600 151114 109640
rect 151114 109600 151135 109640
rect 151217 109600 151238 109640
rect 151238 109600 151278 109640
rect 151278 109600 151303 109640
rect 151049 109577 151135 109600
rect 151217 109577 151303 109600
rect 74209 108884 74295 108907
rect 74377 108884 74463 108907
rect 74209 108844 74234 108884
rect 74234 108844 74274 108884
rect 74274 108844 74295 108884
rect 74377 108844 74398 108884
rect 74398 108844 74438 108884
rect 74438 108844 74463 108884
rect 74209 108821 74295 108844
rect 74377 108821 74463 108844
rect 89329 108884 89415 108907
rect 89497 108884 89583 108907
rect 89329 108844 89354 108884
rect 89354 108844 89394 108884
rect 89394 108844 89415 108884
rect 89497 108844 89518 108884
rect 89518 108844 89558 108884
rect 89558 108844 89583 108884
rect 89329 108821 89415 108844
rect 89497 108821 89583 108844
rect 104449 108884 104535 108907
rect 104617 108884 104703 108907
rect 104449 108844 104474 108884
rect 104474 108844 104514 108884
rect 104514 108844 104535 108884
rect 104617 108844 104638 108884
rect 104638 108844 104678 108884
rect 104678 108844 104703 108884
rect 104449 108821 104535 108844
rect 104617 108821 104703 108844
rect 119569 108884 119655 108907
rect 119737 108884 119823 108907
rect 119569 108844 119594 108884
rect 119594 108844 119634 108884
rect 119634 108844 119655 108884
rect 119737 108844 119758 108884
rect 119758 108844 119798 108884
rect 119798 108844 119823 108884
rect 119569 108821 119655 108844
rect 119737 108821 119823 108844
rect 134689 108884 134775 108907
rect 134857 108884 134943 108907
rect 134689 108844 134714 108884
rect 134714 108844 134754 108884
rect 134754 108844 134775 108884
rect 134857 108844 134878 108884
rect 134878 108844 134918 108884
rect 134918 108844 134943 108884
rect 134689 108821 134775 108844
rect 134857 108821 134943 108844
rect 149809 108884 149895 108907
rect 149977 108884 150063 108907
rect 149809 108844 149834 108884
rect 149834 108844 149874 108884
rect 149874 108844 149895 108884
rect 149977 108844 149998 108884
rect 149998 108844 150038 108884
rect 150038 108844 150063 108884
rect 149809 108821 149895 108844
rect 149977 108821 150063 108844
rect 75449 108128 75535 108151
rect 75617 108128 75703 108151
rect 75449 108088 75474 108128
rect 75474 108088 75514 108128
rect 75514 108088 75535 108128
rect 75617 108088 75638 108128
rect 75638 108088 75678 108128
rect 75678 108088 75703 108128
rect 75449 108065 75535 108088
rect 75617 108065 75703 108088
rect 90569 108128 90655 108151
rect 90737 108128 90823 108151
rect 90569 108088 90594 108128
rect 90594 108088 90634 108128
rect 90634 108088 90655 108128
rect 90737 108088 90758 108128
rect 90758 108088 90798 108128
rect 90798 108088 90823 108128
rect 90569 108065 90655 108088
rect 90737 108065 90823 108088
rect 105689 108128 105775 108151
rect 105857 108128 105943 108151
rect 105689 108088 105714 108128
rect 105714 108088 105754 108128
rect 105754 108088 105775 108128
rect 105857 108088 105878 108128
rect 105878 108088 105918 108128
rect 105918 108088 105943 108128
rect 105689 108065 105775 108088
rect 105857 108065 105943 108088
rect 120809 108128 120895 108151
rect 120977 108128 121063 108151
rect 120809 108088 120834 108128
rect 120834 108088 120874 108128
rect 120874 108088 120895 108128
rect 120977 108088 120998 108128
rect 120998 108088 121038 108128
rect 121038 108088 121063 108128
rect 120809 108065 120895 108088
rect 120977 108065 121063 108088
rect 135929 108128 136015 108151
rect 136097 108128 136183 108151
rect 135929 108088 135954 108128
rect 135954 108088 135994 108128
rect 135994 108088 136015 108128
rect 136097 108088 136118 108128
rect 136118 108088 136158 108128
rect 136158 108088 136183 108128
rect 135929 108065 136015 108088
rect 136097 108065 136183 108088
rect 151049 108128 151135 108151
rect 151217 108128 151303 108151
rect 151049 108088 151074 108128
rect 151074 108088 151114 108128
rect 151114 108088 151135 108128
rect 151217 108088 151238 108128
rect 151238 108088 151278 108128
rect 151278 108088 151303 108128
rect 151049 108065 151135 108088
rect 151217 108065 151303 108088
rect 74209 107372 74295 107395
rect 74377 107372 74463 107395
rect 74209 107332 74234 107372
rect 74234 107332 74274 107372
rect 74274 107332 74295 107372
rect 74377 107332 74398 107372
rect 74398 107332 74438 107372
rect 74438 107332 74463 107372
rect 74209 107309 74295 107332
rect 74377 107309 74463 107332
rect 89329 107372 89415 107395
rect 89497 107372 89583 107395
rect 89329 107332 89354 107372
rect 89354 107332 89394 107372
rect 89394 107332 89415 107372
rect 89497 107332 89518 107372
rect 89518 107332 89558 107372
rect 89558 107332 89583 107372
rect 89329 107309 89415 107332
rect 89497 107309 89583 107332
rect 104449 107372 104535 107395
rect 104617 107372 104703 107395
rect 104449 107332 104474 107372
rect 104474 107332 104514 107372
rect 104514 107332 104535 107372
rect 104617 107332 104638 107372
rect 104638 107332 104678 107372
rect 104678 107332 104703 107372
rect 104449 107309 104535 107332
rect 104617 107309 104703 107332
rect 119569 107372 119655 107395
rect 119737 107372 119823 107395
rect 119569 107332 119594 107372
rect 119594 107332 119634 107372
rect 119634 107332 119655 107372
rect 119737 107332 119758 107372
rect 119758 107332 119798 107372
rect 119798 107332 119823 107372
rect 119569 107309 119655 107332
rect 119737 107309 119823 107332
rect 134689 107372 134775 107395
rect 134857 107372 134943 107395
rect 134689 107332 134714 107372
rect 134714 107332 134754 107372
rect 134754 107332 134775 107372
rect 134857 107332 134878 107372
rect 134878 107332 134918 107372
rect 134918 107332 134943 107372
rect 134689 107309 134775 107332
rect 134857 107309 134943 107332
rect 149809 107372 149895 107395
rect 149977 107372 150063 107395
rect 149809 107332 149834 107372
rect 149834 107332 149874 107372
rect 149874 107332 149895 107372
rect 149977 107332 149998 107372
rect 149998 107332 150038 107372
rect 150038 107332 150063 107372
rect 149809 107309 149895 107332
rect 149977 107309 150063 107332
rect 75449 106616 75535 106639
rect 75617 106616 75703 106639
rect 75449 106576 75474 106616
rect 75474 106576 75514 106616
rect 75514 106576 75535 106616
rect 75617 106576 75638 106616
rect 75638 106576 75678 106616
rect 75678 106576 75703 106616
rect 75449 106553 75535 106576
rect 75617 106553 75703 106576
rect 90569 106616 90655 106639
rect 90737 106616 90823 106639
rect 90569 106576 90594 106616
rect 90594 106576 90634 106616
rect 90634 106576 90655 106616
rect 90737 106576 90758 106616
rect 90758 106576 90798 106616
rect 90798 106576 90823 106616
rect 90569 106553 90655 106576
rect 90737 106553 90823 106576
rect 105689 106616 105775 106639
rect 105857 106616 105943 106639
rect 105689 106576 105714 106616
rect 105714 106576 105754 106616
rect 105754 106576 105775 106616
rect 105857 106576 105878 106616
rect 105878 106576 105918 106616
rect 105918 106576 105943 106616
rect 105689 106553 105775 106576
rect 105857 106553 105943 106576
rect 120809 106616 120895 106639
rect 120977 106616 121063 106639
rect 120809 106576 120834 106616
rect 120834 106576 120874 106616
rect 120874 106576 120895 106616
rect 120977 106576 120998 106616
rect 120998 106576 121038 106616
rect 121038 106576 121063 106616
rect 120809 106553 120895 106576
rect 120977 106553 121063 106576
rect 135929 106616 136015 106639
rect 136097 106616 136183 106639
rect 135929 106576 135954 106616
rect 135954 106576 135994 106616
rect 135994 106576 136015 106616
rect 136097 106576 136118 106616
rect 136118 106576 136158 106616
rect 136158 106576 136183 106616
rect 135929 106553 136015 106576
rect 136097 106553 136183 106576
rect 151049 106616 151135 106639
rect 151217 106616 151303 106639
rect 151049 106576 151074 106616
rect 151074 106576 151114 106616
rect 151114 106576 151135 106616
rect 151217 106576 151238 106616
rect 151238 106576 151278 106616
rect 151278 106576 151303 106616
rect 151049 106553 151135 106576
rect 151217 106553 151303 106576
rect 74209 105860 74295 105883
rect 74377 105860 74463 105883
rect 74209 105820 74234 105860
rect 74234 105820 74274 105860
rect 74274 105820 74295 105860
rect 74377 105820 74398 105860
rect 74398 105820 74438 105860
rect 74438 105820 74463 105860
rect 74209 105797 74295 105820
rect 74377 105797 74463 105820
rect 89329 105860 89415 105883
rect 89497 105860 89583 105883
rect 89329 105820 89354 105860
rect 89354 105820 89394 105860
rect 89394 105820 89415 105860
rect 89497 105820 89518 105860
rect 89518 105820 89558 105860
rect 89558 105820 89583 105860
rect 89329 105797 89415 105820
rect 89497 105797 89583 105820
rect 104449 105860 104535 105883
rect 104617 105860 104703 105883
rect 104449 105820 104474 105860
rect 104474 105820 104514 105860
rect 104514 105820 104535 105860
rect 104617 105820 104638 105860
rect 104638 105820 104678 105860
rect 104678 105820 104703 105860
rect 104449 105797 104535 105820
rect 104617 105797 104703 105820
rect 119569 105860 119655 105883
rect 119737 105860 119823 105883
rect 119569 105820 119594 105860
rect 119594 105820 119634 105860
rect 119634 105820 119655 105860
rect 119737 105820 119758 105860
rect 119758 105820 119798 105860
rect 119798 105820 119823 105860
rect 119569 105797 119655 105820
rect 119737 105797 119823 105820
rect 134689 105860 134775 105883
rect 134857 105860 134943 105883
rect 134689 105820 134714 105860
rect 134714 105820 134754 105860
rect 134754 105820 134775 105860
rect 134857 105820 134878 105860
rect 134878 105820 134918 105860
rect 134918 105820 134943 105860
rect 134689 105797 134775 105820
rect 134857 105797 134943 105820
rect 149809 105860 149895 105883
rect 149977 105860 150063 105883
rect 149809 105820 149834 105860
rect 149834 105820 149874 105860
rect 149874 105820 149895 105860
rect 149977 105820 149998 105860
rect 149998 105820 150038 105860
rect 150038 105820 150063 105860
rect 149809 105797 149895 105820
rect 149977 105797 150063 105820
rect 75449 105104 75535 105127
rect 75617 105104 75703 105127
rect 75449 105064 75474 105104
rect 75474 105064 75514 105104
rect 75514 105064 75535 105104
rect 75617 105064 75638 105104
rect 75638 105064 75678 105104
rect 75678 105064 75703 105104
rect 75449 105041 75535 105064
rect 75617 105041 75703 105064
rect 90569 105104 90655 105127
rect 90737 105104 90823 105127
rect 90569 105064 90594 105104
rect 90594 105064 90634 105104
rect 90634 105064 90655 105104
rect 90737 105064 90758 105104
rect 90758 105064 90798 105104
rect 90798 105064 90823 105104
rect 90569 105041 90655 105064
rect 90737 105041 90823 105064
rect 105689 105104 105775 105127
rect 105857 105104 105943 105127
rect 105689 105064 105714 105104
rect 105714 105064 105754 105104
rect 105754 105064 105775 105104
rect 105857 105064 105878 105104
rect 105878 105064 105918 105104
rect 105918 105064 105943 105104
rect 105689 105041 105775 105064
rect 105857 105041 105943 105064
rect 120809 105104 120895 105127
rect 120977 105104 121063 105127
rect 120809 105064 120834 105104
rect 120834 105064 120874 105104
rect 120874 105064 120895 105104
rect 120977 105064 120998 105104
rect 120998 105064 121038 105104
rect 121038 105064 121063 105104
rect 120809 105041 120895 105064
rect 120977 105041 121063 105064
rect 135929 105104 136015 105127
rect 136097 105104 136183 105127
rect 135929 105064 135954 105104
rect 135954 105064 135994 105104
rect 135994 105064 136015 105104
rect 136097 105064 136118 105104
rect 136118 105064 136158 105104
rect 136158 105064 136183 105104
rect 135929 105041 136015 105064
rect 136097 105041 136183 105064
rect 151049 105104 151135 105127
rect 151217 105104 151303 105127
rect 151049 105064 151074 105104
rect 151074 105064 151114 105104
rect 151114 105064 151135 105104
rect 151217 105064 151238 105104
rect 151238 105064 151278 105104
rect 151278 105064 151303 105104
rect 151049 105041 151135 105064
rect 151217 105041 151303 105064
rect 74209 104348 74295 104371
rect 74377 104348 74463 104371
rect 74209 104308 74234 104348
rect 74234 104308 74274 104348
rect 74274 104308 74295 104348
rect 74377 104308 74398 104348
rect 74398 104308 74438 104348
rect 74438 104308 74463 104348
rect 74209 104285 74295 104308
rect 74377 104285 74463 104308
rect 89329 104348 89415 104371
rect 89497 104348 89583 104371
rect 89329 104308 89354 104348
rect 89354 104308 89394 104348
rect 89394 104308 89415 104348
rect 89497 104308 89518 104348
rect 89518 104308 89558 104348
rect 89558 104308 89583 104348
rect 89329 104285 89415 104308
rect 89497 104285 89583 104308
rect 104449 104348 104535 104371
rect 104617 104348 104703 104371
rect 104449 104308 104474 104348
rect 104474 104308 104514 104348
rect 104514 104308 104535 104348
rect 104617 104308 104638 104348
rect 104638 104308 104678 104348
rect 104678 104308 104703 104348
rect 104449 104285 104535 104308
rect 104617 104285 104703 104308
rect 119569 104348 119655 104371
rect 119737 104348 119823 104371
rect 119569 104308 119594 104348
rect 119594 104308 119634 104348
rect 119634 104308 119655 104348
rect 119737 104308 119758 104348
rect 119758 104308 119798 104348
rect 119798 104308 119823 104348
rect 119569 104285 119655 104308
rect 119737 104285 119823 104308
rect 134689 104348 134775 104371
rect 134857 104348 134943 104371
rect 134689 104308 134714 104348
rect 134714 104308 134754 104348
rect 134754 104308 134775 104348
rect 134857 104308 134878 104348
rect 134878 104308 134918 104348
rect 134918 104308 134943 104348
rect 134689 104285 134775 104308
rect 134857 104285 134943 104308
rect 149809 104348 149895 104371
rect 149977 104348 150063 104371
rect 149809 104308 149834 104348
rect 149834 104308 149874 104348
rect 149874 104308 149895 104348
rect 149977 104308 149998 104348
rect 149998 104308 150038 104348
rect 150038 104308 150063 104348
rect 149809 104285 149895 104308
rect 149977 104285 150063 104308
rect 75449 103592 75535 103615
rect 75617 103592 75703 103615
rect 75449 103552 75474 103592
rect 75474 103552 75514 103592
rect 75514 103552 75535 103592
rect 75617 103552 75638 103592
rect 75638 103552 75678 103592
rect 75678 103552 75703 103592
rect 75449 103529 75535 103552
rect 75617 103529 75703 103552
rect 90569 103592 90655 103615
rect 90737 103592 90823 103615
rect 90569 103552 90594 103592
rect 90594 103552 90634 103592
rect 90634 103552 90655 103592
rect 90737 103552 90758 103592
rect 90758 103552 90798 103592
rect 90798 103552 90823 103592
rect 90569 103529 90655 103552
rect 90737 103529 90823 103552
rect 105689 103592 105775 103615
rect 105857 103592 105943 103615
rect 105689 103552 105714 103592
rect 105714 103552 105754 103592
rect 105754 103552 105775 103592
rect 105857 103552 105878 103592
rect 105878 103552 105918 103592
rect 105918 103552 105943 103592
rect 105689 103529 105775 103552
rect 105857 103529 105943 103552
rect 120809 103592 120895 103615
rect 120977 103592 121063 103615
rect 120809 103552 120834 103592
rect 120834 103552 120874 103592
rect 120874 103552 120895 103592
rect 120977 103552 120998 103592
rect 120998 103552 121038 103592
rect 121038 103552 121063 103592
rect 120809 103529 120895 103552
rect 120977 103529 121063 103552
rect 135929 103592 136015 103615
rect 136097 103592 136183 103615
rect 135929 103552 135954 103592
rect 135954 103552 135994 103592
rect 135994 103552 136015 103592
rect 136097 103552 136118 103592
rect 136118 103552 136158 103592
rect 136158 103552 136183 103592
rect 135929 103529 136015 103552
rect 136097 103529 136183 103552
rect 151049 103592 151135 103615
rect 151217 103592 151303 103615
rect 151049 103552 151074 103592
rect 151074 103552 151114 103592
rect 151114 103552 151135 103592
rect 151217 103552 151238 103592
rect 151238 103552 151278 103592
rect 151278 103552 151303 103592
rect 151049 103529 151135 103552
rect 151217 103529 151303 103552
rect 74209 102836 74295 102859
rect 74377 102836 74463 102859
rect 74209 102796 74234 102836
rect 74234 102796 74274 102836
rect 74274 102796 74295 102836
rect 74377 102796 74398 102836
rect 74398 102796 74438 102836
rect 74438 102796 74463 102836
rect 74209 102773 74295 102796
rect 74377 102773 74463 102796
rect 89329 102836 89415 102859
rect 89497 102836 89583 102859
rect 89329 102796 89354 102836
rect 89354 102796 89394 102836
rect 89394 102796 89415 102836
rect 89497 102796 89518 102836
rect 89518 102796 89558 102836
rect 89558 102796 89583 102836
rect 89329 102773 89415 102796
rect 89497 102773 89583 102796
rect 104449 102836 104535 102859
rect 104617 102836 104703 102859
rect 104449 102796 104474 102836
rect 104474 102796 104514 102836
rect 104514 102796 104535 102836
rect 104617 102796 104638 102836
rect 104638 102796 104678 102836
rect 104678 102796 104703 102836
rect 104449 102773 104535 102796
rect 104617 102773 104703 102796
rect 119569 102836 119655 102859
rect 119737 102836 119823 102859
rect 119569 102796 119594 102836
rect 119594 102796 119634 102836
rect 119634 102796 119655 102836
rect 119737 102796 119758 102836
rect 119758 102796 119798 102836
rect 119798 102796 119823 102836
rect 119569 102773 119655 102796
rect 119737 102773 119823 102796
rect 134689 102836 134775 102859
rect 134857 102836 134943 102859
rect 134689 102796 134714 102836
rect 134714 102796 134754 102836
rect 134754 102796 134775 102836
rect 134857 102796 134878 102836
rect 134878 102796 134918 102836
rect 134918 102796 134943 102836
rect 134689 102773 134775 102796
rect 134857 102773 134943 102796
rect 149809 102836 149895 102859
rect 149977 102836 150063 102859
rect 149809 102796 149834 102836
rect 149834 102796 149874 102836
rect 149874 102796 149895 102836
rect 149977 102796 149998 102836
rect 149998 102796 150038 102836
rect 150038 102796 150063 102836
rect 149809 102773 149895 102796
rect 149977 102773 150063 102796
rect 75449 102080 75535 102103
rect 75617 102080 75703 102103
rect 75449 102040 75474 102080
rect 75474 102040 75514 102080
rect 75514 102040 75535 102080
rect 75617 102040 75638 102080
rect 75638 102040 75678 102080
rect 75678 102040 75703 102080
rect 75449 102017 75535 102040
rect 75617 102017 75703 102040
rect 90569 102080 90655 102103
rect 90737 102080 90823 102103
rect 90569 102040 90594 102080
rect 90594 102040 90634 102080
rect 90634 102040 90655 102080
rect 90737 102040 90758 102080
rect 90758 102040 90798 102080
rect 90798 102040 90823 102080
rect 90569 102017 90655 102040
rect 90737 102017 90823 102040
rect 105689 102080 105775 102103
rect 105857 102080 105943 102103
rect 105689 102040 105714 102080
rect 105714 102040 105754 102080
rect 105754 102040 105775 102080
rect 105857 102040 105878 102080
rect 105878 102040 105918 102080
rect 105918 102040 105943 102080
rect 105689 102017 105775 102040
rect 105857 102017 105943 102040
rect 120809 102080 120895 102103
rect 120977 102080 121063 102103
rect 120809 102040 120834 102080
rect 120834 102040 120874 102080
rect 120874 102040 120895 102080
rect 120977 102040 120998 102080
rect 120998 102040 121038 102080
rect 121038 102040 121063 102080
rect 120809 102017 120895 102040
rect 120977 102017 121063 102040
rect 135929 102080 136015 102103
rect 136097 102080 136183 102103
rect 135929 102040 135954 102080
rect 135954 102040 135994 102080
rect 135994 102040 136015 102080
rect 136097 102040 136118 102080
rect 136118 102040 136158 102080
rect 136158 102040 136183 102080
rect 135929 102017 136015 102040
rect 136097 102017 136183 102040
rect 151049 102080 151135 102103
rect 151217 102080 151303 102103
rect 151049 102040 151074 102080
rect 151074 102040 151114 102080
rect 151114 102040 151135 102080
rect 151217 102040 151238 102080
rect 151238 102040 151278 102080
rect 151278 102040 151303 102080
rect 151049 102017 151135 102040
rect 151217 102017 151303 102040
rect 74209 101324 74295 101347
rect 74377 101324 74463 101347
rect 74209 101284 74234 101324
rect 74234 101284 74274 101324
rect 74274 101284 74295 101324
rect 74377 101284 74398 101324
rect 74398 101284 74438 101324
rect 74438 101284 74463 101324
rect 74209 101261 74295 101284
rect 74377 101261 74463 101284
rect 89329 101324 89415 101347
rect 89497 101324 89583 101347
rect 89329 101284 89354 101324
rect 89354 101284 89394 101324
rect 89394 101284 89415 101324
rect 89497 101284 89518 101324
rect 89518 101284 89558 101324
rect 89558 101284 89583 101324
rect 89329 101261 89415 101284
rect 89497 101261 89583 101284
rect 104449 101324 104535 101347
rect 104617 101324 104703 101347
rect 104449 101284 104474 101324
rect 104474 101284 104514 101324
rect 104514 101284 104535 101324
rect 104617 101284 104638 101324
rect 104638 101284 104678 101324
rect 104678 101284 104703 101324
rect 104449 101261 104535 101284
rect 104617 101261 104703 101284
rect 119569 101324 119655 101347
rect 119737 101324 119823 101347
rect 119569 101284 119594 101324
rect 119594 101284 119634 101324
rect 119634 101284 119655 101324
rect 119737 101284 119758 101324
rect 119758 101284 119798 101324
rect 119798 101284 119823 101324
rect 119569 101261 119655 101284
rect 119737 101261 119823 101284
rect 134689 101324 134775 101347
rect 134857 101324 134943 101347
rect 134689 101284 134714 101324
rect 134714 101284 134754 101324
rect 134754 101284 134775 101324
rect 134857 101284 134878 101324
rect 134878 101284 134918 101324
rect 134918 101284 134943 101324
rect 134689 101261 134775 101284
rect 134857 101261 134943 101284
rect 149809 101324 149895 101347
rect 149977 101324 150063 101347
rect 149809 101284 149834 101324
rect 149834 101284 149874 101324
rect 149874 101284 149895 101324
rect 149977 101284 149998 101324
rect 149998 101284 150038 101324
rect 150038 101284 150063 101324
rect 149809 101261 149895 101284
rect 149977 101261 150063 101284
rect 75449 100568 75535 100591
rect 75617 100568 75703 100591
rect 75449 100528 75474 100568
rect 75474 100528 75514 100568
rect 75514 100528 75535 100568
rect 75617 100528 75638 100568
rect 75638 100528 75678 100568
rect 75678 100528 75703 100568
rect 75449 100505 75535 100528
rect 75617 100505 75703 100528
rect 90569 100568 90655 100591
rect 90737 100568 90823 100591
rect 90569 100528 90594 100568
rect 90594 100528 90634 100568
rect 90634 100528 90655 100568
rect 90737 100528 90758 100568
rect 90758 100528 90798 100568
rect 90798 100528 90823 100568
rect 90569 100505 90655 100528
rect 90737 100505 90823 100528
rect 105689 100568 105775 100591
rect 105857 100568 105943 100591
rect 105689 100528 105714 100568
rect 105714 100528 105754 100568
rect 105754 100528 105775 100568
rect 105857 100528 105878 100568
rect 105878 100528 105918 100568
rect 105918 100528 105943 100568
rect 105689 100505 105775 100528
rect 105857 100505 105943 100528
rect 120809 100568 120895 100591
rect 120977 100568 121063 100591
rect 120809 100528 120834 100568
rect 120834 100528 120874 100568
rect 120874 100528 120895 100568
rect 120977 100528 120998 100568
rect 120998 100528 121038 100568
rect 121038 100528 121063 100568
rect 120809 100505 120895 100528
rect 120977 100505 121063 100528
rect 135929 100568 136015 100591
rect 136097 100568 136183 100591
rect 135929 100528 135954 100568
rect 135954 100528 135994 100568
rect 135994 100528 136015 100568
rect 136097 100528 136118 100568
rect 136118 100528 136158 100568
rect 136158 100528 136183 100568
rect 135929 100505 136015 100528
rect 136097 100505 136183 100528
rect 151049 100568 151135 100591
rect 151217 100568 151303 100591
rect 151049 100528 151074 100568
rect 151074 100528 151114 100568
rect 151114 100528 151135 100568
rect 151217 100528 151238 100568
rect 151238 100528 151278 100568
rect 151278 100528 151303 100568
rect 151049 100505 151135 100528
rect 151217 100505 151303 100528
rect 74209 99812 74295 99835
rect 74377 99812 74463 99835
rect 74209 99772 74234 99812
rect 74234 99772 74274 99812
rect 74274 99772 74295 99812
rect 74377 99772 74398 99812
rect 74398 99772 74438 99812
rect 74438 99772 74463 99812
rect 74209 99749 74295 99772
rect 74377 99749 74463 99772
rect 89329 99812 89415 99835
rect 89497 99812 89583 99835
rect 89329 99772 89354 99812
rect 89354 99772 89394 99812
rect 89394 99772 89415 99812
rect 89497 99772 89518 99812
rect 89518 99772 89558 99812
rect 89558 99772 89583 99812
rect 89329 99749 89415 99772
rect 89497 99749 89583 99772
rect 104449 99812 104535 99835
rect 104617 99812 104703 99835
rect 104449 99772 104474 99812
rect 104474 99772 104514 99812
rect 104514 99772 104535 99812
rect 104617 99772 104638 99812
rect 104638 99772 104678 99812
rect 104678 99772 104703 99812
rect 104449 99749 104535 99772
rect 104617 99749 104703 99772
rect 119569 99812 119655 99835
rect 119737 99812 119823 99835
rect 119569 99772 119594 99812
rect 119594 99772 119634 99812
rect 119634 99772 119655 99812
rect 119737 99772 119758 99812
rect 119758 99772 119798 99812
rect 119798 99772 119823 99812
rect 119569 99749 119655 99772
rect 119737 99749 119823 99772
rect 134689 99812 134775 99835
rect 134857 99812 134943 99835
rect 134689 99772 134714 99812
rect 134714 99772 134754 99812
rect 134754 99772 134775 99812
rect 134857 99772 134878 99812
rect 134878 99772 134918 99812
rect 134918 99772 134943 99812
rect 134689 99749 134775 99772
rect 134857 99749 134943 99772
rect 149809 99812 149895 99835
rect 149977 99812 150063 99835
rect 149809 99772 149834 99812
rect 149834 99772 149874 99812
rect 149874 99772 149895 99812
rect 149977 99772 149998 99812
rect 149998 99772 150038 99812
rect 150038 99772 150063 99812
rect 149809 99749 149895 99772
rect 149977 99749 150063 99772
rect 75449 99056 75535 99079
rect 75617 99056 75703 99079
rect 75449 99016 75474 99056
rect 75474 99016 75514 99056
rect 75514 99016 75535 99056
rect 75617 99016 75638 99056
rect 75638 99016 75678 99056
rect 75678 99016 75703 99056
rect 75449 98993 75535 99016
rect 75617 98993 75703 99016
rect 90569 99056 90655 99079
rect 90737 99056 90823 99079
rect 90569 99016 90594 99056
rect 90594 99016 90634 99056
rect 90634 99016 90655 99056
rect 90737 99016 90758 99056
rect 90758 99016 90798 99056
rect 90798 99016 90823 99056
rect 90569 98993 90655 99016
rect 90737 98993 90823 99016
rect 105689 99056 105775 99079
rect 105857 99056 105943 99079
rect 105689 99016 105714 99056
rect 105714 99016 105754 99056
rect 105754 99016 105775 99056
rect 105857 99016 105878 99056
rect 105878 99016 105918 99056
rect 105918 99016 105943 99056
rect 105689 98993 105775 99016
rect 105857 98993 105943 99016
rect 120809 99056 120895 99079
rect 120977 99056 121063 99079
rect 120809 99016 120834 99056
rect 120834 99016 120874 99056
rect 120874 99016 120895 99056
rect 120977 99016 120998 99056
rect 120998 99016 121038 99056
rect 121038 99016 121063 99056
rect 120809 98993 120895 99016
rect 120977 98993 121063 99016
rect 135929 99056 136015 99079
rect 136097 99056 136183 99079
rect 135929 99016 135954 99056
rect 135954 99016 135994 99056
rect 135994 99016 136015 99056
rect 136097 99016 136118 99056
rect 136118 99016 136158 99056
rect 136158 99016 136183 99056
rect 135929 98993 136015 99016
rect 136097 98993 136183 99016
rect 151049 99056 151135 99079
rect 151217 99056 151303 99079
rect 151049 99016 151074 99056
rect 151074 99016 151114 99056
rect 151114 99016 151135 99056
rect 151217 99016 151238 99056
rect 151238 99016 151278 99056
rect 151278 99016 151303 99056
rect 151049 98993 151135 99016
rect 151217 98993 151303 99016
rect 74209 98300 74295 98323
rect 74377 98300 74463 98323
rect 74209 98260 74234 98300
rect 74234 98260 74274 98300
rect 74274 98260 74295 98300
rect 74377 98260 74398 98300
rect 74398 98260 74438 98300
rect 74438 98260 74463 98300
rect 74209 98237 74295 98260
rect 74377 98237 74463 98260
rect 89329 98300 89415 98323
rect 89497 98300 89583 98323
rect 89329 98260 89354 98300
rect 89354 98260 89394 98300
rect 89394 98260 89415 98300
rect 89497 98260 89518 98300
rect 89518 98260 89558 98300
rect 89558 98260 89583 98300
rect 89329 98237 89415 98260
rect 89497 98237 89583 98260
rect 104449 98300 104535 98323
rect 104617 98300 104703 98323
rect 104449 98260 104474 98300
rect 104474 98260 104514 98300
rect 104514 98260 104535 98300
rect 104617 98260 104638 98300
rect 104638 98260 104678 98300
rect 104678 98260 104703 98300
rect 104449 98237 104535 98260
rect 104617 98237 104703 98260
rect 119569 98300 119655 98323
rect 119737 98300 119823 98323
rect 119569 98260 119594 98300
rect 119594 98260 119634 98300
rect 119634 98260 119655 98300
rect 119737 98260 119758 98300
rect 119758 98260 119798 98300
rect 119798 98260 119823 98300
rect 119569 98237 119655 98260
rect 119737 98237 119823 98260
rect 134689 98300 134775 98323
rect 134857 98300 134943 98323
rect 134689 98260 134714 98300
rect 134714 98260 134754 98300
rect 134754 98260 134775 98300
rect 134857 98260 134878 98300
rect 134878 98260 134918 98300
rect 134918 98260 134943 98300
rect 134689 98237 134775 98260
rect 134857 98237 134943 98260
rect 149809 98300 149895 98323
rect 149977 98300 150063 98323
rect 149809 98260 149834 98300
rect 149834 98260 149874 98300
rect 149874 98260 149895 98300
rect 149977 98260 149998 98300
rect 149998 98260 150038 98300
rect 150038 98260 150063 98300
rect 149809 98237 149895 98260
rect 149977 98237 150063 98260
rect 75449 97544 75535 97567
rect 75617 97544 75703 97567
rect 75449 97504 75474 97544
rect 75474 97504 75514 97544
rect 75514 97504 75535 97544
rect 75617 97504 75638 97544
rect 75638 97504 75678 97544
rect 75678 97504 75703 97544
rect 75449 97481 75535 97504
rect 75617 97481 75703 97504
rect 90569 97544 90655 97567
rect 90737 97544 90823 97567
rect 90569 97504 90594 97544
rect 90594 97504 90634 97544
rect 90634 97504 90655 97544
rect 90737 97504 90758 97544
rect 90758 97504 90798 97544
rect 90798 97504 90823 97544
rect 90569 97481 90655 97504
rect 90737 97481 90823 97504
rect 105689 97544 105775 97567
rect 105857 97544 105943 97567
rect 105689 97504 105714 97544
rect 105714 97504 105754 97544
rect 105754 97504 105775 97544
rect 105857 97504 105878 97544
rect 105878 97504 105918 97544
rect 105918 97504 105943 97544
rect 105689 97481 105775 97504
rect 105857 97481 105943 97504
rect 120809 97544 120895 97567
rect 120977 97544 121063 97567
rect 120809 97504 120834 97544
rect 120834 97504 120874 97544
rect 120874 97504 120895 97544
rect 120977 97504 120998 97544
rect 120998 97504 121038 97544
rect 121038 97504 121063 97544
rect 120809 97481 120895 97504
rect 120977 97481 121063 97504
rect 135929 97544 136015 97567
rect 136097 97544 136183 97567
rect 135929 97504 135954 97544
rect 135954 97504 135994 97544
rect 135994 97504 136015 97544
rect 136097 97504 136118 97544
rect 136118 97504 136158 97544
rect 136158 97504 136183 97544
rect 135929 97481 136015 97504
rect 136097 97481 136183 97504
rect 151049 97544 151135 97567
rect 151217 97544 151303 97567
rect 151049 97504 151074 97544
rect 151074 97504 151114 97544
rect 151114 97504 151135 97544
rect 151217 97504 151238 97544
rect 151238 97504 151278 97544
rect 151278 97504 151303 97544
rect 151049 97481 151135 97504
rect 151217 97481 151303 97504
rect 74209 96788 74295 96811
rect 74377 96788 74463 96811
rect 74209 96748 74234 96788
rect 74234 96748 74274 96788
rect 74274 96748 74295 96788
rect 74377 96748 74398 96788
rect 74398 96748 74438 96788
rect 74438 96748 74463 96788
rect 74209 96725 74295 96748
rect 74377 96725 74463 96748
rect 89329 96788 89415 96811
rect 89497 96788 89583 96811
rect 89329 96748 89354 96788
rect 89354 96748 89394 96788
rect 89394 96748 89415 96788
rect 89497 96748 89518 96788
rect 89518 96748 89558 96788
rect 89558 96748 89583 96788
rect 89329 96725 89415 96748
rect 89497 96725 89583 96748
rect 104449 96788 104535 96811
rect 104617 96788 104703 96811
rect 104449 96748 104474 96788
rect 104474 96748 104514 96788
rect 104514 96748 104535 96788
rect 104617 96748 104638 96788
rect 104638 96748 104678 96788
rect 104678 96748 104703 96788
rect 104449 96725 104535 96748
rect 104617 96725 104703 96748
rect 119569 96788 119655 96811
rect 119737 96788 119823 96811
rect 119569 96748 119594 96788
rect 119594 96748 119634 96788
rect 119634 96748 119655 96788
rect 119737 96748 119758 96788
rect 119758 96748 119798 96788
rect 119798 96748 119823 96788
rect 119569 96725 119655 96748
rect 119737 96725 119823 96748
rect 134689 96788 134775 96811
rect 134857 96788 134943 96811
rect 134689 96748 134714 96788
rect 134714 96748 134754 96788
rect 134754 96748 134775 96788
rect 134857 96748 134878 96788
rect 134878 96748 134918 96788
rect 134918 96748 134943 96788
rect 134689 96725 134775 96748
rect 134857 96725 134943 96748
rect 149809 96788 149895 96811
rect 149977 96788 150063 96811
rect 149809 96748 149834 96788
rect 149834 96748 149874 96788
rect 149874 96748 149895 96788
rect 149977 96748 149998 96788
rect 149998 96748 150038 96788
rect 150038 96748 150063 96788
rect 149809 96725 149895 96748
rect 149977 96725 150063 96748
rect 75449 96032 75535 96055
rect 75617 96032 75703 96055
rect 75449 95992 75474 96032
rect 75474 95992 75514 96032
rect 75514 95992 75535 96032
rect 75617 95992 75638 96032
rect 75638 95992 75678 96032
rect 75678 95992 75703 96032
rect 75449 95969 75535 95992
rect 75617 95969 75703 95992
rect 90569 96032 90655 96055
rect 90737 96032 90823 96055
rect 90569 95992 90594 96032
rect 90594 95992 90634 96032
rect 90634 95992 90655 96032
rect 90737 95992 90758 96032
rect 90758 95992 90798 96032
rect 90798 95992 90823 96032
rect 90569 95969 90655 95992
rect 90737 95969 90823 95992
rect 105689 96032 105775 96055
rect 105857 96032 105943 96055
rect 105689 95992 105714 96032
rect 105714 95992 105754 96032
rect 105754 95992 105775 96032
rect 105857 95992 105878 96032
rect 105878 95992 105918 96032
rect 105918 95992 105943 96032
rect 105689 95969 105775 95992
rect 105857 95969 105943 95992
rect 120809 96032 120895 96055
rect 120977 96032 121063 96055
rect 120809 95992 120834 96032
rect 120834 95992 120874 96032
rect 120874 95992 120895 96032
rect 120977 95992 120998 96032
rect 120998 95992 121038 96032
rect 121038 95992 121063 96032
rect 120809 95969 120895 95992
rect 120977 95969 121063 95992
rect 135929 96032 136015 96055
rect 136097 96032 136183 96055
rect 135929 95992 135954 96032
rect 135954 95992 135994 96032
rect 135994 95992 136015 96032
rect 136097 95992 136118 96032
rect 136118 95992 136158 96032
rect 136158 95992 136183 96032
rect 135929 95969 136015 95992
rect 136097 95969 136183 95992
rect 151049 96032 151135 96055
rect 151217 96032 151303 96055
rect 151049 95992 151074 96032
rect 151074 95992 151114 96032
rect 151114 95992 151135 96032
rect 151217 95992 151238 96032
rect 151238 95992 151278 96032
rect 151278 95992 151303 96032
rect 151049 95969 151135 95992
rect 151217 95969 151303 95992
rect 74209 95276 74295 95299
rect 74377 95276 74463 95299
rect 74209 95236 74234 95276
rect 74234 95236 74274 95276
rect 74274 95236 74295 95276
rect 74377 95236 74398 95276
rect 74398 95236 74438 95276
rect 74438 95236 74463 95276
rect 74209 95213 74295 95236
rect 74377 95213 74463 95236
rect 89329 95276 89415 95299
rect 89497 95276 89583 95299
rect 89329 95236 89354 95276
rect 89354 95236 89394 95276
rect 89394 95236 89415 95276
rect 89497 95236 89518 95276
rect 89518 95236 89558 95276
rect 89558 95236 89583 95276
rect 89329 95213 89415 95236
rect 89497 95213 89583 95236
rect 104449 95276 104535 95299
rect 104617 95276 104703 95299
rect 104449 95236 104474 95276
rect 104474 95236 104514 95276
rect 104514 95236 104535 95276
rect 104617 95236 104638 95276
rect 104638 95236 104678 95276
rect 104678 95236 104703 95276
rect 104449 95213 104535 95236
rect 104617 95213 104703 95236
rect 119569 95276 119655 95299
rect 119737 95276 119823 95299
rect 119569 95236 119594 95276
rect 119594 95236 119634 95276
rect 119634 95236 119655 95276
rect 119737 95236 119758 95276
rect 119758 95236 119798 95276
rect 119798 95236 119823 95276
rect 119569 95213 119655 95236
rect 119737 95213 119823 95236
rect 134689 95276 134775 95299
rect 134857 95276 134943 95299
rect 134689 95236 134714 95276
rect 134714 95236 134754 95276
rect 134754 95236 134775 95276
rect 134857 95236 134878 95276
rect 134878 95236 134918 95276
rect 134918 95236 134943 95276
rect 134689 95213 134775 95236
rect 134857 95213 134943 95236
rect 149809 95276 149895 95299
rect 149977 95276 150063 95299
rect 149809 95236 149834 95276
rect 149834 95236 149874 95276
rect 149874 95236 149895 95276
rect 149977 95236 149998 95276
rect 149998 95236 150038 95276
rect 150038 95236 150063 95276
rect 149809 95213 149895 95236
rect 149977 95213 150063 95236
rect 75449 94520 75535 94543
rect 75617 94520 75703 94543
rect 75449 94480 75474 94520
rect 75474 94480 75514 94520
rect 75514 94480 75535 94520
rect 75617 94480 75638 94520
rect 75638 94480 75678 94520
rect 75678 94480 75703 94520
rect 75449 94457 75535 94480
rect 75617 94457 75703 94480
rect 90569 94520 90655 94543
rect 90737 94520 90823 94543
rect 90569 94480 90594 94520
rect 90594 94480 90634 94520
rect 90634 94480 90655 94520
rect 90737 94480 90758 94520
rect 90758 94480 90798 94520
rect 90798 94480 90823 94520
rect 90569 94457 90655 94480
rect 90737 94457 90823 94480
rect 105689 94520 105775 94543
rect 105857 94520 105943 94543
rect 105689 94480 105714 94520
rect 105714 94480 105754 94520
rect 105754 94480 105775 94520
rect 105857 94480 105878 94520
rect 105878 94480 105918 94520
rect 105918 94480 105943 94520
rect 105689 94457 105775 94480
rect 105857 94457 105943 94480
rect 120809 94520 120895 94543
rect 120977 94520 121063 94543
rect 120809 94480 120834 94520
rect 120834 94480 120874 94520
rect 120874 94480 120895 94520
rect 120977 94480 120998 94520
rect 120998 94480 121038 94520
rect 121038 94480 121063 94520
rect 120809 94457 120895 94480
rect 120977 94457 121063 94480
rect 135929 94520 136015 94543
rect 136097 94520 136183 94543
rect 135929 94480 135954 94520
rect 135954 94480 135994 94520
rect 135994 94480 136015 94520
rect 136097 94480 136118 94520
rect 136118 94480 136158 94520
rect 136158 94480 136183 94520
rect 135929 94457 136015 94480
rect 136097 94457 136183 94480
rect 151049 94520 151135 94543
rect 151217 94520 151303 94543
rect 151049 94480 151074 94520
rect 151074 94480 151114 94520
rect 151114 94480 151135 94520
rect 151217 94480 151238 94520
rect 151238 94480 151278 94520
rect 151278 94480 151303 94520
rect 151049 94457 151135 94480
rect 151217 94457 151303 94480
rect 74209 93764 74295 93787
rect 74377 93764 74463 93787
rect 74209 93724 74234 93764
rect 74234 93724 74274 93764
rect 74274 93724 74295 93764
rect 74377 93724 74398 93764
rect 74398 93724 74438 93764
rect 74438 93724 74463 93764
rect 74209 93701 74295 93724
rect 74377 93701 74463 93724
rect 89329 93764 89415 93787
rect 89497 93764 89583 93787
rect 89329 93724 89354 93764
rect 89354 93724 89394 93764
rect 89394 93724 89415 93764
rect 89497 93724 89518 93764
rect 89518 93724 89558 93764
rect 89558 93724 89583 93764
rect 89329 93701 89415 93724
rect 89497 93701 89583 93724
rect 104449 93764 104535 93787
rect 104617 93764 104703 93787
rect 104449 93724 104474 93764
rect 104474 93724 104514 93764
rect 104514 93724 104535 93764
rect 104617 93724 104638 93764
rect 104638 93724 104678 93764
rect 104678 93724 104703 93764
rect 104449 93701 104535 93724
rect 104617 93701 104703 93724
rect 119569 93764 119655 93787
rect 119737 93764 119823 93787
rect 119569 93724 119594 93764
rect 119594 93724 119634 93764
rect 119634 93724 119655 93764
rect 119737 93724 119758 93764
rect 119758 93724 119798 93764
rect 119798 93724 119823 93764
rect 119569 93701 119655 93724
rect 119737 93701 119823 93724
rect 134689 93764 134775 93787
rect 134857 93764 134943 93787
rect 134689 93724 134714 93764
rect 134714 93724 134754 93764
rect 134754 93724 134775 93764
rect 134857 93724 134878 93764
rect 134878 93724 134918 93764
rect 134918 93724 134943 93764
rect 134689 93701 134775 93724
rect 134857 93701 134943 93724
rect 149809 93764 149895 93787
rect 149977 93764 150063 93787
rect 149809 93724 149834 93764
rect 149834 93724 149874 93764
rect 149874 93724 149895 93764
rect 149977 93724 149998 93764
rect 149998 93724 150038 93764
rect 150038 93724 150063 93764
rect 149809 93701 149895 93724
rect 149977 93701 150063 93724
rect 75449 93008 75535 93031
rect 75617 93008 75703 93031
rect 75449 92968 75474 93008
rect 75474 92968 75514 93008
rect 75514 92968 75535 93008
rect 75617 92968 75638 93008
rect 75638 92968 75678 93008
rect 75678 92968 75703 93008
rect 75449 92945 75535 92968
rect 75617 92945 75703 92968
rect 90569 93008 90655 93031
rect 90737 93008 90823 93031
rect 90569 92968 90594 93008
rect 90594 92968 90634 93008
rect 90634 92968 90655 93008
rect 90737 92968 90758 93008
rect 90758 92968 90798 93008
rect 90798 92968 90823 93008
rect 90569 92945 90655 92968
rect 90737 92945 90823 92968
rect 105689 93008 105775 93031
rect 105857 93008 105943 93031
rect 105689 92968 105714 93008
rect 105714 92968 105754 93008
rect 105754 92968 105775 93008
rect 105857 92968 105878 93008
rect 105878 92968 105918 93008
rect 105918 92968 105943 93008
rect 105689 92945 105775 92968
rect 105857 92945 105943 92968
rect 120809 93008 120895 93031
rect 120977 93008 121063 93031
rect 120809 92968 120834 93008
rect 120834 92968 120874 93008
rect 120874 92968 120895 93008
rect 120977 92968 120998 93008
rect 120998 92968 121038 93008
rect 121038 92968 121063 93008
rect 120809 92945 120895 92968
rect 120977 92945 121063 92968
rect 135929 93008 136015 93031
rect 136097 93008 136183 93031
rect 135929 92968 135954 93008
rect 135954 92968 135994 93008
rect 135994 92968 136015 93008
rect 136097 92968 136118 93008
rect 136118 92968 136158 93008
rect 136158 92968 136183 93008
rect 135929 92945 136015 92968
rect 136097 92945 136183 92968
rect 151049 93008 151135 93031
rect 151217 93008 151303 93031
rect 151049 92968 151074 93008
rect 151074 92968 151114 93008
rect 151114 92968 151135 93008
rect 151217 92968 151238 93008
rect 151238 92968 151278 93008
rect 151278 92968 151303 93008
rect 151049 92945 151135 92968
rect 151217 92945 151303 92968
rect 74209 92252 74295 92275
rect 74377 92252 74463 92275
rect 74209 92212 74234 92252
rect 74234 92212 74274 92252
rect 74274 92212 74295 92252
rect 74377 92212 74398 92252
rect 74398 92212 74438 92252
rect 74438 92212 74463 92252
rect 74209 92189 74295 92212
rect 74377 92189 74463 92212
rect 89329 92252 89415 92275
rect 89497 92252 89583 92275
rect 89329 92212 89354 92252
rect 89354 92212 89394 92252
rect 89394 92212 89415 92252
rect 89497 92212 89518 92252
rect 89518 92212 89558 92252
rect 89558 92212 89583 92252
rect 89329 92189 89415 92212
rect 89497 92189 89583 92212
rect 104449 92252 104535 92275
rect 104617 92252 104703 92275
rect 104449 92212 104474 92252
rect 104474 92212 104514 92252
rect 104514 92212 104535 92252
rect 104617 92212 104638 92252
rect 104638 92212 104678 92252
rect 104678 92212 104703 92252
rect 104449 92189 104535 92212
rect 104617 92189 104703 92212
rect 119569 92252 119655 92275
rect 119737 92252 119823 92275
rect 119569 92212 119594 92252
rect 119594 92212 119634 92252
rect 119634 92212 119655 92252
rect 119737 92212 119758 92252
rect 119758 92212 119798 92252
rect 119798 92212 119823 92252
rect 119569 92189 119655 92212
rect 119737 92189 119823 92212
rect 134689 92252 134775 92275
rect 134857 92252 134943 92275
rect 134689 92212 134714 92252
rect 134714 92212 134754 92252
rect 134754 92212 134775 92252
rect 134857 92212 134878 92252
rect 134878 92212 134918 92252
rect 134918 92212 134943 92252
rect 134689 92189 134775 92212
rect 134857 92189 134943 92212
rect 149809 92252 149895 92275
rect 149977 92252 150063 92275
rect 149809 92212 149834 92252
rect 149834 92212 149874 92252
rect 149874 92212 149895 92252
rect 149977 92212 149998 92252
rect 149998 92212 150038 92252
rect 150038 92212 150063 92252
rect 149809 92189 149895 92212
rect 149977 92189 150063 92212
rect 75449 91496 75535 91519
rect 75617 91496 75703 91519
rect 75449 91456 75474 91496
rect 75474 91456 75514 91496
rect 75514 91456 75535 91496
rect 75617 91456 75638 91496
rect 75638 91456 75678 91496
rect 75678 91456 75703 91496
rect 75449 91433 75535 91456
rect 75617 91433 75703 91456
rect 90569 91496 90655 91519
rect 90737 91496 90823 91519
rect 90569 91456 90594 91496
rect 90594 91456 90634 91496
rect 90634 91456 90655 91496
rect 90737 91456 90758 91496
rect 90758 91456 90798 91496
rect 90798 91456 90823 91496
rect 90569 91433 90655 91456
rect 90737 91433 90823 91456
rect 105689 91496 105775 91519
rect 105857 91496 105943 91519
rect 105689 91456 105714 91496
rect 105714 91456 105754 91496
rect 105754 91456 105775 91496
rect 105857 91456 105878 91496
rect 105878 91456 105918 91496
rect 105918 91456 105943 91496
rect 105689 91433 105775 91456
rect 105857 91433 105943 91456
rect 120809 91496 120895 91519
rect 120977 91496 121063 91519
rect 120809 91456 120834 91496
rect 120834 91456 120874 91496
rect 120874 91456 120895 91496
rect 120977 91456 120998 91496
rect 120998 91456 121038 91496
rect 121038 91456 121063 91496
rect 120809 91433 120895 91456
rect 120977 91433 121063 91456
rect 135929 91496 136015 91519
rect 136097 91496 136183 91519
rect 135929 91456 135954 91496
rect 135954 91456 135994 91496
rect 135994 91456 136015 91496
rect 136097 91456 136118 91496
rect 136118 91456 136158 91496
rect 136158 91456 136183 91496
rect 135929 91433 136015 91456
rect 136097 91433 136183 91456
rect 151049 91496 151135 91519
rect 151217 91496 151303 91519
rect 151049 91456 151074 91496
rect 151074 91456 151114 91496
rect 151114 91456 151135 91496
rect 151217 91456 151238 91496
rect 151238 91456 151278 91496
rect 151278 91456 151303 91496
rect 151049 91433 151135 91456
rect 151217 91433 151303 91456
rect 74209 90740 74295 90763
rect 74377 90740 74463 90763
rect 74209 90700 74234 90740
rect 74234 90700 74274 90740
rect 74274 90700 74295 90740
rect 74377 90700 74398 90740
rect 74398 90700 74438 90740
rect 74438 90700 74463 90740
rect 74209 90677 74295 90700
rect 74377 90677 74463 90700
rect 89329 90740 89415 90763
rect 89497 90740 89583 90763
rect 89329 90700 89354 90740
rect 89354 90700 89394 90740
rect 89394 90700 89415 90740
rect 89497 90700 89518 90740
rect 89518 90700 89558 90740
rect 89558 90700 89583 90740
rect 89329 90677 89415 90700
rect 89497 90677 89583 90700
rect 104449 90740 104535 90763
rect 104617 90740 104703 90763
rect 104449 90700 104474 90740
rect 104474 90700 104514 90740
rect 104514 90700 104535 90740
rect 104617 90700 104638 90740
rect 104638 90700 104678 90740
rect 104678 90700 104703 90740
rect 104449 90677 104535 90700
rect 104617 90677 104703 90700
rect 119569 90740 119655 90763
rect 119737 90740 119823 90763
rect 119569 90700 119594 90740
rect 119594 90700 119634 90740
rect 119634 90700 119655 90740
rect 119737 90700 119758 90740
rect 119758 90700 119798 90740
rect 119798 90700 119823 90740
rect 119569 90677 119655 90700
rect 119737 90677 119823 90700
rect 134689 90740 134775 90763
rect 134857 90740 134943 90763
rect 134689 90700 134714 90740
rect 134714 90700 134754 90740
rect 134754 90700 134775 90740
rect 134857 90700 134878 90740
rect 134878 90700 134918 90740
rect 134918 90700 134943 90740
rect 134689 90677 134775 90700
rect 134857 90677 134943 90700
rect 149809 90740 149895 90763
rect 149977 90740 150063 90763
rect 149809 90700 149834 90740
rect 149834 90700 149874 90740
rect 149874 90700 149895 90740
rect 149977 90700 149998 90740
rect 149998 90700 150038 90740
rect 150038 90700 150063 90740
rect 149809 90677 149895 90700
rect 149977 90677 150063 90700
rect 75449 89984 75535 90007
rect 75617 89984 75703 90007
rect 75449 89944 75474 89984
rect 75474 89944 75514 89984
rect 75514 89944 75535 89984
rect 75617 89944 75638 89984
rect 75638 89944 75678 89984
rect 75678 89944 75703 89984
rect 75449 89921 75535 89944
rect 75617 89921 75703 89944
rect 90569 89984 90655 90007
rect 90737 89984 90823 90007
rect 90569 89944 90594 89984
rect 90594 89944 90634 89984
rect 90634 89944 90655 89984
rect 90737 89944 90758 89984
rect 90758 89944 90798 89984
rect 90798 89944 90823 89984
rect 90569 89921 90655 89944
rect 90737 89921 90823 89944
rect 105689 89984 105775 90007
rect 105857 89984 105943 90007
rect 105689 89944 105714 89984
rect 105714 89944 105754 89984
rect 105754 89944 105775 89984
rect 105857 89944 105878 89984
rect 105878 89944 105918 89984
rect 105918 89944 105943 89984
rect 105689 89921 105775 89944
rect 105857 89921 105943 89944
rect 120809 89984 120895 90007
rect 120977 89984 121063 90007
rect 120809 89944 120834 89984
rect 120834 89944 120874 89984
rect 120874 89944 120895 89984
rect 120977 89944 120998 89984
rect 120998 89944 121038 89984
rect 121038 89944 121063 89984
rect 120809 89921 120895 89944
rect 120977 89921 121063 89944
rect 135929 89984 136015 90007
rect 136097 89984 136183 90007
rect 135929 89944 135954 89984
rect 135954 89944 135994 89984
rect 135994 89944 136015 89984
rect 136097 89944 136118 89984
rect 136118 89944 136158 89984
rect 136158 89944 136183 89984
rect 135929 89921 136015 89944
rect 136097 89921 136183 89944
rect 151049 89984 151135 90007
rect 151217 89984 151303 90007
rect 151049 89944 151074 89984
rect 151074 89944 151114 89984
rect 151114 89944 151135 89984
rect 151217 89944 151238 89984
rect 151238 89944 151278 89984
rect 151278 89944 151303 89984
rect 151049 89921 151135 89944
rect 151217 89921 151303 89944
rect 74209 89228 74295 89251
rect 74377 89228 74463 89251
rect 74209 89188 74234 89228
rect 74234 89188 74274 89228
rect 74274 89188 74295 89228
rect 74377 89188 74398 89228
rect 74398 89188 74438 89228
rect 74438 89188 74463 89228
rect 74209 89165 74295 89188
rect 74377 89165 74463 89188
rect 89329 89228 89415 89251
rect 89497 89228 89583 89251
rect 89329 89188 89354 89228
rect 89354 89188 89394 89228
rect 89394 89188 89415 89228
rect 89497 89188 89518 89228
rect 89518 89188 89558 89228
rect 89558 89188 89583 89228
rect 89329 89165 89415 89188
rect 89497 89165 89583 89188
rect 104449 89228 104535 89251
rect 104617 89228 104703 89251
rect 104449 89188 104474 89228
rect 104474 89188 104514 89228
rect 104514 89188 104535 89228
rect 104617 89188 104638 89228
rect 104638 89188 104678 89228
rect 104678 89188 104703 89228
rect 104449 89165 104535 89188
rect 104617 89165 104703 89188
rect 119569 89228 119655 89251
rect 119737 89228 119823 89251
rect 119569 89188 119594 89228
rect 119594 89188 119634 89228
rect 119634 89188 119655 89228
rect 119737 89188 119758 89228
rect 119758 89188 119798 89228
rect 119798 89188 119823 89228
rect 119569 89165 119655 89188
rect 119737 89165 119823 89188
rect 134689 89228 134775 89251
rect 134857 89228 134943 89251
rect 134689 89188 134714 89228
rect 134714 89188 134754 89228
rect 134754 89188 134775 89228
rect 134857 89188 134878 89228
rect 134878 89188 134918 89228
rect 134918 89188 134943 89228
rect 134689 89165 134775 89188
rect 134857 89165 134943 89188
rect 149809 89228 149895 89251
rect 149977 89228 150063 89251
rect 149809 89188 149834 89228
rect 149834 89188 149874 89228
rect 149874 89188 149895 89228
rect 149977 89188 149998 89228
rect 149998 89188 150038 89228
rect 150038 89188 150063 89228
rect 149809 89165 149895 89188
rect 149977 89165 150063 89188
rect 75449 88472 75535 88495
rect 75617 88472 75703 88495
rect 75449 88432 75474 88472
rect 75474 88432 75514 88472
rect 75514 88432 75535 88472
rect 75617 88432 75638 88472
rect 75638 88432 75678 88472
rect 75678 88432 75703 88472
rect 75449 88409 75535 88432
rect 75617 88409 75703 88432
rect 90569 88472 90655 88495
rect 90737 88472 90823 88495
rect 90569 88432 90594 88472
rect 90594 88432 90634 88472
rect 90634 88432 90655 88472
rect 90737 88432 90758 88472
rect 90758 88432 90798 88472
rect 90798 88432 90823 88472
rect 90569 88409 90655 88432
rect 90737 88409 90823 88432
rect 105689 88472 105775 88495
rect 105857 88472 105943 88495
rect 105689 88432 105714 88472
rect 105714 88432 105754 88472
rect 105754 88432 105775 88472
rect 105857 88432 105878 88472
rect 105878 88432 105918 88472
rect 105918 88432 105943 88472
rect 105689 88409 105775 88432
rect 105857 88409 105943 88432
rect 120809 88472 120895 88495
rect 120977 88472 121063 88495
rect 120809 88432 120834 88472
rect 120834 88432 120874 88472
rect 120874 88432 120895 88472
rect 120977 88432 120998 88472
rect 120998 88432 121038 88472
rect 121038 88432 121063 88472
rect 120809 88409 120895 88432
rect 120977 88409 121063 88432
rect 135929 88472 136015 88495
rect 136097 88472 136183 88495
rect 135929 88432 135954 88472
rect 135954 88432 135994 88472
rect 135994 88432 136015 88472
rect 136097 88432 136118 88472
rect 136118 88432 136158 88472
rect 136158 88432 136183 88472
rect 135929 88409 136015 88432
rect 136097 88409 136183 88432
rect 151049 88472 151135 88495
rect 151217 88472 151303 88495
rect 151049 88432 151074 88472
rect 151074 88432 151114 88472
rect 151114 88432 151135 88472
rect 151217 88432 151238 88472
rect 151238 88432 151278 88472
rect 151278 88432 151303 88472
rect 151049 88409 151135 88432
rect 151217 88409 151303 88432
rect 74209 87716 74295 87739
rect 74377 87716 74463 87739
rect 74209 87676 74234 87716
rect 74234 87676 74274 87716
rect 74274 87676 74295 87716
rect 74377 87676 74398 87716
rect 74398 87676 74438 87716
rect 74438 87676 74463 87716
rect 74209 87653 74295 87676
rect 74377 87653 74463 87676
rect 89329 87716 89415 87739
rect 89497 87716 89583 87739
rect 89329 87676 89354 87716
rect 89354 87676 89394 87716
rect 89394 87676 89415 87716
rect 89497 87676 89518 87716
rect 89518 87676 89558 87716
rect 89558 87676 89583 87716
rect 89329 87653 89415 87676
rect 89497 87653 89583 87676
rect 104449 87716 104535 87739
rect 104617 87716 104703 87739
rect 104449 87676 104474 87716
rect 104474 87676 104514 87716
rect 104514 87676 104535 87716
rect 104617 87676 104638 87716
rect 104638 87676 104678 87716
rect 104678 87676 104703 87716
rect 104449 87653 104535 87676
rect 104617 87653 104703 87676
rect 119569 87716 119655 87739
rect 119737 87716 119823 87739
rect 119569 87676 119594 87716
rect 119594 87676 119634 87716
rect 119634 87676 119655 87716
rect 119737 87676 119758 87716
rect 119758 87676 119798 87716
rect 119798 87676 119823 87716
rect 119569 87653 119655 87676
rect 119737 87653 119823 87676
rect 134689 87716 134775 87739
rect 134857 87716 134943 87739
rect 134689 87676 134714 87716
rect 134714 87676 134754 87716
rect 134754 87676 134775 87716
rect 134857 87676 134878 87716
rect 134878 87676 134918 87716
rect 134918 87676 134943 87716
rect 134689 87653 134775 87676
rect 134857 87653 134943 87676
rect 149809 87716 149895 87739
rect 149977 87716 150063 87739
rect 149809 87676 149834 87716
rect 149834 87676 149874 87716
rect 149874 87676 149895 87716
rect 149977 87676 149998 87716
rect 149998 87676 150038 87716
rect 150038 87676 150063 87716
rect 149809 87653 149895 87676
rect 149977 87653 150063 87676
rect 75449 86960 75535 86983
rect 75617 86960 75703 86983
rect 75449 86920 75474 86960
rect 75474 86920 75514 86960
rect 75514 86920 75535 86960
rect 75617 86920 75638 86960
rect 75638 86920 75678 86960
rect 75678 86920 75703 86960
rect 75449 86897 75535 86920
rect 75617 86897 75703 86920
rect 90569 86960 90655 86983
rect 90737 86960 90823 86983
rect 90569 86920 90594 86960
rect 90594 86920 90634 86960
rect 90634 86920 90655 86960
rect 90737 86920 90758 86960
rect 90758 86920 90798 86960
rect 90798 86920 90823 86960
rect 90569 86897 90655 86920
rect 90737 86897 90823 86920
rect 105689 86960 105775 86983
rect 105857 86960 105943 86983
rect 105689 86920 105714 86960
rect 105714 86920 105754 86960
rect 105754 86920 105775 86960
rect 105857 86920 105878 86960
rect 105878 86920 105918 86960
rect 105918 86920 105943 86960
rect 105689 86897 105775 86920
rect 105857 86897 105943 86920
rect 120809 86960 120895 86983
rect 120977 86960 121063 86983
rect 120809 86920 120834 86960
rect 120834 86920 120874 86960
rect 120874 86920 120895 86960
rect 120977 86920 120998 86960
rect 120998 86920 121038 86960
rect 121038 86920 121063 86960
rect 120809 86897 120895 86920
rect 120977 86897 121063 86920
rect 135929 86960 136015 86983
rect 136097 86960 136183 86983
rect 135929 86920 135954 86960
rect 135954 86920 135994 86960
rect 135994 86920 136015 86960
rect 136097 86920 136118 86960
rect 136118 86920 136158 86960
rect 136158 86920 136183 86960
rect 135929 86897 136015 86920
rect 136097 86897 136183 86920
rect 151049 86960 151135 86983
rect 151217 86960 151303 86983
rect 151049 86920 151074 86960
rect 151074 86920 151114 86960
rect 151114 86920 151135 86960
rect 151217 86920 151238 86960
rect 151238 86920 151278 86960
rect 151278 86920 151303 86960
rect 151049 86897 151135 86920
rect 151217 86897 151303 86920
rect 74209 86204 74295 86227
rect 74377 86204 74463 86227
rect 74209 86164 74234 86204
rect 74234 86164 74274 86204
rect 74274 86164 74295 86204
rect 74377 86164 74398 86204
rect 74398 86164 74438 86204
rect 74438 86164 74463 86204
rect 74209 86141 74295 86164
rect 74377 86141 74463 86164
rect 89329 86204 89415 86227
rect 89497 86204 89583 86227
rect 89329 86164 89354 86204
rect 89354 86164 89394 86204
rect 89394 86164 89415 86204
rect 89497 86164 89518 86204
rect 89518 86164 89558 86204
rect 89558 86164 89583 86204
rect 89329 86141 89415 86164
rect 89497 86141 89583 86164
rect 104449 86204 104535 86227
rect 104617 86204 104703 86227
rect 104449 86164 104474 86204
rect 104474 86164 104514 86204
rect 104514 86164 104535 86204
rect 104617 86164 104638 86204
rect 104638 86164 104678 86204
rect 104678 86164 104703 86204
rect 104449 86141 104535 86164
rect 104617 86141 104703 86164
rect 119569 86204 119655 86227
rect 119737 86204 119823 86227
rect 119569 86164 119594 86204
rect 119594 86164 119634 86204
rect 119634 86164 119655 86204
rect 119737 86164 119758 86204
rect 119758 86164 119798 86204
rect 119798 86164 119823 86204
rect 119569 86141 119655 86164
rect 119737 86141 119823 86164
rect 134689 86204 134775 86227
rect 134857 86204 134943 86227
rect 134689 86164 134714 86204
rect 134714 86164 134754 86204
rect 134754 86164 134775 86204
rect 134857 86164 134878 86204
rect 134878 86164 134918 86204
rect 134918 86164 134943 86204
rect 134689 86141 134775 86164
rect 134857 86141 134943 86164
rect 149809 86204 149895 86227
rect 149977 86204 150063 86227
rect 149809 86164 149834 86204
rect 149834 86164 149874 86204
rect 149874 86164 149895 86204
rect 149977 86164 149998 86204
rect 149998 86164 150038 86204
rect 150038 86164 150063 86204
rect 149809 86141 149895 86164
rect 149977 86141 150063 86164
rect 75449 85448 75535 85471
rect 75617 85448 75703 85471
rect 75449 85408 75474 85448
rect 75474 85408 75514 85448
rect 75514 85408 75535 85448
rect 75617 85408 75638 85448
rect 75638 85408 75678 85448
rect 75678 85408 75703 85448
rect 75449 85385 75535 85408
rect 75617 85385 75703 85408
rect 90569 85448 90655 85471
rect 90737 85448 90823 85471
rect 90569 85408 90594 85448
rect 90594 85408 90634 85448
rect 90634 85408 90655 85448
rect 90737 85408 90758 85448
rect 90758 85408 90798 85448
rect 90798 85408 90823 85448
rect 90569 85385 90655 85408
rect 90737 85385 90823 85408
rect 105689 85448 105775 85471
rect 105857 85448 105943 85471
rect 105689 85408 105714 85448
rect 105714 85408 105754 85448
rect 105754 85408 105775 85448
rect 105857 85408 105878 85448
rect 105878 85408 105918 85448
rect 105918 85408 105943 85448
rect 105689 85385 105775 85408
rect 105857 85385 105943 85408
rect 120809 85448 120895 85471
rect 120977 85448 121063 85471
rect 120809 85408 120834 85448
rect 120834 85408 120874 85448
rect 120874 85408 120895 85448
rect 120977 85408 120998 85448
rect 120998 85408 121038 85448
rect 121038 85408 121063 85448
rect 120809 85385 120895 85408
rect 120977 85385 121063 85408
rect 135929 85448 136015 85471
rect 136097 85448 136183 85471
rect 135929 85408 135954 85448
rect 135954 85408 135994 85448
rect 135994 85408 136015 85448
rect 136097 85408 136118 85448
rect 136118 85408 136158 85448
rect 136158 85408 136183 85448
rect 135929 85385 136015 85408
rect 136097 85385 136183 85408
rect 151049 85448 151135 85471
rect 151217 85448 151303 85471
rect 151049 85408 151074 85448
rect 151074 85408 151114 85448
rect 151114 85408 151135 85448
rect 151217 85408 151238 85448
rect 151238 85408 151278 85448
rect 151278 85408 151303 85448
rect 151049 85385 151135 85408
rect 151217 85385 151303 85408
rect 74209 84692 74295 84715
rect 74377 84692 74463 84715
rect 74209 84652 74234 84692
rect 74234 84652 74274 84692
rect 74274 84652 74295 84692
rect 74377 84652 74398 84692
rect 74398 84652 74438 84692
rect 74438 84652 74463 84692
rect 74209 84629 74295 84652
rect 74377 84629 74463 84652
rect 89329 84692 89415 84715
rect 89497 84692 89583 84715
rect 89329 84652 89354 84692
rect 89354 84652 89394 84692
rect 89394 84652 89415 84692
rect 89497 84652 89518 84692
rect 89518 84652 89558 84692
rect 89558 84652 89583 84692
rect 89329 84629 89415 84652
rect 89497 84629 89583 84652
rect 104449 84692 104535 84715
rect 104617 84692 104703 84715
rect 104449 84652 104474 84692
rect 104474 84652 104514 84692
rect 104514 84652 104535 84692
rect 104617 84652 104638 84692
rect 104638 84652 104678 84692
rect 104678 84652 104703 84692
rect 104449 84629 104535 84652
rect 104617 84629 104703 84652
rect 119569 84692 119655 84715
rect 119737 84692 119823 84715
rect 119569 84652 119594 84692
rect 119594 84652 119634 84692
rect 119634 84652 119655 84692
rect 119737 84652 119758 84692
rect 119758 84652 119798 84692
rect 119798 84652 119823 84692
rect 119569 84629 119655 84652
rect 119737 84629 119823 84652
rect 134689 84692 134775 84715
rect 134857 84692 134943 84715
rect 134689 84652 134714 84692
rect 134714 84652 134754 84692
rect 134754 84652 134775 84692
rect 134857 84652 134878 84692
rect 134878 84652 134918 84692
rect 134918 84652 134943 84692
rect 134689 84629 134775 84652
rect 134857 84629 134943 84652
rect 149809 84692 149895 84715
rect 149977 84692 150063 84715
rect 149809 84652 149834 84692
rect 149834 84652 149874 84692
rect 149874 84652 149895 84692
rect 149977 84652 149998 84692
rect 149998 84652 150038 84692
rect 150038 84652 150063 84692
rect 149809 84629 149895 84652
rect 149977 84629 150063 84652
rect 75449 83936 75535 83959
rect 75617 83936 75703 83959
rect 75449 83896 75474 83936
rect 75474 83896 75514 83936
rect 75514 83896 75535 83936
rect 75617 83896 75638 83936
rect 75638 83896 75678 83936
rect 75678 83896 75703 83936
rect 75449 83873 75535 83896
rect 75617 83873 75703 83896
rect 90569 83936 90655 83959
rect 90737 83936 90823 83959
rect 90569 83896 90594 83936
rect 90594 83896 90634 83936
rect 90634 83896 90655 83936
rect 90737 83896 90758 83936
rect 90758 83896 90798 83936
rect 90798 83896 90823 83936
rect 90569 83873 90655 83896
rect 90737 83873 90823 83896
rect 105689 83936 105775 83959
rect 105857 83936 105943 83959
rect 105689 83896 105714 83936
rect 105714 83896 105754 83936
rect 105754 83896 105775 83936
rect 105857 83896 105878 83936
rect 105878 83896 105918 83936
rect 105918 83896 105943 83936
rect 105689 83873 105775 83896
rect 105857 83873 105943 83896
rect 120809 83936 120895 83959
rect 120977 83936 121063 83959
rect 120809 83896 120834 83936
rect 120834 83896 120874 83936
rect 120874 83896 120895 83936
rect 120977 83896 120998 83936
rect 120998 83896 121038 83936
rect 121038 83896 121063 83936
rect 120809 83873 120895 83896
rect 120977 83873 121063 83896
rect 135929 83936 136015 83959
rect 136097 83936 136183 83959
rect 135929 83896 135954 83936
rect 135954 83896 135994 83936
rect 135994 83896 136015 83936
rect 136097 83896 136118 83936
rect 136118 83896 136158 83936
rect 136158 83896 136183 83936
rect 135929 83873 136015 83896
rect 136097 83873 136183 83896
rect 151049 83936 151135 83959
rect 151217 83936 151303 83959
rect 151049 83896 151074 83936
rect 151074 83896 151114 83936
rect 151114 83896 151135 83936
rect 151217 83896 151238 83936
rect 151238 83896 151278 83936
rect 151278 83896 151303 83936
rect 151049 83873 151135 83896
rect 151217 83873 151303 83896
rect 74209 83180 74295 83203
rect 74377 83180 74463 83203
rect 74209 83140 74234 83180
rect 74234 83140 74274 83180
rect 74274 83140 74295 83180
rect 74377 83140 74398 83180
rect 74398 83140 74438 83180
rect 74438 83140 74463 83180
rect 74209 83117 74295 83140
rect 74377 83117 74463 83140
rect 89329 83180 89415 83203
rect 89497 83180 89583 83203
rect 89329 83140 89354 83180
rect 89354 83140 89394 83180
rect 89394 83140 89415 83180
rect 89497 83140 89518 83180
rect 89518 83140 89558 83180
rect 89558 83140 89583 83180
rect 89329 83117 89415 83140
rect 89497 83117 89583 83140
rect 104449 83180 104535 83203
rect 104617 83180 104703 83203
rect 104449 83140 104474 83180
rect 104474 83140 104514 83180
rect 104514 83140 104535 83180
rect 104617 83140 104638 83180
rect 104638 83140 104678 83180
rect 104678 83140 104703 83180
rect 104449 83117 104535 83140
rect 104617 83117 104703 83140
rect 119569 83180 119655 83203
rect 119737 83180 119823 83203
rect 119569 83140 119594 83180
rect 119594 83140 119634 83180
rect 119634 83140 119655 83180
rect 119737 83140 119758 83180
rect 119758 83140 119798 83180
rect 119798 83140 119823 83180
rect 119569 83117 119655 83140
rect 119737 83117 119823 83140
rect 134689 83180 134775 83203
rect 134857 83180 134943 83203
rect 134689 83140 134714 83180
rect 134714 83140 134754 83180
rect 134754 83140 134775 83180
rect 134857 83140 134878 83180
rect 134878 83140 134918 83180
rect 134918 83140 134943 83180
rect 134689 83117 134775 83140
rect 134857 83117 134943 83140
rect 149809 83180 149895 83203
rect 149977 83180 150063 83203
rect 149809 83140 149834 83180
rect 149834 83140 149874 83180
rect 149874 83140 149895 83180
rect 149977 83140 149998 83180
rect 149998 83140 150038 83180
rect 150038 83140 150063 83180
rect 149809 83117 149895 83140
rect 149977 83117 150063 83140
rect 75449 82424 75535 82447
rect 75617 82424 75703 82447
rect 75449 82384 75474 82424
rect 75474 82384 75514 82424
rect 75514 82384 75535 82424
rect 75617 82384 75638 82424
rect 75638 82384 75678 82424
rect 75678 82384 75703 82424
rect 75449 82361 75535 82384
rect 75617 82361 75703 82384
rect 90569 82424 90655 82447
rect 90737 82424 90823 82447
rect 90569 82384 90594 82424
rect 90594 82384 90634 82424
rect 90634 82384 90655 82424
rect 90737 82384 90758 82424
rect 90758 82384 90798 82424
rect 90798 82384 90823 82424
rect 90569 82361 90655 82384
rect 90737 82361 90823 82384
rect 105689 82424 105775 82447
rect 105857 82424 105943 82447
rect 105689 82384 105714 82424
rect 105714 82384 105754 82424
rect 105754 82384 105775 82424
rect 105857 82384 105878 82424
rect 105878 82384 105918 82424
rect 105918 82384 105943 82424
rect 105689 82361 105775 82384
rect 105857 82361 105943 82384
rect 120809 82424 120895 82447
rect 120977 82424 121063 82447
rect 120809 82384 120834 82424
rect 120834 82384 120874 82424
rect 120874 82384 120895 82424
rect 120977 82384 120998 82424
rect 120998 82384 121038 82424
rect 121038 82384 121063 82424
rect 120809 82361 120895 82384
rect 120977 82361 121063 82384
rect 135929 82424 136015 82447
rect 136097 82424 136183 82447
rect 135929 82384 135954 82424
rect 135954 82384 135994 82424
rect 135994 82384 136015 82424
rect 136097 82384 136118 82424
rect 136118 82384 136158 82424
rect 136158 82384 136183 82424
rect 135929 82361 136015 82384
rect 136097 82361 136183 82384
rect 151049 82424 151135 82447
rect 151217 82424 151303 82447
rect 151049 82384 151074 82424
rect 151074 82384 151114 82424
rect 151114 82384 151135 82424
rect 151217 82384 151238 82424
rect 151238 82384 151278 82424
rect 151278 82384 151303 82424
rect 151049 82361 151135 82384
rect 151217 82361 151303 82384
rect 74209 81668 74295 81691
rect 74377 81668 74463 81691
rect 74209 81628 74234 81668
rect 74234 81628 74274 81668
rect 74274 81628 74295 81668
rect 74377 81628 74398 81668
rect 74398 81628 74438 81668
rect 74438 81628 74463 81668
rect 74209 81605 74295 81628
rect 74377 81605 74463 81628
rect 89329 81668 89415 81691
rect 89497 81668 89583 81691
rect 89329 81628 89354 81668
rect 89354 81628 89394 81668
rect 89394 81628 89415 81668
rect 89497 81628 89518 81668
rect 89518 81628 89558 81668
rect 89558 81628 89583 81668
rect 89329 81605 89415 81628
rect 89497 81605 89583 81628
rect 104449 81668 104535 81691
rect 104617 81668 104703 81691
rect 104449 81628 104474 81668
rect 104474 81628 104514 81668
rect 104514 81628 104535 81668
rect 104617 81628 104638 81668
rect 104638 81628 104678 81668
rect 104678 81628 104703 81668
rect 104449 81605 104535 81628
rect 104617 81605 104703 81628
rect 119569 81668 119655 81691
rect 119737 81668 119823 81691
rect 119569 81628 119594 81668
rect 119594 81628 119634 81668
rect 119634 81628 119655 81668
rect 119737 81628 119758 81668
rect 119758 81628 119798 81668
rect 119798 81628 119823 81668
rect 119569 81605 119655 81628
rect 119737 81605 119823 81628
rect 134689 81668 134775 81691
rect 134857 81668 134943 81691
rect 134689 81628 134714 81668
rect 134714 81628 134754 81668
rect 134754 81628 134775 81668
rect 134857 81628 134878 81668
rect 134878 81628 134918 81668
rect 134918 81628 134943 81668
rect 134689 81605 134775 81628
rect 134857 81605 134943 81628
rect 149809 81668 149895 81691
rect 149977 81668 150063 81691
rect 149809 81628 149834 81668
rect 149834 81628 149874 81668
rect 149874 81628 149895 81668
rect 149977 81628 149998 81668
rect 149998 81628 150038 81668
rect 150038 81628 150063 81668
rect 149809 81605 149895 81628
rect 149977 81605 150063 81628
rect 75449 80912 75535 80935
rect 75617 80912 75703 80935
rect 75449 80872 75474 80912
rect 75474 80872 75514 80912
rect 75514 80872 75535 80912
rect 75617 80872 75638 80912
rect 75638 80872 75678 80912
rect 75678 80872 75703 80912
rect 75449 80849 75535 80872
rect 75617 80849 75703 80872
rect 90569 80912 90655 80935
rect 90737 80912 90823 80935
rect 90569 80872 90594 80912
rect 90594 80872 90634 80912
rect 90634 80872 90655 80912
rect 90737 80872 90758 80912
rect 90758 80872 90798 80912
rect 90798 80872 90823 80912
rect 90569 80849 90655 80872
rect 90737 80849 90823 80872
rect 105689 80912 105775 80935
rect 105857 80912 105943 80935
rect 105689 80872 105714 80912
rect 105714 80872 105754 80912
rect 105754 80872 105775 80912
rect 105857 80872 105878 80912
rect 105878 80872 105918 80912
rect 105918 80872 105943 80912
rect 105689 80849 105775 80872
rect 105857 80849 105943 80872
rect 120809 80912 120895 80935
rect 120977 80912 121063 80935
rect 120809 80872 120834 80912
rect 120834 80872 120874 80912
rect 120874 80872 120895 80912
rect 120977 80872 120998 80912
rect 120998 80872 121038 80912
rect 121038 80872 121063 80912
rect 120809 80849 120895 80872
rect 120977 80849 121063 80872
rect 135929 80912 136015 80935
rect 136097 80912 136183 80935
rect 135929 80872 135954 80912
rect 135954 80872 135994 80912
rect 135994 80872 136015 80912
rect 136097 80872 136118 80912
rect 136118 80872 136158 80912
rect 136158 80872 136183 80912
rect 135929 80849 136015 80872
rect 136097 80849 136183 80872
rect 151049 80912 151135 80935
rect 151217 80912 151303 80935
rect 151049 80872 151074 80912
rect 151074 80872 151114 80912
rect 151114 80872 151135 80912
rect 151217 80872 151238 80912
rect 151238 80872 151278 80912
rect 151278 80872 151303 80912
rect 151049 80849 151135 80872
rect 151217 80849 151303 80872
rect 74209 80156 74295 80179
rect 74377 80156 74463 80179
rect 74209 80116 74234 80156
rect 74234 80116 74274 80156
rect 74274 80116 74295 80156
rect 74377 80116 74398 80156
rect 74398 80116 74438 80156
rect 74438 80116 74463 80156
rect 74209 80093 74295 80116
rect 74377 80093 74463 80116
rect 89329 80156 89415 80179
rect 89497 80156 89583 80179
rect 89329 80116 89354 80156
rect 89354 80116 89394 80156
rect 89394 80116 89415 80156
rect 89497 80116 89518 80156
rect 89518 80116 89558 80156
rect 89558 80116 89583 80156
rect 89329 80093 89415 80116
rect 89497 80093 89583 80116
rect 104449 80156 104535 80179
rect 104617 80156 104703 80179
rect 104449 80116 104474 80156
rect 104474 80116 104514 80156
rect 104514 80116 104535 80156
rect 104617 80116 104638 80156
rect 104638 80116 104678 80156
rect 104678 80116 104703 80156
rect 104449 80093 104535 80116
rect 104617 80093 104703 80116
rect 119569 80156 119655 80179
rect 119737 80156 119823 80179
rect 119569 80116 119594 80156
rect 119594 80116 119634 80156
rect 119634 80116 119655 80156
rect 119737 80116 119758 80156
rect 119758 80116 119798 80156
rect 119798 80116 119823 80156
rect 119569 80093 119655 80116
rect 119737 80093 119823 80116
rect 134689 80156 134775 80179
rect 134857 80156 134943 80179
rect 134689 80116 134714 80156
rect 134714 80116 134754 80156
rect 134754 80116 134775 80156
rect 134857 80116 134878 80156
rect 134878 80116 134918 80156
rect 134918 80116 134943 80156
rect 134689 80093 134775 80116
rect 134857 80093 134943 80116
rect 149809 80156 149895 80179
rect 149977 80156 150063 80179
rect 149809 80116 149834 80156
rect 149834 80116 149874 80156
rect 149874 80116 149895 80156
rect 149977 80116 149998 80156
rect 149998 80116 150038 80156
rect 150038 80116 150063 80156
rect 149809 80093 149895 80116
rect 149977 80093 150063 80116
rect 75449 79400 75535 79423
rect 75617 79400 75703 79423
rect 75449 79360 75474 79400
rect 75474 79360 75514 79400
rect 75514 79360 75535 79400
rect 75617 79360 75638 79400
rect 75638 79360 75678 79400
rect 75678 79360 75703 79400
rect 75449 79337 75535 79360
rect 75617 79337 75703 79360
rect 90569 79400 90655 79423
rect 90737 79400 90823 79423
rect 90569 79360 90594 79400
rect 90594 79360 90634 79400
rect 90634 79360 90655 79400
rect 90737 79360 90758 79400
rect 90758 79360 90798 79400
rect 90798 79360 90823 79400
rect 90569 79337 90655 79360
rect 90737 79337 90823 79360
rect 105689 79400 105775 79423
rect 105857 79400 105943 79423
rect 105689 79360 105714 79400
rect 105714 79360 105754 79400
rect 105754 79360 105775 79400
rect 105857 79360 105878 79400
rect 105878 79360 105918 79400
rect 105918 79360 105943 79400
rect 105689 79337 105775 79360
rect 105857 79337 105943 79360
rect 120809 79400 120895 79423
rect 120977 79400 121063 79423
rect 120809 79360 120834 79400
rect 120834 79360 120874 79400
rect 120874 79360 120895 79400
rect 120977 79360 120998 79400
rect 120998 79360 121038 79400
rect 121038 79360 121063 79400
rect 120809 79337 120895 79360
rect 120977 79337 121063 79360
rect 135929 79400 136015 79423
rect 136097 79400 136183 79423
rect 135929 79360 135954 79400
rect 135954 79360 135994 79400
rect 135994 79360 136015 79400
rect 136097 79360 136118 79400
rect 136118 79360 136158 79400
rect 136158 79360 136183 79400
rect 135929 79337 136015 79360
rect 136097 79337 136183 79360
rect 151049 79400 151135 79423
rect 151217 79400 151303 79423
rect 151049 79360 151074 79400
rect 151074 79360 151114 79400
rect 151114 79360 151135 79400
rect 151217 79360 151238 79400
rect 151238 79360 151278 79400
rect 151278 79360 151303 79400
rect 151049 79337 151135 79360
rect 151217 79337 151303 79360
rect 74209 78644 74295 78667
rect 74377 78644 74463 78667
rect 74209 78604 74234 78644
rect 74234 78604 74274 78644
rect 74274 78604 74295 78644
rect 74377 78604 74398 78644
rect 74398 78604 74438 78644
rect 74438 78604 74463 78644
rect 74209 78581 74295 78604
rect 74377 78581 74463 78604
rect 89329 78644 89415 78667
rect 89497 78644 89583 78667
rect 89329 78604 89354 78644
rect 89354 78604 89394 78644
rect 89394 78604 89415 78644
rect 89497 78604 89518 78644
rect 89518 78604 89558 78644
rect 89558 78604 89583 78644
rect 89329 78581 89415 78604
rect 89497 78581 89583 78604
rect 104449 78644 104535 78667
rect 104617 78644 104703 78667
rect 104449 78604 104474 78644
rect 104474 78604 104514 78644
rect 104514 78604 104535 78644
rect 104617 78604 104638 78644
rect 104638 78604 104678 78644
rect 104678 78604 104703 78644
rect 104449 78581 104535 78604
rect 104617 78581 104703 78604
rect 119569 78644 119655 78667
rect 119737 78644 119823 78667
rect 119569 78604 119594 78644
rect 119594 78604 119634 78644
rect 119634 78604 119655 78644
rect 119737 78604 119758 78644
rect 119758 78604 119798 78644
rect 119798 78604 119823 78644
rect 119569 78581 119655 78604
rect 119737 78581 119823 78604
rect 134689 78644 134775 78667
rect 134857 78644 134943 78667
rect 134689 78604 134714 78644
rect 134714 78604 134754 78644
rect 134754 78604 134775 78644
rect 134857 78604 134878 78644
rect 134878 78604 134918 78644
rect 134918 78604 134943 78644
rect 134689 78581 134775 78604
rect 134857 78581 134943 78604
rect 149809 78644 149895 78667
rect 149977 78644 150063 78667
rect 149809 78604 149834 78644
rect 149834 78604 149874 78644
rect 149874 78604 149895 78644
rect 149977 78604 149998 78644
rect 149998 78604 150038 78644
rect 150038 78604 150063 78644
rect 149809 78581 149895 78604
rect 149977 78581 150063 78604
rect 75449 77888 75535 77911
rect 75617 77888 75703 77911
rect 75449 77848 75474 77888
rect 75474 77848 75514 77888
rect 75514 77848 75535 77888
rect 75617 77848 75638 77888
rect 75638 77848 75678 77888
rect 75678 77848 75703 77888
rect 75449 77825 75535 77848
rect 75617 77825 75703 77848
rect 90569 77888 90655 77911
rect 90737 77888 90823 77911
rect 90569 77848 90594 77888
rect 90594 77848 90634 77888
rect 90634 77848 90655 77888
rect 90737 77848 90758 77888
rect 90758 77848 90798 77888
rect 90798 77848 90823 77888
rect 90569 77825 90655 77848
rect 90737 77825 90823 77848
rect 105689 77888 105775 77911
rect 105857 77888 105943 77911
rect 105689 77848 105714 77888
rect 105714 77848 105754 77888
rect 105754 77848 105775 77888
rect 105857 77848 105878 77888
rect 105878 77848 105918 77888
rect 105918 77848 105943 77888
rect 105689 77825 105775 77848
rect 105857 77825 105943 77848
rect 120809 77888 120895 77911
rect 120977 77888 121063 77911
rect 120809 77848 120834 77888
rect 120834 77848 120874 77888
rect 120874 77848 120895 77888
rect 120977 77848 120998 77888
rect 120998 77848 121038 77888
rect 121038 77848 121063 77888
rect 120809 77825 120895 77848
rect 120977 77825 121063 77848
rect 135929 77888 136015 77911
rect 136097 77888 136183 77911
rect 135929 77848 135954 77888
rect 135954 77848 135994 77888
rect 135994 77848 136015 77888
rect 136097 77848 136118 77888
rect 136118 77848 136158 77888
rect 136158 77848 136183 77888
rect 135929 77825 136015 77848
rect 136097 77825 136183 77848
rect 151049 77888 151135 77911
rect 151217 77888 151303 77911
rect 151049 77848 151074 77888
rect 151074 77848 151114 77888
rect 151114 77848 151135 77888
rect 151217 77848 151238 77888
rect 151238 77848 151278 77888
rect 151278 77848 151303 77888
rect 151049 77825 151135 77848
rect 151217 77825 151303 77848
rect 74209 77132 74295 77155
rect 74377 77132 74463 77155
rect 74209 77092 74234 77132
rect 74234 77092 74274 77132
rect 74274 77092 74295 77132
rect 74377 77092 74398 77132
rect 74398 77092 74438 77132
rect 74438 77092 74463 77132
rect 74209 77069 74295 77092
rect 74377 77069 74463 77092
rect 89329 77132 89415 77155
rect 89497 77132 89583 77155
rect 89329 77092 89354 77132
rect 89354 77092 89394 77132
rect 89394 77092 89415 77132
rect 89497 77092 89518 77132
rect 89518 77092 89558 77132
rect 89558 77092 89583 77132
rect 89329 77069 89415 77092
rect 89497 77069 89583 77092
rect 104449 77132 104535 77155
rect 104617 77132 104703 77155
rect 104449 77092 104474 77132
rect 104474 77092 104514 77132
rect 104514 77092 104535 77132
rect 104617 77092 104638 77132
rect 104638 77092 104678 77132
rect 104678 77092 104703 77132
rect 104449 77069 104535 77092
rect 104617 77069 104703 77092
rect 119569 77132 119655 77155
rect 119737 77132 119823 77155
rect 119569 77092 119594 77132
rect 119594 77092 119634 77132
rect 119634 77092 119655 77132
rect 119737 77092 119758 77132
rect 119758 77092 119798 77132
rect 119798 77092 119823 77132
rect 119569 77069 119655 77092
rect 119737 77069 119823 77092
rect 134689 77132 134775 77155
rect 134857 77132 134943 77155
rect 134689 77092 134714 77132
rect 134714 77092 134754 77132
rect 134754 77092 134775 77132
rect 134857 77092 134878 77132
rect 134878 77092 134918 77132
rect 134918 77092 134943 77132
rect 134689 77069 134775 77092
rect 134857 77069 134943 77092
rect 149809 77132 149895 77155
rect 149977 77132 150063 77155
rect 149809 77092 149834 77132
rect 149834 77092 149874 77132
rect 149874 77092 149895 77132
rect 149977 77092 149998 77132
rect 149998 77092 150038 77132
rect 150038 77092 150063 77132
rect 149809 77069 149895 77092
rect 149977 77069 150063 77092
rect 75449 76376 75535 76399
rect 75617 76376 75703 76399
rect 75449 76336 75474 76376
rect 75474 76336 75514 76376
rect 75514 76336 75535 76376
rect 75617 76336 75638 76376
rect 75638 76336 75678 76376
rect 75678 76336 75703 76376
rect 75449 76313 75535 76336
rect 75617 76313 75703 76336
rect 90569 76376 90655 76399
rect 90737 76376 90823 76399
rect 90569 76336 90594 76376
rect 90594 76336 90634 76376
rect 90634 76336 90655 76376
rect 90737 76336 90758 76376
rect 90758 76336 90798 76376
rect 90798 76336 90823 76376
rect 90569 76313 90655 76336
rect 90737 76313 90823 76336
rect 105689 76376 105775 76399
rect 105857 76376 105943 76399
rect 105689 76336 105714 76376
rect 105714 76336 105754 76376
rect 105754 76336 105775 76376
rect 105857 76336 105878 76376
rect 105878 76336 105918 76376
rect 105918 76336 105943 76376
rect 105689 76313 105775 76336
rect 105857 76313 105943 76336
rect 120809 76376 120895 76399
rect 120977 76376 121063 76399
rect 120809 76336 120834 76376
rect 120834 76336 120874 76376
rect 120874 76336 120895 76376
rect 120977 76336 120998 76376
rect 120998 76336 121038 76376
rect 121038 76336 121063 76376
rect 120809 76313 120895 76336
rect 120977 76313 121063 76336
rect 135929 76376 136015 76399
rect 136097 76376 136183 76399
rect 135929 76336 135954 76376
rect 135954 76336 135994 76376
rect 135994 76336 136015 76376
rect 136097 76336 136118 76376
rect 136118 76336 136158 76376
rect 136158 76336 136183 76376
rect 135929 76313 136015 76336
rect 136097 76313 136183 76336
rect 151049 76376 151135 76399
rect 151217 76376 151303 76399
rect 151049 76336 151074 76376
rect 151074 76336 151114 76376
rect 151114 76336 151135 76376
rect 151217 76336 151238 76376
rect 151238 76336 151278 76376
rect 151278 76336 151303 76376
rect 151049 76313 151135 76336
rect 151217 76313 151303 76336
rect 74209 75620 74295 75643
rect 74377 75620 74463 75643
rect 74209 75580 74234 75620
rect 74234 75580 74274 75620
rect 74274 75580 74295 75620
rect 74377 75580 74398 75620
rect 74398 75580 74438 75620
rect 74438 75580 74463 75620
rect 74209 75557 74295 75580
rect 74377 75557 74463 75580
rect 89329 75620 89415 75643
rect 89497 75620 89583 75643
rect 89329 75580 89354 75620
rect 89354 75580 89394 75620
rect 89394 75580 89415 75620
rect 89497 75580 89518 75620
rect 89518 75580 89558 75620
rect 89558 75580 89583 75620
rect 89329 75557 89415 75580
rect 89497 75557 89583 75580
rect 104449 75620 104535 75643
rect 104617 75620 104703 75643
rect 104449 75580 104474 75620
rect 104474 75580 104514 75620
rect 104514 75580 104535 75620
rect 104617 75580 104638 75620
rect 104638 75580 104678 75620
rect 104678 75580 104703 75620
rect 104449 75557 104535 75580
rect 104617 75557 104703 75580
rect 119569 75620 119655 75643
rect 119737 75620 119823 75643
rect 119569 75580 119594 75620
rect 119594 75580 119634 75620
rect 119634 75580 119655 75620
rect 119737 75580 119758 75620
rect 119758 75580 119798 75620
rect 119798 75580 119823 75620
rect 119569 75557 119655 75580
rect 119737 75557 119823 75580
rect 134689 75620 134775 75643
rect 134857 75620 134943 75643
rect 134689 75580 134714 75620
rect 134714 75580 134754 75620
rect 134754 75580 134775 75620
rect 134857 75580 134878 75620
rect 134878 75580 134918 75620
rect 134918 75580 134943 75620
rect 134689 75557 134775 75580
rect 134857 75557 134943 75580
rect 149809 75620 149895 75643
rect 149977 75620 150063 75643
rect 149809 75580 149834 75620
rect 149834 75580 149874 75620
rect 149874 75580 149895 75620
rect 149977 75580 149998 75620
rect 149998 75580 150038 75620
rect 150038 75580 150063 75620
rect 149809 75557 149895 75580
rect 149977 75557 150063 75580
rect 75449 74864 75535 74887
rect 75617 74864 75703 74887
rect 75449 74824 75474 74864
rect 75474 74824 75514 74864
rect 75514 74824 75535 74864
rect 75617 74824 75638 74864
rect 75638 74824 75678 74864
rect 75678 74824 75703 74864
rect 75449 74801 75535 74824
rect 75617 74801 75703 74824
rect 90569 74864 90655 74887
rect 90737 74864 90823 74887
rect 90569 74824 90594 74864
rect 90594 74824 90634 74864
rect 90634 74824 90655 74864
rect 90737 74824 90758 74864
rect 90758 74824 90798 74864
rect 90798 74824 90823 74864
rect 90569 74801 90655 74824
rect 90737 74801 90823 74824
rect 105689 74864 105775 74887
rect 105857 74864 105943 74887
rect 105689 74824 105714 74864
rect 105714 74824 105754 74864
rect 105754 74824 105775 74864
rect 105857 74824 105878 74864
rect 105878 74824 105918 74864
rect 105918 74824 105943 74864
rect 105689 74801 105775 74824
rect 105857 74801 105943 74824
rect 120809 74864 120895 74887
rect 120977 74864 121063 74887
rect 120809 74824 120834 74864
rect 120834 74824 120874 74864
rect 120874 74824 120895 74864
rect 120977 74824 120998 74864
rect 120998 74824 121038 74864
rect 121038 74824 121063 74864
rect 120809 74801 120895 74824
rect 120977 74801 121063 74824
rect 135929 74864 136015 74887
rect 136097 74864 136183 74887
rect 135929 74824 135954 74864
rect 135954 74824 135994 74864
rect 135994 74824 136015 74864
rect 136097 74824 136118 74864
rect 136118 74824 136158 74864
rect 136158 74824 136183 74864
rect 135929 74801 136015 74824
rect 136097 74801 136183 74824
rect 151049 74864 151135 74887
rect 151217 74864 151303 74887
rect 151049 74824 151074 74864
rect 151074 74824 151114 74864
rect 151114 74824 151135 74864
rect 151217 74824 151238 74864
rect 151238 74824 151278 74864
rect 151278 74824 151303 74864
rect 151049 74801 151135 74824
rect 151217 74801 151303 74824
rect 74209 74108 74295 74131
rect 74377 74108 74463 74131
rect 74209 74068 74234 74108
rect 74234 74068 74274 74108
rect 74274 74068 74295 74108
rect 74377 74068 74398 74108
rect 74398 74068 74438 74108
rect 74438 74068 74463 74108
rect 74209 74045 74295 74068
rect 74377 74045 74463 74068
rect 89329 74108 89415 74131
rect 89497 74108 89583 74131
rect 89329 74068 89354 74108
rect 89354 74068 89394 74108
rect 89394 74068 89415 74108
rect 89497 74068 89518 74108
rect 89518 74068 89558 74108
rect 89558 74068 89583 74108
rect 89329 74045 89415 74068
rect 89497 74045 89583 74068
rect 104449 74108 104535 74131
rect 104617 74108 104703 74131
rect 104449 74068 104474 74108
rect 104474 74068 104514 74108
rect 104514 74068 104535 74108
rect 104617 74068 104638 74108
rect 104638 74068 104678 74108
rect 104678 74068 104703 74108
rect 104449 74045 104535 74068
rect 104617 74045 104703 74068
rect 119569 74108 119655 74131
rect 119737 74108 119823 74131
rect 119569 74068 119594 74108
rect 119594 74068 119634 74108
rect 119634 74068 119655 74108
rect 119737 74068 119758 74108
rect 119758 74068 119798 74108
rect 119798 74068 119823 74108
rect 119569 74045 119655 74068
rect 119737 74045 119823 74068
rect 134689 74108 134775 74131
rect 134857 74108 134943 74131
rect 134689 74068 134714 74108
rect 134714 74068 134754 74108
rect 134754 74068 134775 74108
rect 134857 74068 134878 74108
rect 134878 74068 134918 74108
rect 134918 74068 134943 74108
rect 134689 74045 134775 74068
rect 134857 74045 134943 74068
rect 149809 74108 149895 74131
rect 149977 74108 150063 74131
rect 149809 74068 149834 74108
rect 149834 74068 149874 74108
rect 149874 74068 149895 74108
rect 149977 74068 149998 74108
rect 149998 74068 150038 74108
rect 150038 74068 150063 74108
rect 149809 74045 149895 74068
rect 149977 74045 150063 74068
rect 75449 73352 75535 73375
rect 75617 73352 75703 73375
rect 75449 73312 75474 73352
rect 75474 73312 75514 73352
rect 75514 73312 75535 73352
rect 75617 73312 75638 73352
rect 75638 73312 75678 73352
rect 75678 73312 75703 73352
rect 75449 73289 75535 73312
rect 75617 73289 75703 73312
rect 90569 73352 90655 73375
rect 90737 73352 90823 73375
rect 90569 73312 90594 73352
rect 90594 73312 90634 73352
rect 90634 73312 90655 73352
rect 90737 73312 90758 73352
rect 90758 73312 90798 73352
rect 90798 73312 90823 73352
rect 90569 73289 90655 73312
rect 90737 73289 90823 73312
rect 105689 73352 105775 73375
rect 105857 73352 105943 73375
rect 105689 73312 105714 73352
rect 105714 73312 105754 73352
rect 105754 73312 105775 73352
rect 105857 73312 105878 73352
rect 105878 73312 105918 73352
rect 105918 73312 105943 73352
rect 105689 73289 105775 73312
rect 105857 73289 105943 73312
rect 120809 73352 120895 73375
rect 120977 73352 121063 73375
rect 120809 73312 120834 73352
rect 120834 73312 120874 73352
rect 120874 73312 120895 73352
rect 120977 73312 120998 73352
rect 120998 73312 121038 73352
rect 121038 73312 121063 73352
rect 120809 73289 120895 73312
rect 120977 73289 121063 73312
rect 135929 73352 136015 73375
rect 136097 73352 136183 73375
rect 135929 73312 135954 73352
rect 135954 73312 135994 73352
rect 135994 73312 136015 73352
rect 136097 73312 136118 73352
rect 136118 73312 136158 73352
rect 136158 73312 136183 73352
rect 135929 73289 136015 73312
rect 136097 73289 136183 73312
rect 151049 73352 151135 73375
rect 151217 73352 151303 73375
rect 151049 73312 151074 73352
rect 151074 73312 151114 73352
rect 151114 73312 151135 73352
rect 151217 73312 151238 73352
rect 151238 73312 151278 73352
rect 151278 73312 151303 73352
rect 151049 73289 151135 73312
rect 151217 73289 151303 73312
rect 74209 72596 74295 72619
rect 74377 72596 74463 72619
rect 74209 72556 74234 72596
rect 74234 72556 74274 72596
rect 74274 72556 74295 72596
rect 74377 72556 74398 72596
rect 74398 72556 74438 72596
rect 74438 72556 74463 72596
rect 74209 72533 74295 72556
rect 74377 72533 74463 72556
rect 89329 72596 89415 72619
rect 89497 72596 89583 72619
rect 89329 72556 89354 72596
rect 89354 72556 89394 72596
rect 89394 72556 89415 72596
rect 89497 72556 89518 72596
rect 89518 72556 89558 72596
rect 89558 72556 89583 72596
rect 89329 72533 89415 72556
rect 89497 72533 89583 72556
rect 104449 72596 104535 72619
rect 104617 72596 104703 72619
rect 104449 72556 104474 72596
rect 104474 72556 104514 72596
rect 104514 72556 104535 72596
rect 104617 72556 104638 72596
rect 104638 72556 104678 72596
rect 104678 72556 104703 72596
rect 104449 72533 104535 72556
rect 104617 72533 104703 72556
rect 119569 72596 119655 72619
rect 119737 72596 119823 72619
rect 119569 72556 119594 72596
rect 119594 72556 119634 72596
rect 119634 72556 119655 72596
rect 119737 72556 119758 72596
rect 119758 72556 119798 72596
rect 119798 72556 119823 72596
rect 119569 72533 119655 72556
rect 119737 72533 119823 72556
rect 134689 72596 134775 72619
rect 134857 72596 134943 72619
rect 134689 72556 134714 72596
rect 134714 72556 134754 72596
rect 134754 72556 134775 72596
rect 134857 72556 134878 72596
rect 134878 72556 134918 72596
rect 134918 72556 134943 72596
rect 134689 72533 134775 72556
rect 134857 72533 134943 72556
rect 149809 72596 149895 72619
rect 149977 72596 150063 72619
rect 149809 72556 149834 72596
rect 149834 72556 149874 72596
rect 149874 72556 149895 72596
rect 149977 72556 149998 72596
rect 149998 72556 150038 72596
rect 150038 72556 150063 72596
rect 149809 72533 149895 72556
rect 149977 72533 150063 72556
rect 75449 71840 75535 71863
rect 75617 71840 75703 71863
rect 75449 71800 75474 71840
rect 75474 71800 75514 71840
rect 75514 71800 75535 71840
rect 75617 71800 75638 71840
rect 75638 71800 75678 71840
rect 75678 71800 75703 71840
rect 75449 71777 75535 71800
rect 75617 71777 75703 71800
rect 90569 71840 90655 71863
rect 90737 71840 90823 71863
rect 90569 71800 90594 71840
rect 90594 71800 90634 71840
rect 90634 71800 90655 71840
rect 90737 71800 90758 71840
rect 90758 71800 90798 71840
rect 90798 71800 90823 71840
rect 90569 71777 90655 71800
rect 90737 71777 90823 71800
rect 105689 71840 105775 71863
rect 105857 71840 105943 71863
rect 105689 71800 105714 71840
rect 105714 71800 105754 71840
rect 105754 71800 105775 71840
rect 105857 71800 105878 71840
rect 105878 71800 105918 71840
rect 105918 71800 105943 71840
rect 105689 71777 105775 71800
rect 105857 71777 105943 71800
rect 120809 71840 120895 71863
rect 120977 71840 121063 71863
rect 120809 71800 120834 71840
rect 120834 71800 120874 71840
rect 120874 71800 120895 71840
rect 120977 71800 120998 71840
rect 120998 71800 121038 71840
rect 121038 71800 121063 71840
rect 120809 71777 120895 71800
rect 120977 71777 121063 71800
rect 135929 71840 136015 71863
rect 136097 71840 136183 71863
rect 135929 71800 135954 71840
rect 135954 71800 135994 71840
rect 135994 71800 136015 71840
rect 136097 71800 136118 71840
rect 136118 71800 136158 71840
rect 136158 71800 136183 71840
rect 135929 71777 136015 71800
rect 136097 71777 136183 71800
rect 151049 71840 151135 71863
rect 151217 71840 151303 71863
rect 151049 71800 151074 71840
rect 151074 71800 151114 71840
rect 151114 71800 151135 71840
rect 151217 71800 151238 71840
rect 151238 71800 151278 71840
rect 151278 71800 151303 71840
rect 151049 71777 151135 71800
rect 151217 71777 151303 71800
<< metal6 >>
rect 82666 167958 85332 168000
rect 82666 167578 82829 167958
rect 83209 167578 83221 167958
rect 83601 167578 83613 167958
rect 83993 167578 84005 167958
rect 84385 167578 84397 167958
rect 84777 167578 84789 167958
rect 85169 167578 85332 167958
rect 82666 167566 85332 167578
rect 82666 167186 82829 167566
rect 83209 167186 83221 167566
rect 83601 167186 83613 167566
rect 83993 167186 84005 167566
rect 84385 167186 84397 167566
rect 84777 167186 84789 167566
rect 85169 167186 85332 167566
rect 82666 167174 85332 167186
rect 82666 166794 82829 167174
rect 83209 166794 83221 167174
rect 83601 166794 83613 167174
rect 83993 166794 84005 167174
rect 84385 166794 84397 167174
rect 84777 166794 84789 167174
rect 85169 166794 85332 167174
rect 82666 166782 85332 166794
rect 82666 166402 82829 166782
rect 83209 166402 83221 166782
rect 83601 166402 83613 166782
rect 83993 166402 84005 166782
rect 84385 166402 84397 166782
rect 84777 166402 84789 166782
rect 85169 166402 85332 166782
rect 82666 166390 85332 166402
rect 82666 166010 82829 166390
rect 83209 166010 83221 166390
rect 83601 166010 83613 166390
rect 83993 166010 84005 166390
rect 84385 166010 84397 166390
rect 84777 166010 84789 166390
rect 85169 166010 85332 166390
rect 82666 165998 85332 166010
rect 82666 165618 82829 165998
rect 83209 165618 83221 165998
rect 83601 165618 83613 165998
rect 83993 165618 84005 165998
rect 84385 165618 84397 165998
rect 84777 165618 84789 165998
rect 85169 165618 85332 165998
rect 82666 165606 85332 165618
rect 82666 165226 82829 165606
rect 83209 165226 83221 165606
rect 83601 165226 83613 165606
rect 83993 165226 84005 165606
rect 84385 165226 84397 165606
rect 84777 165226 84789 165606
rect 85169 165226 85332 165606
rect 82666 165214 85332 165226
rect 82666 164834 82829 165214
rect 83209 164834 83221 165214
rect 83601 164834 83613 165214
rect 83993 164834 84005 165214
rect 84385 164834 84397 165214
rect 84777 164834 84789 165214
rect 85169 164834 85332 165214
rect 82666 164822 85332 164834
rect 82666 164442 82829 164822
rect 83209 164442 83221 164822
rect 83601 164442 83613 164822
rect 83993 164442 84005 164822
rect 84385 164442 84397 164822
rect 84777 164442 84789 164822
rect 85169 164442 85332 164822
rect 82666 164400 85332 164442
rect 98666 167958 101332 168000
rect 98666 167578 98829 167958
rect 99209 167578 99221 167958
rect 99601 167578 99613 167958
rect 99993 167578 100005 167958
rect 100385 167578 100397 167958
rect 100777 167578 100789 167958
rect 101169 167578 101332 167958
rect 98666 167566 101332 167578
rect 98666 167186 98829 167566
rect 99209 167186 99221 167566
rect 99601 167186 99613 167566
rect 99993 167186 100005 167566
rect 100385 167186 100397 167566
rect 100777 167186 100789 167566
rect 101169 167186 101332 167566
rect 98666 167174 101332 167186
rect 98666 166794 98829 167174
rect 99209 166794 99221 167174
rect 99601 166794 99613 167174
rect 99993 166794 100005 167174
rect 100385 166794 100397 167174
rect 100777 166794 100789 167174
rect 101169 166794 101332 167174
rect 98666 166782 101332 166794
rect 98666 166402 98829 166782
rect 99209 166402 99221 166782
rect 99601 166402 99613 166782
rect 99993 166402 100005 166782
rect 100385 166402 100397 166782
rect 100777 166402 100789 166782
rect 101169 166402 101332 166782
rect 98666 166390 101332 166402
rect 98666 166010 98829 166390
rect 99209 166010 99221 166390
rect 99601 166010 99613 166390
rect 99993 166010 100005 166390
rect 100385 166010 100397 166390
rect 100777 166010 100789 166390
rect 101169 166010 101332 166390
rect 98666 165998 101332 166010
rect 98666 165618 98829 165998
rect 99209 165618 99221 165998
rect 99601 165618 99613 165998
rect 99993 165618 100005 165998
rect 100385 165618 100397 165998
rect 100777 165618 100789 165998
rect 101169 165618 101332 165998
rect 98666 165606 101332 165618
rect 98666 165226 98829 165606
rect 99209 165226 99221 165606
rect 99601 165226 99613 165606
rect 99993 165226 100005 165606
rect 100385 165226 100397 165606
rect 100777 165226 100789 165606
rect 101169 165226 101332 165606
rect 98666 165214 101332 165226
rect 98666 164834 98829 165214
rect 99209 164834 99221 165214
rect 99601 164834 99613 165214
rect 99993 164834 100005 165214
rect 100385 164834 100397 165214
rect 100777 164834 100789 165214
rect 101169 164834 101332 165214
rect 98666 164822 101332 164834
rect 98666 164442 98829 164822
rect 99209 164442 99221 164822
rect 99601 164442 99613 164822
rect 99993 164442 100005 164822
rect 100385 164442 100397 164822
rect 100777 164442 100789 164822
rect 101169 164442 101332 164822
rect 98666 164400 101332 164442
rect 114666 167958 117332 168000
rect 114666 167578 114829 167958
rect 115209 167578 115221 167958
rect 115601 167578 115613 167958
rect 115993 167578 116005 167958
rect 116385 167578 116397 167958
rect 116777 167578 116789 167958
rect 117169 167578 117332 167958
rect 114666 167566 117332 167578
rect 114666 167186 114829 167566
rect 115209 167186 115221 167566
rect 115601 167186 115613 167566
rect 115993 167186 116005 167566
rect 116385 167186 116397 167566
rect 116777 167186 116789 167566
rect 117169 167186 117332 167566
rect 114666 167174 117332 167186
rect 114666 166794 114829 167174
rect 115209 166794 115221 167174
rect 115601 166794 115613 167174
rect 115993 166794 116005 167174
rect 116385 166794 116397 167174
rect 116777 166794 116789 167174
rect 117169 166794 117332 167174
rect 114666 166782 117332 166794
rect 114666 166402 114829 166782
rect 115209 166402 115221 166782
rect 115601 166402 115613 166782
rect 115993 166402 116005 166782
rect 116385 166402 116397 166782
rect 116777 166402 116789 166782
rect 117169 166402 117332 166782
rect 114666 166390 117332 166402
rect 114666 166010 114829 166390
rect 115209 166010 115221 166390
rect 115601 166010 115613 166390
rect 115993 166010 116005 166390
rect 116385 166010 116397 166390
rect 116777 166010 116789 166390
rect 117169 166010 117332 166390
rect 114666 165998 117332 166010
rect 114666 165618 114829 165998
rect 115209 165618 115221 165998
rect 115601 165618 115613 165998
rect 115993 165618 116005 165998
rect 116385 165618 116397 165998
rect 116777 165618 116789 165998
rect 117169 165618 117332 165998
rect 114666 165606 117332 165618
rect 114666 165226 114829 165606
rect 115209 165226 115221 165606
rect 115601 165226 115613 165606
rect 115993 165226 116005 165606
rect 116385 165226 116397 165606
rect 116777 165226 116789 165606
rect 117169 165226 117332 165606
rect 114666 165214 117332 165226
rect 114666 164834 114829 165214
rect 115209 164834 115221 165214
rect 115601 164834 115613 165214
rect 115993 164834 116005 165214
rect 116385 164834 116397 165214
rect 116777 164834 116789 165214
rect 117169 164834 117332 165214
rect 114666 164822 117332 164834
rect 114666 164442 114829 164822
rect 115209 164442 115221 164822
rect 115601 164442 115613 164822
rect 115993 164442 116005 164822
rect 116385 164442 116397 164822
rect 116777 164442 116789 164822
rect 117169 164442 117332 164822
rect 114666 164400 117332 164442
rect 130666 167958 133332 168000
rect 130666 167578 130829 167958
rect 131209 167578 131221 167958
rect 131601 167578 131613 167958
rect 131993 167578 132005 167958
rect 132385 167578 132397 167958
rect 132777 167578 132789 167958
rect 133169 167578 133332 167958
rect 130666 167566 133332 167578
rect 130666 167186 130829 167566
rect 131209 167186 131221 167566
rect 131601 167186 131613 167566
rect 131993 167186 132005 167566
rect 132385 167186 132397 167566
rect 132777 167186 132789 167566
rect 133169 167186 133332 167566
rect 130666 167174 133332 167186
rect 130666 166794 130829 167174
rect 131209 166794 131221 167174
rect 131601 166794 131613 167174
rect 131993 166794 132005 167174
rect 132385 166794 132397 167174
rect 132777 166794 132789 167174
rect 133169 166794 133332 167174
rect 130666 166782 133332 166794
rect 130666 166402 130829 166782
rect 131209 166402 131221 166782
rect 131601 166402 131613 166782
rect 131993 166402 132005 166782
rect 132385 166402 132397 166782
rect 132777 166402 132789 166782
rect 133169 166402 133332 166782
rect 130666 166390 133332 166402
rect 130666 166010 130829 166390
rect 131209 166010 131221 166390
rect 131601 166010 131613 166390
rect 131993 166010 132005 166390
rect 132385 166010 132397 166390
rect 132777 166010 132789 166390
rect 133169 166010 133332 166390
rect 130666 165998 133332 166010
rect 130666 165618 130829 165998
rect 131209 165618 131221 165998
rect 131601 165618 131613 165998
rect 131993 165618 132005 165998
rect 132385 165618 132397 165998
rect 132777 165618 132789 165998
rect 133169 165618 133332 165998
rect 130666 165606 133332 165618
rect 130666 165226 130829 165606
rect 131209 165226 131221 165606
rect 131601 165226 131613 165606
rect 131993 165226 132005 165606
rect 132385 165226 132397 165606
rect 132777 165226 132789 165606
rect 133169 165226 133332 165606
rect 130666 165214 133332 165226
rect 130666 164834 130829 165214
rect 131209 164834 131221 165214
rect 131601 164834 131613 165214
rect 131993 164834 132005 165214
rect 132385 164834 132397 165214
rect 132777 164834 132789 165214
rect 133169 164834 133332 165214
rect 130666 164822 133332 164834
rect 130666 164442 130829 164822
rect 131209 164442 131221 164822
rect 131601 164442 131613 164822
rect 131993 164442 132005 164822
rect 132385 164442 132397 164822
rect 132777 164442 132789 164822
rect 133169 164442 133332 164822
rect 130666 164400 133332 164442
rect 146666 167958 149332 168000
rect 146666 167578 146829 167958
rect 147209 167578 147221 167958
rect 147601 167578 147613 167958
rect 147993 167578 148005 167958
rect 148385 167578 148397 167958
rect 148777 167578 148789 167958
rect 149169 167578 149332 167958
rect 146666 167566 149332 167578
rect 146666 167186 146829 167566
rect 147209 167186 147221 167566
rect 147601 167186 147613 167566
rect 147993 167186 148005 167566
rect 148385 167186 148397 167566
rect 148777 167186 148789 167566
rect 149169 167186 149332 167566
rect 146666 167174 149332 167186
rect 146666 166794 146829 167174
rect 147209 166794 147221 167174
rect 147601 166794 147613 167174
rect 147993 166794 148005 167174
rect 148385 166794 148397 167174
rect 148777 166794 148789 167174
rect 149169 166794 149332 167174
rect 146666 166782 149332 166794
rect 146666 166402 146829 166782
rect 147209 166402 147221 166782
rect 147601 166402 147613 166782
rect 147993 166402 148005 166782
rect 148385 166402 148397 166782
rect 148777 166402 148789 166782
rect 149169 166402 149332 166782
rect 146666 166390 149332 166402
rect 146666 166010 146829 166390
rect 147209 166010 147221 166390
rect 147601 166010 147613 166390
rect 147993 166010 148005 166390
rect 148385 166010 148397 166390
rect 148777 166010 148789 166390
rect 149169 166010 149332 166390
rect 146666 165998 149332 166010
rect 146666 165618 146829 165998
rect 147209 165618 147221 165998
rect 147601 165618 147613 165998
rect 147993 165618 148005 165998
rect 148385 165618 148397 165998
rect 148777 165618 148789 165998
rect 149169 165618 149332 165998
rect 146666 165606 149332 165618
rect 146666 165226 146829 165606
rect 147209 165226 147221 165606
rect 147601 165226 147613 165606
rect 147993 165226 148005 165606
rect 148385 165226 148397 165606
rect 148777 165226 148789 165606
rect 149169 165226 149332 165606
rect 146666 165214 149332 165226
rect 146666 164834 146829 165214
rect 147209 164834 147221 165214
rect 147601 164834 147613 165214
rect 147993 164834 148005 165214
rect 148385 164834 148397 165214
rect 148777 164834 148789 165214
rect 149169 164834 149332 165214
rect 146666 164822 149332 164834
rect 146666 164442 146829 164822
rect 147209 164442 147221 164822
rect 147601 164442 147613 164822
rect 147993 164442 148005 164822
rect 148385 164442 148397 164822
rect 148777 164442 148789 164822
rect 149169 164442 149332 164822
rect 146666 164400 149332 164442
rect 71998 163958 74664 164000
rect 71998 163578 72161 163958
rect 72541 163578 72553 163958
rect 72933 163578 72945 163958
rect 73325 163578 73337 163958
rect 73717 163578 73729 163958
rect 74109 163578 74121 163958
rect 74501 163578 74664 163958
rect 71998 163566 74664 163578
rect 71998 163186 72161 163566
rect 72541 163186 72553 163566
rect 72933 163186 72945 163566
rect 73325 163186 73337 163566
rect 73717 163186 73729 163566
rect 74109 163186 74121 163566
rect 74501 163186 74664 163566
rect 71998 163174 74664 163186
rect 71998 162794 72161 163174
rect 72541 162794 72553 163174
rect 72933 162794 72945 163174
rect 73325 162794 73337 163174
rect 73717 162794 73729 163174
rect 74109 162794 74121 163174
rect 74501 162794 74664 163174
rect 71998 162782 74664 162794
rect 71998 162402 72161 162782
rect 72541 162402 72553 162782
rect 72933 162402 72945 162782
rect 73325 162402 73337 162782
rect 73717 162402 73729 162782
rect 74109 162402 74121 162782
rect 74501 162402 74664 162782
rect 71998 162390 74664 162402
rect 71998 162010 72161 162390
rect 72541 162010 72553 162390
rect 72933 162010 72945 162390
rect 73325 162010 73337 162390
rect 73717 162010 73729 162390
rect 74109 162010 74121 162390
rect 74501 162010 74664 162390
rect 71998 161998 74664 162010
rect 71998 161618 72161 161998
rect 72541 161618 72553 161998
rect 72933 161618 72945 161998
rect 73325 161618 73337 161998
rect 73717 161618 73729 161998
rect 74109 161618 74121 161998
rect 74501 161618 74664 161998
rect 71998 161606 74664 161618
rect 71998 161226 72161 161606
rect 72541 161226 72553 161606
rect 72933 161226 72945 161606
rect 73325 161226 73337 161606
rect 73717 161226 73729 161606
rect 74109 161226 74121 161606
rect 74501 161226 74664 161606
rect 71998 161214 74664 161226
rect 71998 160834 72161 161214
rect 72541 160834 72553 161214
rect 72933 160834 72945 161214
rect 73325 160834 73337 161214
rect 73717 160834 73729 161214
rect 74109 160834 74121 161214
rect 74501 160834 74664 161214
rect 71998 160822 74664 160834
rect 71998 160442 72161 160822
rect 72541 160442 72553 160822
rect 72933 160442 72945 160822
rect 73325 160442 73337 160822
rect 73717 160442 73729 160822
rect 74109 160442 74121 160822
rect 74501 160442 74664 160822
rect 71998 160400 74664 160442
rect 87998 163958 90664 164000
rect 87998 163578 88161 163958
rect 88541 163578 88553 163958
rect 88933 163578 88945 163958
rect 89325 163578 89337 163958
rect 89717 163578 89729 163958
rect 90109 163578 90121 163958
rect 90501 163578 90664 163958
rect 87998 163566 90664 163578
rect 87998 163186 88161 163566
rect 88541 163186 88553 163566
rect 88933 163186 88945 163566
rect 89325 163186 89337 163566
rect 89717 163186 89729 163566
rect 90109 163186 90121 163566
rect 90501 163186 90664 163566
rect 87998 163174 90664 163186
rect 87998 162794 88161 163174
rect 88541 162794 88553 163174
rect 88933 162794 88945 163174
rect 89325 162794 89337 163174
rect 89717 162794 89729 163174
rect 90109 162794 90121 163174
rect 90501 162794 90664 163174
rect 87998 162782 90664 162794
rect 87998 162402 88161 162782
rect 88541 162402 88553 162782
rect 88933 162402 88945 162782
rect 89325 162402 89337 162782
rect 89717 162402 89729 162782
rect 90109 162402 90121 162782
rect 90501 162402 90664 162782
rect 87998 162390 90664 162402
rect 87998 162010 88161 162390
rect 88541 162010 88553 162390
rect 88933 162010 88945 162390
rect 89325 162010 89337 162390
rect 89717 162010 89729 162390
rect 90109 162010 90121 162390
rect 90501 162010 90664 162390
rect 87998 161998 90664 162010
rect 87998 161618 88161 161998
rect 88541 161618 88553 161998
rect 88933 161618 88945 161998
rect 89325 161618 89337 161998
rect 89717 161618 89729 161998
rect 90109 161618 90121 161998
rect 90501 161618 90664 161998
rect 87998 161606 90664 161618
rect 87998 161226 88161 161606
rect 88541 161226 88553 161606
rect 88933 161226 88945 161606
rect 89325 161226 89337 161606
rect 89717 161226 89729 161606
rect 90109 161226 90121 161606
rect 90501 161226 90664 161606
rect 87998 161214 90664 161226
rect 87998 160834 88161 161214
rect 88541 160834 88553 161214
rect 88933 160834 88945 161214
rect 89325 160834 89337 161214
rect 89717 160834 89729 161214
rect 90109 160834 90121 161214
rect 90501 160834 90664 161214
rect 87998 160822 90664 160834
rect 87998 160442 88161 160822
rect 88541 160442 88553 160822
rect 88933 160442 88945 160822
rect 89325 160442 89337 160822
rect 89717 160442 89729 160822
rect 90109 160442 90121 160822
rect 90501 160442 90664 160822
rect 87998 160400 90664 160442
rect 103998 163958 106664 164000
rect 103998 163578 104161 163958
rect 104541 163578 104553 163958
rect 104933 163578 104945 163958
rect 105325 163578 105337 163958
rect 105717 163578 105729 163958
rect 106109 163578 106121 163958
rect 106501 163578 106664 163958
rect 103998 163566 106664 163578
rect 103998 163186 104161 163566
rect 104541 163186 104553 163566
rect 104933 163186 104945 163566
rect 105325 163186 105337 163566
rect 105717 163186 105729 163566
rect 106109 163186 106121 163566
rect 106501 163186 106664 163566
rect 103998 163174 106664 163186
rect 103998 162794 104161 163174
rect 104541 162794 104553 163174
rect 104933 162794 104945 163174
rect 105325 162794 105337 163174
rect 105717 162794 105729 163174
rect 106109 162794 106121 163174
rect 106501 162794 106664 163174
rect 103998 162782 106664 162794
rect 103998 162402 104161 162782
rect 104541 162402 104553 162782
rect 104933 162402 104945 162782
rect 105325 162402 105337 162782
rect 105717 162402 105729 162782
rect 106109 162402 106121 162782
rect 106501 162402 106664 162782
rect 103998 162390 106664 162402
rect 103998 162010 104161 162390
rect 104541 162010 104553 162390
rect 104933 162010 104945 162390
rect 105325 162010 105337 162390
rect 105717 162010 105729 162390
rect 106109 162010 106121 162390
rect 106501 162010 106664 162390
rect 103998 161998 106664 162010
rect 103998 161618 104161 161998
rect 104541 161618 104553 161998
rect 104933 161618 104945 161998
rect 105325 161618 105337 161998
rect 105717 161618 105729 161998
rect 106109 161618 106121 161998
rect 106501 161618 106664 161998
rect 103998 161606 106664 161618
rect 103998 161226 104161 161606
rect 104541 161226 104553 161606
rect 104933 161226 104945 161606
rect 105325 161226 105337 161606
rect 105717 161226 105729 161606
rect 106109 161226 106121 161606
rect 106501 161226 106664 161606
rect 103998 161214 106664 161226
rect 103998 160834 104161 161214
rect 104541 160834 104553 161214
rect 104933 160834 104945 161214
rect 105325 160834 105337 161214
rect 105717 160834 105729 161214
rect 106109 160834 106121 161214
rect 106501 160834 106664 161214
rect 103998 160822 106664 160834
rect 103998 160442 104161 160822
rect 104541 160442 104553 160822
rect 104933 160442 104945 160822
rect 105325 160442 105337 160822
rect 105717 160442 105729 160822
rect 106109 160442 106121 160822
rect 106501 160442 106664 160822
rect 103998 160400 106664 160442
rect 119998 163958 122664 164000
rect 119998 163578 120161 163958
rect 120541 163578 120553 163958
rect 120933 163578 120945 163958
rect 121325 163578 121337 163958
rect 121717 163578 121729 163958
rect 122109 163578 122121 163958
rect 122501 163578 122664 163958
rect 119998 163566 122664 163578
rect 119998 163186 120161 163566
rect 120541 163186 120553 163566
rect 120933 163186 120945 163566
rect 121325 163186 121337 163566
rect 121717 163186 121729 163566
rect 122109 163186 122121 163566
rect 122501 163186 122664 163566
rect 119998 163174 122664 163186
rect 119998 162794 120161 163174
rect 120541 162794 120553 163174
rect 120933 162794 120945 163174
rect 121325 162794 121337 163174
rect 121717 162794 121729 163174
rect 122109 162794 122121 163174
rect 122501 162794 122664 163174
rect 119998 162782 122664 162794
rect 119998 162402 120161 162782
rect 120541 162402 120553 162782
rect 120933 162402 120945 162782
rect 121325 162402 121337 162782
rect 121717 162402 121729 162782
rect 122109 162402 122121 162782
rect 122501 162402 122664 162782
rect 119998 162390 122664 162402
rect 119998 162010 120161 162390
rect 120541 162010 120553 162390
rect 120933 162010 120945 162390
rect 121325 162010 121337 162390
rect 121717 162010 121729 162390
rect 122109 162010 122121 162390
rect 122501 162010 122664 162390
rect 119998 161998 122664 162010
rect 119998 161618 120161 161998
rect 120541 161618 120553 161998
rect 120933 161618 120945 161998
rect 121325 161618 121337 161998
rect 121717 161618 121729 161998
rect 122109 161618 122121 161998
rect 122501 161618 122664 161998
rect 119998 161606 122664 161618
rect 119998 161226 120161 161606
rect 120541 161226 120553 161606
rect 120933 161226 120945 161606
rect 121325 161226 121337 161606
rect 121717 161226 121729 161606
rect 122109 161226 122121 161606
rect 122501 161226 122664 161606
rect 119998 161214 122664 161226
rect 119998 160834 120161 161214
rect 120541 160834 120553 161214
rect 120933 160834 120945 161214
rect 121325 160834 121337 161214
rect 121717 160834 121729 161214
rect 122109 160834 122121 161214
rect 122501 160834 122664 161214
rect 119998 160822 122664 160834
rect 119998 160442 120161 160822
rect 120541 160442 120553 160822
rect 120933 160442 120945 160822
rect 121325 160442 121337 160822
rect 121717 160442 121729 160822
rect 122109 160442 122121 160822
rect 122501 160442 122664 160822
rect 119998 160400 122664 160442
rect 135998 163958 138664 164000
rect 135998 163578 136161 163958
rect 136541 163578 136553 163958
rect 136933 163578 136945 163958
rect 137325 163578 137337 163958
rect 137717 163578 137729 163958
rect 138109 163578 138121 163958
rect 138501 163578 138664 163958
rect 135998 163566 138664 163578
rect 135998 163186 136161 163566
rect 136541 163186 136553 163566
rect 136933 163186 136945 163566
rect 137325 163186 137337 163566
rect 137717 163186 137729 163566
rect 138109 163186 138121 163566
rect 138501 163186 138664 163566
rect 135998 163174 138664 163186
rect 135998 162794 136161 163174
rect 136541 162794 136553 163174
rect 136933 162794 136945 163174
rect 137325 162794 137337 163174
rect 137717 162794 137729 163174
rect 138109 162794 138121 163174
rect 138501 162794 138664 163174
rect 135998 162782 138664 162794
rect 135998 162402 136161 162782
rect 136541 162402 136553 162782
rect 136933 162402 136945 162782
rect 137325 162402 137337 162782
rect 137717 162402 137729 162782
rect 138109 162402 138121 162782
rect 138501 162402 138664 162782
rect 135998 162390 138664 162402
rect 135998 162010 136161 162390
rect 136541 162010 136553 162390
rect 136933 162010 136945 162390
rect 137325 162010 137337 162390
rect 137717 162010 137729 162390
rect 138109 162010 138121 162390
rect 138501 162010 138664 162390
rect 135998 161998 138664 162010
rect 135998 161618 136161 161998
rect 136541 161618 136553 161998
rect 136933 161618 136945 161998
rect 137325 161618 137337 161998
rect 137717 161618 137729 161998
rect 138109 161618 138121 161998
rect 138501 161618 138664 161998
rect 135998 161606 138664 161618
rect 135998 161226 136161 161606
rect 136541 161226 136553 161606
rect 136933 161226 136945 161606
rect 137325 161226 137337 161606
rect 137717 161226 137729 161606
rect 138109 161226 138121 161606
rect 138501 161226 138664 161606
rect 135998 161214 138664 161226
rect 135998 160834 136161 161214
rect 136541 160834 136553 161214
rect 136933 160834 136945 161214
rect 137325 160834 137337 161214
rect 137717 160834 137729 161214
rect 138109 160834 138121 161214
rect 138501 160834 138664 161214
rect 135998 160822 138664 160834
rect 135998 160442 136161 160822
rect 136541 160442 136553 160822
rect 136933 160442 136945 160822
rect 137325 160442 137337 160822
rect 137717 160442 137729 160822
rect 138109 160442 138121 160822
rect 138501 160442 138664 160822
rect 135998 160400 138664 160442
rect 151998 163958 154664 164000
rect 151998 163578 152161 163958
rect 152541 163578 152553 163958
rect 152933 163578 152945 163958
rect 153325 163578 153337 163958
rect 153717 163578 153729 163958
rect 154109 163578 154121 163958
rect 154501 163578 154664 163958
rect 151998 163566 154664 163578
rect 151998 163186 152161 163566
rect 152541 163186 152553 163566
rect 152933 163186 152945 163566
rect 153325 163186 153337 163566
rect 153717 163186 153729 163566
rect 154109 163186 154121 163566
rect 154501 163186 154664 163566
rect 151998 163174 154664 163186
rect 151998 162794 152161 163174
rect 152541 162794 152553 163174
rect 152933 162794 152945 163174
rect 153325 162794 153337 163174
rect 153717 162794 153729 163174
rect 154109 162794 154121 163174
rect 154501 162794 154664 163174
rect 151998 162782 154664 162794
rect 151998 162402 152161 162782
rect 152541 162402 152553 162782
rect 152933 162402 152945 162782
rect 153325 162402 153337 162782
rect 153717 162402 153729 162782
rect 154109 162402 154121 162782
rect 154501 162402 154664 162782
rect 151998 162390 154664 162402
rect 151998 162010 152161 162390
rect 152541 162010 152553 162390
rect 152933 162010 152945 162390
rect 153325 162010 153337 162390
rect 153717 162010 153729 162390
rect 154109 162010 154121 162390
rect 154501 162010 154664 162390
rect 151998 161998 154664 162010
rect 151998 161618 152161 161998
rect 152541 161618 152553 161998
rect 152933 161618 152945 161998
rect 153325 161618 153337 161998
rect 153717 161618 153729 161998
rect 154109 161618 154121 161998
rect 154501 161618 154664 161998
rect 151998 161606 154664 161618
rect 151998 161226 152161 161606
rect 152541 161226 152553 161606
rect 152933 161226 152945 161606
rect 153325 161226 153337 161606
rect 153717 161226 153729 161606
rect 154109 161226 154121 161606
rect 154501 161226 154664 161606
rect 151998 161214 154664 161226
rect 151998 160834 152161 161214
rect 152541 160834 152553 161214
rect 152933 160834 152945 161214
rect 153325 160834 153337 161214
rect 153717 160834 153729 161214
rect 154109 160834 154121 161214
rect 154501 160834 154664 161214
rect 151998 160822 154664 160834
rect 151998 160442 152161 160822
rect 152541 160442 152553 160822
rect 152933 160442 152945 160822
rect 153325 160442 153337 160822
rect 153717 160442 153729 160822
rect 154109 160442 154121 160822
rect 154501 160442 154664 160822
rect 151998 160400 154664 160442
rect 68316 155142 69316 155256
rect 68316 154762 68430 155142
rect 68810 154762 68822 155142
rect 69202 154762 69316 155142
rect 68316 154750 69316 154762
rect 60000 154501 63600 154664
rect 60000 154121 60042 154501
rect 60422 154121 60434 154501
rect 60814 154121 60826 154501
rect 61206 154121 61218 154501
rect 61598 154121 61610 154501
rect 61990 154121 62002 154501
rect 62382 154121 62394 154501
rect 62774 154121 62786 154501
rect 63166 154121 63178 154501
rect 63558 154121 63600 154501
rect 60000 154109 63600 154121
rect 60000 153729 60042 154109
rect 60422 153729 60434 154109
rect 60814 153729 60826 154109
rect 61206 153729 61218 154109
rect 61598 153729 61610 154109
rect 61990 153729 62002 154109
rect 62382 153729 62394 154109
rect 62774 153729 62786 154109
rect 63166 153729 63178 154109
rect 63558 153729 63600 154109
rect 60000 153717 63600 153729
rect 60000 153337 60042 153717
rect 60422 153337 60434 153717
rect 60814 153337 60826 153717
rect 61206 153337 61218 153717
rect 61598 153337 61610 153717
rect 61990 153337 62002 153717
rect 62382 153337 62394 153717
rect 62774 153337 62786 153717
rect 63166 153337 63178 153717
rect 63558 153337 63600 153717
rect 60000 153325 63600 153337
rect 60000 152945 60042 153325
rect 60422 152945 60434 153325
rect 60814 152945 60826 153325
rect 61206 152945 61218 153325
rect 61598 152945 61610 153325
rect 61990 152945 62002 153325
rect 62382 152945 62394 153325
rect 62774 152945 62786 153325
rect 63166 152945 63178 153325
rect 63558 152945 63600 153325
rect 60000 152933 63600 152945
rect 60000 152553 60042 152933
rect 60422 152553 60434 152933
rect 60814 152553 60826 152933
rect 61206 152553 61218 152933
rect 61598 152553 61610 152933
rect 61990 152553 62002 152933
rect 62382 152553 62394 152933
rect 62774 152553 62786 152933
rect 63166 152553 63178 152933
rect 63558 152553 63600 152933
rect 60000 152541 63600 152553
rect 60000 152161 60042 152541
rect 60422 152161 60434 152541
rect 60814 152161 60826 152541
rect 61206 152161 61218 152541
rect 61598 152161 61610 152541
rect 61990 152161 62002 152541
rect 62382 152161 62394 152541
rect 62774 152161 62786 152541
rect 63166 152161 63178 152541
rect 63558 152161 63600 152541
rect 60000 151998 63600 152161
rect 68316 154370 68430 154750
rect 68810 154370 68822 154750
rect 69202 154370 69316 154750
rect 68316 151570 69316 154370
rect 68316 151190 68430 151570
rect 68810 151190 68822 151570
rect 69202 151190 69316 151570
rect 56000 149169 59600 149332
rect 56000 148789 56042 149169
rect 56422 148789 56434 149169
rect 56814 148789 56826 149169
rect 57206 148789 57218 149169
rect 57598 148789 57610 149169
rect 57990 148789 58002 149169
rect 58382 148789 58394 149169
rect 58774 148789 58786 149169
rect 59166 148789 59178 149169
rect 59558 148789 59600 149169
rect 56000 148777 59600 148789
rect 56000 148397 56042 148777
rect 56422 148397 56434 148777
rect 56814 148397 56826 148777
rect 57206 148397 57218 148777
rect 57598 148397 57610 148777
rect 57990 148397 58002 148777
rect 58382 148397 58394 148777
rect 58774 148397 58786 148777
rect 59166 148397 59178 148777
rect 59558 148397 59600 148777
rect 56000 148385 59600 148397
rect 56000 148005 56042 148385
rect 56422 148005 56434 148385
rect 56814 148005 56826 148385
rect 57206 148005 57218 148385
rect 57598 148005 57610 148385
rect 57990 148005 58002 148385
rect 58382 148005 58394 148385
rect 58774 148005 58786 148385
rect 59166 148005 59178 148385
rect 59558 148005 59600 148385
rect 56000 147993 59600 148005
rect 56000 147613 56042 147993
rect 56422 147613 56434 147993
rect 56814 147613 56826 147993
rect 57206 147613 57218 147993
rect 57598 147613 57610 147993
rect 57990 147613 58002 147993
rect 58382 147613 58394 147993
rect 58774 147613 58786 147993
rect 59166 147613 59178 147993
rect 59558 147613 59600 147993
rect 56000 147601 59600 147613
rect 56000 147221 56042 147601
rect 56422 147221 56434 147601
rect 56814 147221 56826 147601
rect 57206 147221 57218 147601
rect 57598 147221 57610 147601
rect 57990 147221 58002 147601
rect 58382 147221 58394 147601
rect 58774 147221 58786 147601
rect 59166 147221 59178 147601
rect 59558 147221 59600 147601
rect 56000 147209 59600 147221
rect 56000 146829 56042 147209
rect 56422 146829 56434 147209
rect 56814 146829 56826 147209
rect 57206 146829 57218 147209
rect 57598 146829 57610 147209
rect 57990 146829 58002 147209
rect 58382 146829 58394 147209
rect 58774 146829 58786 147209
rect 59166 146829 59178 147209
rect 59558 146829 59600 147209
rect 56000 146666 59600 146829
rect 60000 138501 63600 138664
rect 60000 138121 60042 138501
rect 60422 138121 60434 138501
rect 60814 138121 60826 138501
rect 61206 138121 61218 138501
rect 61598 138121 61610 138501
rect 61990 138121 62002 138501
rect 62382 138121 62394 138501
rect 62774 138121 62786 138501
rect 63166 138121 63178 138501
rect 63558 138121 63600 138501
rect 60000 138109 63600 138121
rect 60000 137729 60042 138109
rect 60422 137729 60434 138109
rect 60814 137729 60826 138109
rect 61206 137729 61218 138109
rect 61598 137729 61610 138109
rect 61990 137729 62002 138109
rect 62382 137729 62394 138109
rect 62774 137729 62786 138109
rect 63166 137729 63178 138109
rect 63558 137729 63600 138109
rect 60000 137717 63600 137729
rect 60000 137337 60042 137717
rect 60422 137337 60434 137717
rect 60814 137337 60826 137717
rect 61206 137337 61218 137717
rect 61598 137337 61610 137717
rect 61990 137337 62002 137717
rect 62382 137337 62394 137717
rect 62774 137337 62786 137717
rect 63166 137337 63178 137717
rect 63558 137337 63600 137717
rect 60000 137325 63600 137337
rect 60000 136945 60042 137325
rect 60422 136945 60434 137325
rect 60814 136945 60826 137325
rect 61206 136945 61218 137325
rect 61598 136945 61610 137325
rect 61990 136945 62002 137325
rect 62382 136945 62394 137325
rect 62774 136945 62786 137325
rect 63166 136945 63178 137325
rect 63558 136945 63600 137325
rect 60000 136933 63600 136945
rect 60000 136553 60042 136933
rect 60422 136553 60434 136933
rect 60814 136553 60826 136933
rect 61206 136553 61218 136933
rect 61598 136553 61610 136933
rect 61990 136553 62002 136933
rect 62382 136553 62394 136933
rect 62774 136553 62786 136933
rect 63166 136553 63178 136933
rect 63558 136553 63600 136933
rect 60000 136541 63600 136553
rect 60000 136161 60042 136541
rect 60422 136161 60434 136541
rect 60814 136161 60826 136541
rect 61206 136161 61218 136541
rect 61598 136161 61610 136541
rect 61990 136161 62002 136541
rect 62382 136161 62394 136541
rect 62774 136161 62786 136541
rect 63166 136161 63178 136541
rect 63558 136161 63600 136541
rect 60000 135998 63600 136161
rect 68316 138501 69316 151190
rect 68316 138121 68430 138501
rect 68810 138121 68822 138501
rect 69202 138121 69316 138501
rect 68316 138109 69316 138121
rect 68316 137729 68430 138109
rect 68810 137729 68822 138109
rect 69202 137729 69316 138109
rect 68316 137717 69316 137729
rect 68316 137337 68430 137717
rect 68810 137337 68822 137717
rect 69202 137337 69316 137717
rect 68316 137325 69316 137337
rect 68316 136945 68430 137325
rect 68810 136945 68822 137325
rect 69202 136945 69316 137325
rect 68316 136933 69316 136945
rect 68316 136553 68430 136933
rect 68810 136553 68822 136933
rect 69202 136553 69316 136933
rect 68316 136541 69316 136553
rect 68316 136161 68430 136541
rect 68810 136161 68822 136541
rect 69202 136161 69316 136541
rect 56000 133169 59600 133332
rect 56000 132789 56042 133169
rect 56422 132789 56434 133169
rect 56814 132789 56826 133169
rect 57206 132789 57218 133169
rect 57598 132789 57610 133169
rect 57990 132789 58002 133169
rect 58382 132789 58394 133169
rect 58774 132789 58786 133169
rect 59166 132789 59178 133169
rect 59558 132789 59600 133169
rect 56000 132777 59600 132789
rect 56000 132397 56042 132777
rect 56422 132397 56434 132777
rect 56814 132397 56826 132777
rect 57206 132397 57218 132777
rect 57598 132397 57610 132777
rect 57990 132397 58002 132777
rect 58382 132397 58394 132777
rect 58774 132397 58786 132777
rect 59166 132397 59178 132777
rect 59558 132397 59600 132777
rect 56000 132385 59600 132397
rect 56000 132005 56042 132385
rect 56422 132005 56434 132385
rect 56814 132005 56826 132385
rect 57206 132005 57218 132385
rect 57598 132005 57610 132385
rect 57990 132005 58002 132385
rect 58382 132005 58394 132385
rect 58774 132005 58786 132385
rect 59166 132005 59178 132385
rect 59558 132005 59600 132385
rect 56000 131993 59600 132005
rect 56000 131613 56042 131993
rect 56422 131613 56434 131993
rect 56814 131613 56826 131993
rect 57206 131613 57218 131993
rect 57598 131613 57610 131993
rect 57990 131613 58002 131993
rect 58382 131613 58394 131993
rect 58774 131613 58786 131993
rect 59166 131613 59178 131993
rect 59558 131613 59600 131993
rect 56000 131601 59600 131613
rect 56000 131221 56042 131601
rect 56422 131221 56434 131601
rect 56814 131221 56826 131601
rect 57206 131221 57218 131601
rect 57598 131221 57610 131601
rect 57990 131221 58002 131601
rect 58382 131221 58394 131601
rect 58774 131221 58786 131601
rect 59166 131221 59178 131601
rect 59558 131221 59600 131601
rect 56000 131209 59600 131221
rect 56000 130829 56042 131209
rect 56422 130829 56434 131209
rect 56814 130829 56826 131209
rect 57206 130829 57218 131209
rect 57598 130829 57610 131209
rect 57990 130829 58002 131209
rect 58382 130829 58394 131209
rect 58774 130829 58786 131209
rect 59166 130829 59178 131209
rect 59558 130829 59600 131209
rect 56000 130666 59600 130829
rect 60000 122501 63600 122664
rect 60000 122121 60042 122501
rect 60422 122121 60434 122501
rect 60814 122121 60826 122501
rect 61206 122121 61218 122501
rect 61598 122121 61610 122501
rect 61990 122121 62002 122501
rect 62382 122121 62394 122501
rect 62774 122121 62786 122501
rect 63166 122121 63178 122501
rect 63558 122121 63600 122501
rect 60000 122109 63600 122121
rect 60000 121729 60042 122109
rect 60422 121729 60434 122109
rect 60814 121729 60826 122109
rect 61206 121729 61218 122109
rect 61598 121729 61610 122109
rect 61990 121729 62002 122109
rect 62382 121729 62394 122109
rect 62774 121729 62786 122109
rect 63166 121729 63178 122109
rect 63558 121729 63600 122109
rect 60000 121717 63600 121729
rect 60000 121337 60042 121717
rect 60422 121337 60434 121717
rect 60814 121337 60826 121717
rect 61206 121337 61218 121717
rect 61598 121337 61610 121717
rect 61990 121337 62002 121717
rect 62382 121337 62394 121717
rect 62774 121337 62786 121717
rect 63166 121337 63178 121717
rect 63558 121337 63600 121717
rect 60000 121325 63600 121337
rect 60000 120945 60042 121325
rect 60422 120945 60434 121325
rect 60814 120945 60826 121325
rect 61206 120945 61218 121325
rect 61598 120945 61610 121325
rect 61990 120945 62002 121325
rect 62382 120945 62394 121325
rect 62774 120945 62786 121325
rect 63166 120945 63178 121325
rect 63558 120945 63600 121325
rect 60000 120933 63600 120945
rect 60000 120553 60042 120933
rect 60422 120553 60434 120933
rect 60814 120553 60826 120933
rect 61206 120553 61218 120933
rect 61598 120553 61610 120933
rect 61990 120553 62002 120933
rect 62382 120553 62394 120933
rect 62774 120553 62786 120933
rect 63166 120553 63178 120933
rect 63558 120553 63600 120933
rect 60000 120541 63600 120553
rect 60000 120161 60042 120541
rect 60422 120161 60434 120541
rect 60814 120161 60826 120541
rect 61206 120161 61218 120541
rect 61598 120161 61610 120541
rect 61990 120161 62002 120541
rect 62382 120161 62394 120541
rect 62774 120161 62786 120541
rect 63166 120161 63178 120541
rect 63558 120161 63600 120541
rect 60000 119998 63600 120161
rect 68316 122501 69316 136161
rect 68316 122121 68430 122501
rect 68810 122121 68822 122501
rect 69202 122121 69316 122501
rect 68316 122109 69316 122121
rect 68316 121729 68430 122109
rect 68810 121729 68822 122109
rect 69202 121729 69316 122109
rect 68316 121717 69316 121729
rect 68316 121337 68430 121717
rect 68810 121337 68822 121717
rect 69202 121337 69316 121717
rect 68316 121325 69316 121337
rect 68316 120945 68430 121325
rect 68810 120945 68822 121325
rect 69202 120945 69316 121325
rect 68316 120933 69316 120945
rect 68316 120553 68430 120933
rect 68810 120553 68822 120933
rect 69202 120553 69316 120933
rect 68316 120541 69316 120553
rect 68316 120161 68430 120541
rect 68810 120161 68822 120541
rect 69202 120161 69316 120541
rect 56000 117169 59600 117332
rect 56000 116789 56042 117169
rect 56422 116789 56434 117169
rect 56814 116789 56826 117169
rect 57206 116789 57218 117169
rect 57598 116789 57610 117169
rect 57990 116789 58002 117169
rect 58382 116789 58394 117169
rect 58774 116789 58786 117169
rect 59166 116789 59178 117169
rect 59558 116789 59600 117169
rect 56000 116777 59600 116789
rect 56000 116397 56042 116777
rect 56422 116397 56434 116777
rect 56814 116397 56826 116777
rect 57206 116397 57218 116777
rect 57598 116397 57610 116777
rect 57990 116397 58002 116777
rect 58382 116397 58394 116777
rect 58774 116397 58786 116777
rect 59166 116397 59178 116777
rect 59558 116397 59600 116777
rect 56000 116385 59600 116397
rect 56000 116005 56042 116385
rect 56422 116005 56434 116385
rect 56814 116005 56826 116385
rect 57206 116005 57218 116385
rect 57598 116005 57610 116385
rect 57990 116005 58002 116385
rect 58382 116005 58394 116385
rect 58774 116005 58786 116385
rect 59166 116005 59178 116385
rect 59558 116005 59600 116385
rect 56000 115993 59600 116005
rect 56000 115613 56042 115993
rect 56422 115613 56434 115993
rect 56814 115613 56826 115993
rect 57206 115613 57218 115993
rect 57598 115613 57610 115993
rect 57990 115613 58002 115993
rect 58382 115613 58394 115993
rect 58774 115613 58786 115993
rect 59166 115613 59178 115993
rect 59558 115613 59600 115993
rect 56000 115601 59600 115613
rect 56000 115221 56042 115601
rect 56422 115221 56434 115601
rect 56814 115221 56826 115601
rect 57206 115221 57218 115601
rect 57598 115221 57610 115601
rect 57990 115221 58002 115601
rect 58382 115221 58394 115601
rect 58774 115221 58786 115601
rect 59166 115221 59178 115601
rect 59558 115221 59600 115601
rect 56000 115209 59600 115221
rect 56000 114829 56042 115209
rect 56422 114829 56434 115209
rect 56814 114829 56826 115209
rect 57206 114829 57218 115209
rect 57598 114829 57610 115209
rect 57990 114829 58002 115209
rect 58382 114829 58394 115209
rect 58774 114829 58786 115209
rect 59166 114829 59178 115209
rect 59558 114829 59600 115209
rect 56000 114666 59600 114829
rect 60000 106501 63600 106664
rect 60000 106121 60042 106501
rect 60422 106121 60434 106501
rect 60814 106121 60826 106501
rect 61206 106121 61218 106501
rect 61598 106121 61610 106501
rect 61990 106121 62002 106501
rect 62382 106121 62394 106501
rect 62774 106121 62786 106501
rect 63166 106121 63178 106501
rect 63558 106121 63600 106501
rect 60000 106109 63600 106121
rect 60000 105729 60042 106109
rect 60422 105729 60434 106109
rect 60814 105729 60826 106109
rect 61206 105729 61218 106109
rect 61598 105729 61610 106109
rect 61990 105729 62002 106109
rect 62382 105729 62394 106109
rect 62774 105729 62786 106109
rect 63166 105729 63178 106109
rect 63558 105729 63600 106109
rect 60000 105717 63600 105729
rect 60000 105337 60042 105717
rect 60422 105337 60434 105717
rect 60814 105337 60826 105717
rect 61206 105337 61218 105717
rect 61598 105337 61610 105717
rect 61990 105337 62002 105717
rect 62382 105337 62394 105717
rect 62774 105337 62786 105717
rect 63166 105337 63178 105717
rect 63558 105337 63600 105717
rect 60000 105325 63600 105337
rect 60000 104945 60042 105325
rect 60422 104945 60434 105325
rect 60814 104945 60826 105325
rect 61206 104945 61218 105325
rect 61598 104945 61610 105325
rect 61990 104945 62002 105325
rect 62382 104945 62394 105325
rect 62774 104945 62786 105325
rect 63166 104945 63178 105325
rect 63558 104945 63600 105325
rect 60000 104933 63600 104945
rect 60000 104553 60042 104933
rect 60422 104553 60434 104933
rect 60814 104553 60826 104933
rect 61206 104553 61218 104933
rect 61598 104553 61610 104933
rect 61990 104553 62002 104933
rect 62382 104553 62394 104933
rect 62774 104553 62786 104933
rect 63166 104553 63178 104933
rect 63558 104553 63600 104933
rect 60000 104541 63600 104553
rect 60000 104161 60042 104541
rect 60422 104161 60434 104541
rect 60814 104161 60826 104541
rect 61206 104161 61218 104541
rect 61598 104161 61610 104541
rect 61990 104161 62002 104541
rect 62382 104161 62394 104541
rect 62774 104161 62786 104541
rect 63166 104161 63178 104541
rect 63558 104161 63600 104541
rect 60000 103998 63600 104161
rect 68316 106501 69316 120161
rect 68316 106121 68430 106501
rect 68810 106121 68822 106501
rect 69202 106121 69316 106501
rect 68316 106109 69316 106121
rect 68316 105729 68430 106109
rect 68810 105729 68822 106109
rect 69202 105729 69316 106109
rect 68316 105717 69316 105729
rect 68316 105337 68430 105717
rect 68810 105337 68822 105717
rect 69202 105337 69316 105717
rect 68316 105325 69316 105337
rect 68316 104945 68430 105325
rect 68810 104945 68822 105325
rect 69202 104945 69316 105325
rect 68316 104933 69316 104945
rect 68316 104553 68430 104933
rect 68810 104553 68822 104933
rect 69202 104553 69316 104933
rect 68316 104541 69316 104553
rect 68316 104161 68430 104541
rect 68810 104161 68822 104541
rect 69202 104161 69316 104541
rect 56000 101169 59600 101332
rect 56000 100789 56042 101169
rect 56422 100789 56434 101169
rect 56814 100789 56826 101169
rect 57206 100789 57218 101169
rect 57598 100789 57610 101169
rect 57990 100789 58002 101169
rect 58382 100789 58394 101169
rect 58774 100789 58786 101169
rect 59166 100789 59178 101169
rect 59558 100789 59600 101169
rect 56000 100777 59600 100789
rect 56000 100397 56042 100777
rect 56422 100397 56434 100777
rect 56814 100397 56826 100777
rect 57206 100397 57218 100777
rect 57598 100397 57610 100777
rect 57990 100397 58002 100777
rect 58382 100397 58394 100777
rect 58774 100397 58786 100777
rect 59166 100397 59178 100777
rect 59558 100397 59600 100777
rect 56000 100385 59600 100397
rect 56000 100005 56042 100385
rect 56422 100005 56434 100385
rect 56814 100005 56826 100385
rect 57206 100005 57218 100385
rect 57598 100005 57610 100385
rect 57990 100005 58002 100385
rect 58382 100005 58394 100385
rect 58774 100005 58786 100385
rect 59166 100005 59178 100385
rect 59558 100005 59600 100385
rect 56000 99993 59600 100005
rect 56000 99613 56042 99993
rect 56422 99613 56434 99993
rect 56814 99613 56826 99993
rect 57206 99613 57218 99993
rect 57598 99613 57610 99993
rect 57990 99613 58002 99993
rect 58382 99613 58394 99993
rect 58774 99613 58786 99993
rect 59166 99613 59178 99993
rect 59558 99613 59600 99993
rect 56000 99601 59600 99613
rect 56000 99221 56042 99601
rect 56422 99221 56434 99601
rect 56814 99221 56826 99601
rect 57206 99221 57218 99601
rect 57598 99221 57610 99601
rect 57990 99221 58002 99601
rect 58382 99221 58394 99601
rect 58774 99221 58786 99601
rect 59166 99221 59178 99601
rect 59558 99221 59600 99601
rect 56000 99209 59600 99221
rect 56000 98829 56042 99209
rect 56422 98829 56434 99209
rect 56814 98829 56826 99209
rect 57206 98829 57218 99209
rect 57598 98829 57610 99209
rect 57990 98829 58002 99209
rect 58382 98829 58394 99209
rect 58774 98829 58786 99209
rect 59166 98829 59178 99209
rect 59558 98829 59600 99209
rect 56000 98666 59600 98829
rect 60000 90501 63600 90664
rect 60000 90121 60042 90501
rect 60422 90121 60434 90501
rect 60814 90121 60826 90501
rect 61206 90121 61218 90501
rect 61598 90121 61610 90501
rect 61990 90121 62002 90501
rect 62382 90121 62394 90501
rect 62774 90121 62786 90501
rect 63166 90121 63178 90501
rect 63558 90121 63600 90501
rect 60000 90109 63600 90121
rect 60000 89729 60042 90109
rect 60422 89729 60434 90109
rect 60814 89729 60826 90109
rect 61206 89729 61218 90109
rect 61598 89729 61610 90109
rect 61990 89729 62002 90109
rect 62382 89729 62394 90109
rect 62774 89729 62786 90109
rect 63166 89729 63178 90109
rect 63558 89729 63600 90109
rect 60000 89717 63600 89729
rect 60000 89337 60042 89717
rect 60422 89337 60434 89717
rect 60814 89337 60826 89717
rect 61206 89337 61218 89717
rect 61598 89337 61610 89717
rect 61990 89337 62002 89717
rect 62382 89337 62394 89717
rect 62774 89337 62786 89717
rect 63166 89337 63178 89717
rect 63558 89337 63600 89717
rect 60000 89325 63600 89337
rect 60000 88945 60042 89325
rect 60422 88945 60434 89325
rect 60814 88945 60826 89325
rect 61206 88945 61218 89325
rect 61598 88945 61610 89325
rect 61990 88945 62002 89325
rect 62382 88945 62394 89325
rect 62774 88945 62786 89325
rect 63166 88945 63178 89325
rect 63558 88945 63600 89325
rect 60000 88933 63600 88945
rect 60000 88553 60042 88933
rect 60422 88553 60434 88933
rect 60814 88553 60826 88933
rect 61206 88553 61218 88933
rect 61598 88553 61610 88933
rect 61990 88553 62002 88933
rect 62382 88553 62394 88933
rect 62774 88553 62786 88933
rect 63166 88553 63178 88933
rect 63558 88553 63600 88933
rect 60000 88541 63600 88553
rect 60000 88161 60042 88541
rect 60422 88161 60434 88541
rect 60814 88161 60826 88541
rect 61206 88161 61218 88541
rect 61598 88161 61610 88541
rect 61990 88161 62002 88541
rect 62382 88161 62394 88541
rect 62774 88161 62786 88541
rect 63166 88161 63178 88541
rect 63558 88161 63600 88541
rect 60000 87998 63600 88161
rect 68316 90501 69316 104161
rect 68316 90121 68430 90501
rect 68810 90121 68822 90501
rect 69202 90121 69316 90501
rect 68316 90109 69316 90121
rect 68316 89729 68430 90109
rect 68810 89729 68822 90109
rect 69202 89729 69316 90109
rect 68316 89717 69316 89729
rect 68316 89337 68430 89717
rect 68810 89337 68822 89717
rect 69202 89337 69316 89717
rect 68316 89325 69316 89337
rect 68316 88945 68430 89325
rect 68810 88945 68822 89325
rect 69202 88945 69316 89325
rect 68316 88933 69316 88945
rect 68316 88553 68430 88933
rect 68810 88553 68822 88933
rect 69202 88553 69316 88933
rect 68316 88541 69316 88553
rect 68316 88161 68430 88541
rect 68810 88161 68822 88541
rect 69202 88161 69316 88541
rect 56000 85169 59600 85332
rect 56000 84789 56042 85169
rect 56422 84789 56434 85169
rect 56814 84789 56826 85169
rect 57206 84789 57218 85169
rect 57598 84789 57610 85169
rect 57990 84789 58002 85169
rect 58382 84789 58394 85169
rect 58774 84789 58786 85169
rect 59166 84789 59178 85169
rect 59558 84789 59600 85169
rect 56000 84777 59600 84789
rect 56000 84397 56042 84777
rect 56422 84397 56434 84777
rect 56814 84397 56826 84777
rect 57206 84397 57218 84777
rect 57598 84397 57610 84777
rect 57990 84397 58002 84777
rect 58382 84397 58394 84777
rect 58774 84397 58786 84777
rect 59166 84397 59178 84777
rect 59558 84397 59600 84777
rect 56000 84385 59600 84397
rect 56000 84005 56042 84385
rect 56422 84005 56434 84385
rect 56814 84005 56826 84385
rect 57206 84005 57218 84385
rect 57598 84005 57610 84385
rect 57990 84005 58002 84385
rect 58382 84005 58394 84385
rect 58774 84005 58786 84385
rect 59166 84005 59178 84385
rect 59558 84005 59600 84385
rect 56000 83993 59600 84005
rect 56000 83613 56042 83993
rect 56422 83613 56434 83993
rect 56814 83613 56826 83993
rect 57206 83613 57218 83993
rect 57598 83613 57610 83993
rect 57990 83613 58002 83993
rect 58382 83613 58394 83993
rect 58774 83613 58786 83993
rect 59166 83613 59178 83993
rect 59558 83613 59600 83993
rect 56000 83601 59600 83613
rect 56000 83221 56042 83601
rect 56422 83221 56434 83601
rect 56814 83221 56826 83601
rect 57206 83221 57218 83601
rect 57598 83221 57610 83601
rect 57990 83221 58002 83601
rect 58382 83221 58394 83601
rect 58774 83221 58786 83601
rect 59166 83221 59178 83601
rect 59558 83221 59600 83601
rect 56000 83209 59600 83221
rect 56000 82829 56042 83209
rect 56422 82829 56434 83209
rect 56814 82829 56826 83209
rect 57206 82829 57218 83209
rect 57598 82829 57610 83209
rect 57990 82829 58002 83209
rect 58382 82829 58394 83209
rect 58774 82829 58786 83209
rect 59166 82829 59178 83209
rect 59558 82829 59600 83209
rect 56000 82666 59600 82829
rect 68316 75970 69316 88161
rect 68316 75590 68430 75970
rect 68810 75590 68822 75970
rect 69202 75590 69316 75970
rect 60000 74501 63600 74664
rect 60000 74121 60042 74501
rect 60422 74121 60434 74501
rect 60814 74121 60826 74501
rect 61206 74121 61218 74501
rect 61598 74121 61610 74501
rect 61990 74121 62002 74501
rect 62382 74121 62394 74501
rect 62774 74121 62786 74501
rect 63166 74121 63178 74501
rect 63558 74121 63600 74501
rect 60000 74109 63600 74121
rect 60000 73729 60042 74109
rect 60422 73729 60434 74109
rect 60814 73729 60826 74109
rect 61206 73729 61218 74109
rect 61598 73729 61610 74109
rect 61990 73729 62002 74109
rect 62382 73729 62394 74109
rect 62774 73729 62786 74109
rect 63166 73729 63178 74109
rect 63558 73729 63600 74109
rect 60000 73717 63600 73729
rect 60000 73337 60042 73717
rect 60422 73337 60434 73717
rect 60814 73337 60826 73717
rect 61206 73337 61218 73717
rect 61598 73337 61610 73717
rect 61990 73337 62002 73717
rect 62382 73337 62394 73717
rect 62774 73337 62786 73717
rect 63166 73337 63178 73717
rect 63558 73337 63600 73717
rect 60000 73325 63600 73337
rect 60000 72945 60042 73325
rect 60422 72945 60434 73325
rect 60814 72945 60826 73325
rect 61206 72945 61218 73325
rect 61598 72945 61610 73325
rect 61990 72945 62002 73325
rect 62382 72945 62394 73325
rect 62774 72945 62786 73325
rect 63166 72945 63178 73325
rect 63558 72945 63600 73325
rect 60000 72933 63600 72945
rect 60000 72553 60042 72933
rect 60422 72553 60434 72933
rect 60814 72553 60826 72933
rect 61206 72553 61218 72933
rect 61598 72553 61610 72933
rect 61990 72553 62002 72933
rect 62382 72553 62394 72933
rect 62774 72553 62786 72933
rect 63166 72553 63178 72933
rect 63558 72553 63600 72933
rect 60000 72541 63600 72553
rect 60000 72161 60042 72541
rect 60422 72161 60434 72541
rect 60814 72161 60826 72541
rect 61206 72161 61218 72541
rect 61598 72161 61610 72541
rect 61990 72161 62002 72541
rect 62382 72161 62394 72541
rect 62774 72161 62786 72541
rect 63166 72161 63178 72541
rect 63558 72161 63600 72541
rect 60000 71998 63600 72161
rect 68316 74501 69316 75590
rect 68316 74121 68430 74501
rect 68810 74121 68822 74501
rect 69202 74121 69316 74501
rect 68316 74109 69316 74121
rect 68316 73729 68430 74109
rect 68810 73729 68822 74109
rect 69202 73729 69316 74109
rect 68316 73717 69316 73729
rect 68316 73337 68430 73717
rect 68810 73337 68822 73717
rect 69202 73337 69316 73717
rect 68316 73325 69316 73337
rect 68316 72945 68430 73325
rect 68810 72945 68822 73325
rect 69202 72945 69316 73325
rect 68316 72933 69316 72945
rect 68316 72553 68430 72933
rect 68810 72553 68822 72933
rect 69202 72553 69316 72933
rect 68316 72541 69316 72553
rect 68316 72161 68430 72541
rect 68810 72161 68822 72541
rect 69202 72161 69316 72541
rect 68316 69406 69316 72161
rect 69716 153742 70716 153856
rect 69716 153362 69830 153742
rect 70210 153362 70222 153742
rect 70602 153362 70716 153742
rect 69716 153350 70716 153362
rect 69716 152970 69830 153350
rect 70210 152970 70222 153350
rect 70602 152970 70716 153350
rect 69716 149169 70716 152970
rect 69716 148789 69830 149169
rect 70210 148789 70222 149169
rect 70602 148789 70716 149169
rect 69716 148777 70716 148789
rect 69716 148397 69830 148777
rect 70210 148397 70222 148777
rect 70602 148397 70716 148777
rect 69716 148385 70716 148397
rect 69716 148005 69830 148385
rect 70210 148005 70222 148385
rect 70602 148005 70716 148385
rect 69716 147993 70716 148005
rect 69716 147613 69830 147993
rect 70210 147613 70222 147993
rect 70602 147613 70716 147993
rect 69716 147601 70716 147613
rect 69716 147221 69830 147601
rect 70210 147221 70222 147601
rect 70602 147221 70716 147601
rect 69716 147209 70716 147221
rect 69716 146829 69830 147209
rect 70210 146829 70222 147209
rect 70602 146829 70716 147209
rect 69716 135210 70716 146829
rect 69716 134830 69830 135210
rect 70210 134830 70222 135210
rect 70602 134830 70716 135210
rect 69716 133169 70716 134830
rect 69716 132789 69830 133169
rect 70210 132789 70222 133169
rect 70602 132789 70716 133169
rect 69716 132777 70716 132789
rect 69716 132397 69830 132777
rect 70210 132397 70222 132777
rect 70602 132397 70716 132777
rect 69716 132385 70716 132397
rect 69716 132005 69830 132385
rect 70210 132005 70222 132385
rect 70602 132005 70716 132385
rect 69716 131993 70716 132005
rect 69716 131613 69830 131993
rect 70210 131613 70222 131993
rect 70602 131613 70716 131993
rect 69716 131601 70716 131613
rect 69716 131221 69830 131601
rect 70210 131221 70222 131601
rect 70602 131221 70716 131601
rect 69716 131209 70716 131221
rect 69716 130829 69830 131209
rect 70210 130829 70222 131209
rect 70602 130829 70716 131209
rect 69716 120090 70716 130829
rect 69716 119710 69830 120090
rect 70210 119710 70222 120090
rect 70602 119710 70716 120090
rect 69716 117169 70716 119710
rect 69716 116789 69830 117169
rect 70210 116789 70222 117169
rect 70602 116789 70716 117169
rect 69716 116777 70716 116789
rect 69716 116397 69830 116777
rect 70210 116397 70222 116777
rect 70602 116397 70716 116777
rect 69716 116385 70716 116397
rect 69716 116005 69830 116385
rect 70210 116005 70222 116385
rect 70602 116005 70716 116385
rect 69716 115993 70716 116005
rect 69716 115613 69830 115993
rect 70210 115613 70222 115993
rect 70602 115613 70716 115993
rect 69716 115601 70716 115613
rect 69716 115221 69830 115601
rect 70210 115221 70222 115601
rect 70602 115221 70716 115601
rect 69716 115209 70716 115221
rect 69716 114829 69830 115209
rect 70210 114829 70222 115209
rect 70602 114829 70716 115209
rect 69716 104970 70716 114829
rect 69716 104590 69830 104970
rect 70210 104590 70222 104970
rect 70602 104590 70716 104970
rect 69716 101169 70716 104590
rect 69716 100789 69830 101169
rect 70210 100789 70222 101169
rect 70602 100789 70716 101169
rect 69716 100777 70716 100789
rect 69716 100397 69830 100777
rect 70210 100397 70222 100777
rect 70602 100397 70716 100777
rect 69716 100385 70716 100397
rect 69716 100005 69830 100385
rect 70210 100005 70222 100385
rect 70602 100005 70716 100385
rect 69716 99993 70716 100005
rect 69716 99613 69830 99993
rect 70210 99613 70222 99993
rect 70602 99613 70716 99993
rect 69716 99601 70716 99613
rect 69716 99221 69830 99601
rect 70210 99221 70222 99601
rect 70602 99221 70716 99601
rect 69716 99209 70716 99221
rect 69716 98829 69830 99209
rect 70210 98829 70222 99209
rect 70602 98829 70716 99209
rect 69716 89850 70716 98829
rect 69716 89470 69830 89850
rect 70210 89470 70222 89850
rect 70602 89470 70716 89850
rect 69716 85169 70716 89470
rect 69716 84789 69830 85169
rect 70210 84789 70222 85169
rect 70602 84789 70716 85169
rect 69716 84777 70716 84789
rect 69716 84397 69830 84777
rect 70210 84397 70222 84777
rect 70602 84397 70716 84777
rect 69716 84385 70716 84397
rect 69716 84005 69830 84385
rect 70210 84005 70222 84385
rect 70602 84005 70716 84385
rect 69716 83993 70716 84005
rect 69716 83613 69830 83993
rect 70210 83613 70222 83993
rect 70602 83613 70716 83993
rect 69716 83601 70716 83613
rect 69716 83221 69830 83601
rect 70210 83221 70222 83601
rect 70602 83221 70716 83601
rect 69716 83209 70716 83221
rect 69716 82829 69830 83209
rect 70210 82829 70222 83209
rect 70602 82829 70716 83209
rect 69716 74730 70716 82829
rect 69716 74350 69830 74730
rect 70210 74350 70222 74730
rect 70602 74350 70716 74730
rect 69716 70806 70716 74350
rect 69716 70426 69830 70806
rect 70210 70426 70222 70806
rect 70602 70426 70716 70806
rect 69716 70414 70716 70426
rect 69716 70034 69830 70414
rect 70210 70034 70222 70414
rect 70602 70034 70716 70414
rect 69716 69920 70716 70034
rect 74116 153742 74556 155256
rect 74116 153362 74146 153742
rect 74526 153362 74556 153742
rect 74116 153350 74556 153362
rect 74116 152970 74146 153350
rect 74526 152970 74556 153350
rect 74116 151243 74556 152970
rect 74116 151157 74209 151243
rect 74295 151157 74377 151243
rect 74463 151157 74556 151243
rect 74116 150330 74556 151157
rect 74116 149950 74146 150330
rect 74526 149950 74556 150330
rect 74116 149731 74556 149950
rect 74116 149645 74209 149731
rect 74295 149645 74377 149731
rect 74463 149645 74556 149731
rect 74116 148219 74556 149645
rect 74116 148133 74209 148219
rect 74295 148133 74377 148219
rect 74463 148133 74556 148219
rect 74116 146707 74556 148133
rect 74116 146621 74209 146707
rect 74295 146621 74377 146707
rect 74463 146621 74556 146707
rect 74116 145195 74556 146621
rect 74116 145109 74209 145195
rect 74295 145109 74377 145195
rect 74463 145109 74556 145195
rect 74116 143683 74556 145109
rect 74116 143597 74209 143683
rect 74295 143597 74377 143683
rect 74463 143597 74556 143683
rect 74116 142171 74556 143597
rect 74116 142085 74209 142171
rect 74295 142085 74377 142171
rect 74463 142085 74556 142171
rect 74116 140659 74556 142085
rect 74116 140573 74209 140659
rect 74295 140573 74377 140659
rect 74463 140573 74556 140659
rect 74116 139147 74556 140573
rect 74116 139061 74209 139147
rect 74295 139061 74377 139147
rect 74463 139061 74556 139147
rect 74116 137635 74556 139061
rect 74116 137549 74209 137635
rect 74295 137549 74377 137635
rect 74463 137549 74556 137635
rect 74116 136123 74556 137549
rect 74116 136037 74209 136123
rect 74295 136037 74377 136123
rect 74463 136037 74556 136123
rect 74116 135210 74556 136037
rect 74116 134830 74146 135210
rect 74526 134830 74556 135210
rect 74116 134611 74556 134830
rect 74116 134525 74209 134611
rect 74295 134525 74377 134611
rect 74463 134525 74556 134611
rect 74116 133099 74556 134525
rect 74116 133013 74209 133099
rect 74295 133013 74377 133099
rect 74463 133013 74556 133099
rect 74116 131587 74556 133013
rect 74116 131501 74209 131587
rect 74295 131501 74377 131587
rect 74463 131501 74556 131587
rect 74116 130075 74556 131501
rect 74116 129989 74209 130075
rect 74295 129989 74377 130075
rect 74463 129989 74556 130075
rect 74116 128563 74556 129989
rect 74116 128477 74209 128563
rect 74295 128477 74377 128563
rect 74463 128477 74556 128563
rect 74116 127051 74556 128477
rect 74116 126965 74209 127051
rect 74295 126965 74377 127051
rect 74463 126965 74556 127051
rect 74116 125539 74556 126965
rect 74116 125453 74209 125539
rect 74295 125453 74377 125539
rect 74463 125453 74556 125539
rect 74116 124027 74556 125453
rect 74116 123941 74209 124027
rect 74295 123941 74377 124027
rect 74463 123941 74556 124027
rect 74116 122515 74556 123941
rect 74116 122429 74209 122515
rect 74295 122429 74377 122515
rect 74463 122429 74556 122515
rect 74116 121003 74556 122429
rect 74116 120917 74209 121003
rect 74295 120917 74377 121003
rect 74463 120917 74556 121003
rect 74116 120090 74556 120917
rect 74116 119710 74146 120090
rect 74526 119710 74556 120090
rect 74116 119491 74556 119710
rect 74116 119405 74209 119491
rect 74295 119405 74377 119491
rect 74463 119405 74556 119491
rect 74116 117979 74556 119405
rect 74116 117893 74209 117979
rect 74295 117893 74377 117979
rect 74463 117893 74556 117979
rect 74116 116467 74556 117893
rect 74116 116381 74209 116467
rect 74295 116381 74377 116467
rect 74463 116381 74556 116467
rect 74116 114955 74556 116381
rect 74116 114869 74209 114955
rect 74295 114869 74377 114955
rect 74463 114869 74556 114955
rect 74116 113443 74556 114869
rect 74116 113357 74209 113443
rect 74295 113357 74377 113443
rect 74463 113357 74556 113443
rect 74116 111931 74556 113357
rect 74116 111845 74209 111931
rect 74295 111845 74377 111931
rect 74463 111845 74556 111931
rect 74116 110419 74556 111845
rect 74116 110333 74209 110419
rect 74295 110333 74377 110419
rect 74463 110333 74556 110419
rect 74116 108907 74556 110333
rect 74116 108821 74209 108907
rect 74295 108821 74377 108907
rect 74463 108821 74556 108907
rect 74116 107395 74556 108821
rect 74116 107309 74209 107395
rect 74295 107309 74377 107395
rect 74463 107309 74556 107395
rect 74116 105883 74556 107309
rect 74116 105797 74209 105883
rect 74295 105797 74377 105883
rect 74463 105797 74556 105883
rect 74116 104970 74556 105797
rect 74116 104590 74146 104970
rect 74526 104590 74556 104970
rect 74116 104371 74556 104590
rect 74116 104285 74209 104371
rect 74295 104285 74377 104371
rect 74463 104285 74556 104371
rect 74116 102859 74556 104285
rect 74116 102773 74209 102859
rect 74295 102773 74377 102859
rect 74463 102773 74556 102859
rect 74116 101347 74556 102773
rect 74116 101261 74209 101347
rect 74295 101261 74377 101347
rect 74463 101261 74556 101347
rect 74116 99835 74556 101261
rect 74116 99749 74209 99835
rect 74295 99749 74377 99835
rect 74463 99749 74556 99835
rect 74116 98323 74556 99749
rect 74116 98237 74209 98323
rect 74295 98237 74377 98323
rect 74463 98237 74556 98323
rect 74116 96811 74556 98237
rect 74116 96725 74209 96811
rect 74295 96725 74377 96811
rect 74463 96725 74556 96811
rect 74116 95299 74556 96725
rect 74116 95213 74209 95299
rect 74295 95213 74377 95299
rect 74463 95213 74556 95299
rect 74116 93787 74556 95213
rect 74116 93701 74209 93787
rect 74295 93701 74377 93787
rect 74463 93701 74556 93787
rect 74116 92275 74556 93701
rect 74116 92189 74209 92275
rect 74295 92189 74377 92275
rect 74463 92189 74556 92275
rect 74116 90763 74556 92189
rect 74116 90677 74209 90763
rect 74295 90677 74377 90763
rect 74463 90677 74556 90763
rect 74116 89850 74556 90677
rect 74116 89470 74146 89850
rect 74526 89470 74556 89850
rect 74116 89251 74556 89470
rect 74116 89165 74209 89251
rect 74295 89165 74377 89251
rect 74463 89165 74556 89251
rect 74116 87739 74556 89165
rect 74116 87653 74209 87739
rect 74295 87653 74377 87739
rect 74463 87653 74556 87739
rect 74116 86227 74556 87653
rect 74116 86141 74209 86227
rect 74295 86141 74377 86227
rect 74463 86141 74556 86227
rect 74116 84715 74556 86141
rect 74116 84629 74209 84715
rect 74295 84629 74377 84715
rect 74463 84629 74556 84715
rect 74116 83203 74556 84629
rect 74116 83117 74209 83203
rect 74295 83117 74377 83203
rect 74463 83117 74556 83203
rect 74116 81691 74556 83117
rect 74116 81605 74209 81691
rect 74295 81605 74377 81691
rect 74463 81605 74556 81691
rect 74116 80179 74556 81605
rect 74116 80093 74209 80179
rect 74295 80093 74377 80179
rect 74463 80093 74556 80179
rect 74116 78667 74556 80093
rect 74116 78581 74209 78667
rect 74295 78581 74377 78667
rect 74463 78581 74556 78667
rect 74116 77155 74556 78581
rect 74116 77069 74209 77155
rect 74295 77069 74377 77155
rect 74463 77069 74556 77155
rect 74116 75643 74556 77069
rect 74116 75557 74209 75643
rect 74295 75557 74377 75643
rect 74463 75557 74556 75643
rect 74116 74730 74556 75557
rect 74116 74350 74146 74730
rect 74526 74350 74556 74730
rect 74116 74131 74556 74350
rect 74116 74045 74209 74131
rect 74295 74045 74377 74131
rect 74463 74045 74556 74131
rect 74116 72619 74556 74045
rect 74116 72533 74209 72619
rect 74295 72533 74377 72619
rect 74463 72533 74556 72619
rect 74116 70806 74556 72533
rect 74116 70426 74146 70806
rect 74526 70426 74556 70806
rect 74116 70414 74556 70426
rect 74116 70034 74146 70414
rect 74526 70034 74556 70414
rect 68316 69026 68430 69406
rect 68810 69026 68822 69406
rect 69202 69026 69316 69406
rect 68316 69014 69316 69026
rect 68316 68634 68430 69014
rect 68810 68634 68822 69014
rect 69202 68634 69316 69014
rect 68316 68520 69316 68634
rect 74116 68520 74556 70034
rect 75356 155142 75796 155256
rect 75356 154762 75386 155142
rect 75766 154762 75796 155142
rect 75356 154750 75796 154762
rect 75356 154370 75386 154750
rect 75766 154370 75796 154750
rect 75356 151999 75796 154370
rect 75356 151913 75449 151999
rect 75535 151913 75617 151999
rect 75703 151913 75796 151999
rect 75356 151570 75796 151913
rect 75356 151190 75386 151570
rect 75766 151190 75796 151570
rect 75356 150487 75796 151190
rect 75356 150401 75449 150487
rect 75535 150401 75617 150487
rect 75703 150401 75796 150487
rect 75356 148975 75796 150401
rect 75356 148889 75449 148975
rect 75535 148889 75617 148975
rect 75703 148889 75796 148975
rect 75356 147463 75796 148889
rect 75356 147377 75449 147463
rect 75535 147377 75617 147463
rect 75703 147377 75796 147463
rect 75356 145951 75796 147377
rect 75356 145865 75449 145951
rect 75535 145865 75617 145951
rect 75703 145865 75796 145951
rect 75356 144439 75796 145865
rect 75356 144353 75449 144439
rect 75535 144353 75617 144439
rect 75703 144353 75796 144439
rect 75356 142927 75796 144353
rect 75356 142841 75449 142927
rect 75535 142841 75617 142927
rect 75703 142841 75796 142927
rect 75356 141415 75796 142841
rect 75356 141329 75449 141415
rect 75535 141329 75617 141415
rect 75703 141329 75796 141415
rect 75356 139903 75796 141329
rect 75356 139817 75449 139903
rect 75535 139817 75617 139903
rect 75703 139817 75796 139903
rect 75356 138391 75796 139817
rect 75356 138305 75449 138391
rect 75535 138305 75617 138391
rect 75703 138305 75796 138391
rect 75356 136879 75796 138305
rect 75356 136793 75449 136879
rect 75535 136793 75617 136879
rect 75703 136793 75796 136879
rect 75356 136450 75796 136793
rect 75356 136070 75386 136450
rect 75766 136070 75796 136450
rect 75356 135367 75796 136070
rect 75356 135281 75449 135367
rect 75535 135281 75617 135367
rect 75703 135281 75796 135367
rect 75356 133855 75796 135281
rect 75356 133769 75449 133855
rect 75535 133769 75617 133855
rect 75703 133769 75796 133855
rect 75356 132343 75796 133769
rect 75356 132257 75449 132343
rect 75535 132257 75617 132343
rect 75703 132257 75796 132343
rect 75356 130831 75796 132257
rect 75356 130745 75449 130831
rect 75535 130745 75617 130831
rect 75703 130745 75796 130831
rect 75356 129319 75796 130745
rect 75356 129233 75449 129319
rect 75535 129233 75617 129319
rect 75703 129233 75796 129319
rect 75356 127807 75796 129233
rect 75356 127721 75449 127807
rect 75535 127721 75617 127807
rect 75703 127721 75796 127807
rect 75356 126295 75796 127721
rect 75356 126209 75449 126295
rect 75535 126209 75617 126295
rect 75703 126209 75796 126295
rect 75356 124783 75796 126209
rect 75356 124697 75449 124783
rect 75535 124697 75617 124783
rect 75703 124697 75796 124783
rect 75356 123271 75796 124697
rect 75356 123185 75449 123271
rect 75535 123185 75617 123271
rect 75703 123185 75796 123271
rect 75356 121759 75796 123185
rect 75356 121673 75449 121759
rect 75535 121673 75617 121759
rect 75703 121673 75796 121759
rect 75356 121330 75796 121673
rect 75356 120950 75386 121330
rect 75766 120950 75796 121330
rect 75356 120247 75796 120950
rect 75356 120161 75449 120247
rect 75535 120161 75617 120247
rect 75703 120161 75796 120247
rect 75356 118735 75796 120161
rect 75356 118649 75449 118735
rect 75535 118649 75617 118735
rect 75703 118649 75796 118735
rect 75356 117223 75796 118649
rect 75356 117137 75449 117223
rect 75535 117137 75617 117223
rect 75703 117137 75796 117223
rect 75356 115711 75796 117137
rect 75356 115625 75449 115711
rect 75535 115625 75617 115711
rect 75703 115625 75796 115711
rect 75356 114199 75796 115625
rect 75356 114113 75449 114199
rect 75535 114113 75617 114199
rect 75703 114113 75796 114199
rect 75356 112687 75796 114113
rect 75356 112601 75449 112687
rect 75535 112601 75617 112687
rect 75703 112601 75796 112687
rect 75356 111175 75796 112601
rect 75356 111089 75449 111175
rect 75535 111089 75617 111175
rect 75703 111089 75796 111175
rect 75356 109663 75796 111089
rect 75356 109577 75449 109663
rect 75535 109577 75617 109663
rect 75703 109577 75796 109663
rect 75356 108151 75796 109577
rect 75356 108065 75449 108151
rect 75535 108065 75617 108151
rect 75703 108065 75796 108151
rect 75356 106639 75796 108065
rect 75356 106553 75449 106639
rect 75535 106553 75617 106639
rect 75703 106553 75796 106639
rect 75356 106210 75796 106553
rect 75356 105830 75386 106210
rect 75766 105830 75796 106210
rect 75356 105127 75796 105830
rect 75356 105041 75449 105127
rect 75535 105041 75617 105127
rect 75703 105041 75796 105127
rect 75356 103615 75796 105041
rect 75356 103529 75449 103615
rect 75535 103529 75617 103615
rect 75703 103529 75796 103615
rect 75356 102103 75796 103529
rect 75356 102017 75449 102103
rect 75535 102017 75617 102103
rect 75703 102017 75796 102103
rect 75356 100591 75796 102017
rect 75356 100505 75449 100591
rect 75535 100505 75617 100591
rect 75703 100505 75796 100591
rect 75356 99079 75796 100505
rect 75356 98993 75449 99079
rect 75535 98993 75617 99079
rect 75703 98993 75796 99079
rect 75356 97567 75796 98993
rect 75356 97481 75449 97567
rect 75535 97481 75617 97567
rect 75703 97481 75796 97567
rect 75356 96055 75796 97481
rect 75356 95969 75449 96055
rect 75535 95969 75617 96055
rect 75703 95969 75796 96055
rect 75356 94543 75796 95969
rect 75356 94457 75449 94543
rect 75535 94457 75617 94543
rect 75703 94457 75796 94543
rect 75356 93031 75796 94457
rect 75356 92945 75449 93031
rect 75535 92945 75617 93031
rect 75703 92945 75796 93031
rect 75356 91519 75796 92945
rect 75356 91433 75449 91519
rect 75535 91433 75617 91519
rect 75703 91433 75796 91519
rect 75356 91090 75796 91433
rect 75356 90710 75386 91090
rect 75766 90710 75796 91090
rect 75356 90007 75796 90710
rect 75356 89921 75449 90007
rect 75535 89921 75617 90007
rect 75703 89921 75796 90007
rect 75356 88495 75796 89921
rect 75356 88409 75449 88495
rect 75535 88409 75617 88495
rect 75703 88409 75796 88495
rect 75356 86983 75796 88409
rect 75356 86897 75449 86983
rect 75535 86897 75617 86983
rect 75703 86897 75796 86983
rect 75356 85471 75796 86897
rect 75356 85385 75449 85471
rect 75535 85385 75617 85471
rect 75703 85385 75796 85471
rect 75356 83959 75796 85385
rect 75356 83873 75449 83959
rect 75535 83873 75617 83959
rect 75703 83873 75796 83959
rect 75356 82447 75796 83873
rect 75356 82361 75449 82447
rect 75535 82361 75617 82447
rect 75703 82361 75796 82447
rect 75356 80935 75796 82361
rect 75356 80849 75449 80935
rect 75535 80849 75617 80935
rect 75703 80849 75796 80935
rect 75356 79423 75796 80849
rect 75356 79337 75449 79423
rect 75535 79337 75617 79423
rect 75703 79337 75796 79423
rect 75356 77911 75796 79337
rect 75356 77825 75449 77911
rect 75535 77825 75617 77911
rect 75703 77825 75796 77911
rect 75356 76399 75796 77825
rect 75356 76313 75449 76399
rect 75535 76313 75617 76399
rect 75703 76313 75796 76399
rect 75356 75970 75796 76313
rect 75356 75590 75386 75970
rect 75766 75590 75796 75970
rect 75356 74887 75796 75590
rect 75356 74801 75449 74887
rect 75535 74801 75617 74887
rect 75703 74801 75796 74887
rect 75356 73375 75796 74801
rect 75356 73289 75449 73375
rect 75535 73289 75617 73375
rect 75703 73289 75796 73375
rect 75356 71863 75796 73289
rect 75356 71777 75449 71863
rect 75535 71777 75617 71863
rect 75703 71777 75796 71863
rect 75356 69406 75796 71777
rect 75356 69026 75386 69406
rect 75766 69026 75796 69406
rect 75356 69014 75796 69026
rect 75356 68634 75386 69014
rect 75766 68634 75796 69014
rect 75356 68520 75796 68634
rect 89236 153742 89676 155256
rect 89236 153362 89266 153742
rect 89646 153362 89676 153742
rect 89236 153350 89676 153362
rect 89236 152970 89266 153350
rect 89646 152970 89676 153350
rect 89236 151243 89676 152970
rect 89236 151157 89329 151243
rect 89415 151157 89497 151243
rect 89583 151157 89676 151243
rect 89236 150330 89676 151157
rect 89236 149950 89266 150330
rect 89646 149950 89676 150330
rect 89236 149731 89676 149950
rect 89236 149645 89329 149731
rect 89415 149645 89497 149731
rect 89583 149645 89676 149731
rect 89236 148219 89676 149645
rect 89236 148133 89329 148219
rect 89415 148133 89497 148219
rect 89583 148133 89676 148219
rect 89236 146707 89676 148133
rect 89236 146621 89329 146707
rect 89415 146621 89497 146707
rect 89583 146621 89676 146707
rect 89236 145195 89676 146621
rect 89236 145109 89329 145195
rect 89415 145109 89497 145195
rect 89583 145109 89676 145195
rect 89236 143683 89676 145109
rect 89236 143597 89329 143683
rect 89415 143597 89497 143683
rect 89583 143597 89676 143683
rect 89236 142171 89676 143597
rect 89236 142085 89329 142171
rect 89415 142085 89497 142171
rect 89583 142085 89676 142171
rect 89236 140659 89676 142085
rect 89236 140573 89329 140659
rect 89415 140573 89497 140659
rect 89583 140573 89676 140659
rect 89236 139147 89676 140573
rect 89236 139061 89329 139147
rect 89415 139061 89497 139147
rect 89583 139061 89676 139147
rect 89236 137635 89676 139061
rect 89236 137549 89329 137635
rect 89415 137549 89497 137635
rect 89583 137549 89676 137635
rect 89236 136123 89676 137549
rect 89236 136037 89329 136123
rect 89415 136037 89497 136123
rect 89583 136037 89676 136123
rect 89236 135210 89676 136037
rect 89236 134830 89266 135210
rect 89646 134830 89676 135210
rect 89236 134611 89676 134830
rect 89236 134525 89329 134611
rect 89415 134525 89497 134611
rect 89583 134525 89676 134611
rect 89236 133099 89676 134525
rect 89236 133013 89329 133099
rect 89415 133013 89497 133099
rect 89583 133013 89676 133099
rect 89236 131587 89676 133013
rect 89236 131501 89329 131587
rect 89415 131501 89497 131587
rect 89583 131501 89676 131587
rect 89236 130075 89676 131501
rect 89236 129989 89329 130075
rect 89415 129989 89497 130075
rect 89583 129989 89676 130075
rect 89236 128563 89676 129989
rect 89236 128477 89329 128563
rect 89415 128477 89497 128563
rect 89583 128477 89676 128563
rect 89236 127051 89676 128477
rect 89236 126965 89329 127051
rect 89415 126965 89497 127051
rect 89583 126965 89676 127051
rect 89236 125539 89676 126965
rect 89236 125453 89329 125539
rect 89415 125453 89497 125539
rect 89583 125453 89676 125539
rect 89236 124027 89676 125453
rect 89236 123941 89329 124027
rect 89415 123941 89497 124027
rect 89583 123941 89676 124027
rect 89236 122515 89676 123941
rect 89236 122429 89329 122515
rect 89415 122429 89497 122515
rect 89583 122429 89676 122515
rect 89236 121003 89676 122429
rect 89236 120917 89329 121003
rect 89415 120917 89497 121003
rect 89583 120917 89676 121003
rect 89236 120090 89676 120917
rect 89236 119710 89266 120090
rect 89646 119710 89676 120090
rect 89236 119491 89676 119710
rect 89236 119405 89329 119491
rect 89415 119405 89497 119491
rect 89583 119405 89676 119491
rect 89236 117979 89676 119405
rect 89236 117893 89329 117979
rect 89415 117893 89497 117979
rect 89583 117893 89676 117979
rect 89236 116467 89676 117893
rect 89236 116381 89329 116467
rect 89415 116381 89497 116467
rect 89583 116381 89676 116467
rect 89236 114955 89676 116381
rect 89236 114869 89329 114955
rect 89415 114869 89497 114955
rect 89583 114869 89676 114955
rect 89236 113443 89676 114869
rect 89236 113357 89329 113443
rect 89415 113357 89497 113443
rect 89583 113357 89676 113443
rect 89236 111931 89676 113357
rect 89236 111845 89329 111931
rect 89415 111845 89497 111931
rect 89583 111845 89676 111931
rect 89236 110419 89676 111845
rect 89236 110333 89329 110419
rect 89415 110333 89497 110419
rect 89583 110333 89676 110419
rect 89236 108907 89676 110333
rect 89236 108821 89329 108907
rect 89415 108821 89497 108907
rect 89583 108821 89676 108907
rect 89236 107395 89676 108821
rect 89236 107309 89329 107395
rect 89415 107309 89497 107395
rect 89583 107309 89676 107395
rect 89236 105883 89676 107309
rect 89236 105797 89329 105883
rect 89415 105797 89497 105883
rect 89583 105797 89676 105883
rect 89236 104970 89676 105797
rect 89236 104590 89266 104970
rect 89646 104590 89676 104970
rect 89236 104371 89676 104590
rect 89236 104285 89329 104371
rect 89415 104285 89497 104371
rect 89583 104285 89676 104371
rect 89236 102859 89676 104285
rect 89236 102773 89329 102859
rect 89415 102773 89497 102859
rect 89583 102773 89676 102859
rect 89236 101347 89676 102773
rect 89236 101261 89329 101347
rect 89415 101261 89497 101347
rect 89583 101261 89676 101347
rect 89236 99835 89676 101261
rect 89236 99749 89329 99835
rect 89415 99749 89497 99835
rect 89583 99749 89676 99835
rect 89236 98323 89676 99749
rect 89236 98237 89329 98323
rect 89415 98237 89497 98323
rect 89583 98237 89676 98323
rect 89236 96811 89676 98237
rect 89236 96725 89329 96811
rect 89415 96725 89497 96811
rect 89583 96725 89676 96811
rect 89236 95299 89676 96725
rect 89236 95213 89329 95299
rect 89415 95213 89497 95299
rect 89583 95213 89676 95299
rect 89236 93787 89676 95213
rect 89236 93701 89329 93787
rect 89415 93701 89497 93787
rect 89583 93701 89676 93787
rect 89236 92275 89676 93701
rect 89236 92189 89329 92275
rect 89415 92189 89497 92275
rect 89583 92189 89676 92275
rect 89236 90763 89676 92189
rect 89236 90677 89329 90763
rect 89415 90677 89497 90763
rect 89583 90677 89676 90763
rect 89236 89850 89676 90677
rect 89236 89470 89266 89850
rect 89646 89470 89676 89850
rect 89236 89251 89676 89470
rect 89236 89165 89329 89251
rect 89415 89165 89497 89251
rect 89583 89165 89676 89251
rect 89236 87739 89676 89165
rect 89236 87653 89329 87739
rect 89415 87653 89497 87739
rect 89583 87653 89676 87739
rect 89236 86227 89676 87653
rect 89236 86141 89329 86227
rect 89415 86141 89497 86227
rect 89583 86141 89676 86227
rect 89236 84715 89676 86141
rect 89236 84629 89329 84715
rect 89415 84629 89497 84715
rect 89583 84629 89676 84715
rect 89236 83203 89676 84629
rect 89236 83117 89329 83203
rect 89415 83117 89497 83203
rect 89583 83117 89676 83203
rect 89236 81691 89676 83117
rect 89236 81605 89329 81691
rect 89415 81605 89497 81691
rect 89583 81605 89676 81691
rect 89236 80179 89676 81605
rect 89236 80093 89329 80179
rect 89415 80093 89497 80179
rect 89583 80093 89676 80179
rect 89236 78667 89676 80093
rect 89236 78581 89329 78667
rect 89415 78581 89497 78667
rect 89583 78581 89676 78667
rect 89236 77155 89676 78581
rect 89236 77069 89329 77155
rect 89415 77069 89497 77155
rect 89583 77069 89676 77155
rect 89236 75643 89676 77069
rect 89236 75557 89329 75643
rect 89415 75557 89497 75643
rect 89583 75557 89676 75643
rect 89236 74730 89676 75557
rect 89236 74350 89266 74730
rect 89646 74350 89676 74730
rect 89236 74131 89676 74350
rect 89236 74045 89329 74131
rect 89415 74045 89497 74131
rect 89583 74045 89676 74131
rect 89236 72619 89676 74045
rect 89236 72533 89329 72619
rect 89415 72533 89497 72619
rect 89583 72533 89676 72619
rect 89236 70806 89676 72533
rect 89236 70426 89266 70806
rect 89646 70426 89676 70806
rect 89236 70414 89676 70426
rect 89236 70034 89266 70414
rect 89646 70034 89676 70414
rect 89236 68520 89676 70034
rect 90476 155142 90916 155256
rect 90476 154762 90506 155142
rect 90886 154762 90916 155142
rect 90476 154750 90916 154762
rect 90476 154370 90506 154750
rect 90886 154370 90916 154750
rect 90476 151999 90916 154370
rect 90476 151913 90569 151999
rect 90655 151913 90737 151999
rect 90823 151913 90916 151999
rect 90476 151570 90916 151913
rect 90476 151190 90506 151570
rect 90886 151190 90916 151570
rect 90476 150487 90916 151190
rect 90476 150401 90569 150487
rect 90655 150401 90737 150487
rect 90823 150401 90916 150487
rect 90476 148975 90916 150401
rect 90476 148889 90569 148975
rect 90655 148889 90737 148975
rect 90823 148889 90916 148975
rect 90476 147463 90916 148889
rect 90476 147377 90569 147463
rect 90655 147377 90737 147463
rect 90823 147377 90916 147463
rect 90476 145951 90916 147377
rect 90476 145865 90569 145951
rect 90655 145865 90737 145951
rect 90823 145865 90916 145951
rect 90476 144439 90916 145865
rect 90476 144353 90569 144439
rect 90655 144353 90737 144439
rect 90823 144353 90916 144439
rect 90476 142927 90916 144353
rect 90476 142841 90569 142927
rect 90655 142841 90737 142927
rect 90823 142841 90916 142927
rect 90476 141415 90916 142841
rect 90476 141329 90569 141415
rect 90655 141329 90737 141415
rect 90823 141329 90916 141415
rect 90476 139903 90916 141329
rect 90476 139817 90569 139903
rect 90655 139817 90737 139903
rect 90823 139817 90916 139903
rect 90476 138391 90916 139817
rect 90476 138305 90569 138391
rect 90655 138305 90737 138391
rect 90823 138305 90916 138391
rect 90476 136879 90916 138305
rect 90476 136793 90569 136879
rect 90655 136793 90737 136879
rect 90823 136793 90916 136879
rect 90476 136450 90916 136793
rect 90476 136070 90506 136450
rect 90886 136070 90916 136450
rect 90476 135367 90916 136070
rect 90476 135281 90569 135367
rect 90655 135281 90737 135367
rect 90823 135281 90916 135367
rect 90476 133855 90916 135281
rect 90476 133769 90569 133855
rect 90655 133769 90737 133855
rect 90823 133769 90916 133855
rect 90476 132343 90916 133769
rect 90476 132257 90569 132343
rect 90655 132257 90737 132343
rect 90823 132257 90916 132343
rect 90476 130831 90916 132257
rect 90476 130745 90569 130831
rect 90655 130745 90737 130831
rect 90823 130745 90916 130831
rect 90476 129319 90916 130745
rect 90476 129233 90569 129319
rect 90655 129233 90737 129319
rect 90823 129233 90916 129319
rect 90476 127807 90916 129233
rect 90476 127721 90569 127807
rect 90655 127721 90737 127807
rect 90823 127721 90916 127807
rect 90476 126295 90916 127721
rect 90476 126209 90569 126295
rect 90655 126209 90737 126295
rect 90823 126209 90916 126295
rect 90476 124783 90916 126209
rect 90476 124697 90569 124783
rect 90655 124697 90737 124783
rect 90823 124697 90916 124783
rect 90476 123271 90916 124697
rect 90476 123185 90569 123271
rect 90655 123185 90737 123271
rect 90823 123185 90916 123271
rect 90476 121759 90916 123185
rect 90476 121673 90569 121759
rect 90655 121673 90737 121759
rect 90823 121673 90916 121759
rect 90476 121330 90916 121673
rect 90476 120950 90506 121330
rect 90886 120950 90916 121330
rect 90476 120247 90916 120950
rect 90476 120161 90569 120247
rect 90655 120161 90737 120247
rect 90823 120161 90916 120247
rect 90476 118735 90916 120161
rect 90476 118649 90569 118735
rect 90655 118649 90737 118735
rect 90823 118649 90916 118735
rect 90476 117223 90916 118649
rect 90476 117137 90569 117223
rect 90655 117137 90737 117223
rect 90823 117137 90916 117223
rect 90476 115711 90916 117137
rect 90476 115625 90569 115711
rect 90655 115625 90737 115711
rect 90823 115625 90916 115711
rect 90476 114199 90916 115625
rect 90476 114113 90569 114199
rect 90655 114113 90737 114199
rect 90823 114113 90916 114199
rect 90476 112687 90916 114113
rect 90476 112601 90569 112687
rect 90655 112601 90737 112687
rect 90823 112601 90916 112687
rect 90476 111175 90916 112601
rect 90476 111089 90569 111175
rect 90655 111089 90737 111175
rect 90823 111089 90916 111175
rect 90476 109663 90916 111089
rect 90476 109577 90569 109663
rect 90655 109577 90737 109663
rect 90823 109577 90916 109663
rect 90476 108151 90916 109577
rect 90476 108065 90569 108151
rect 90655 108065 90737 108151
rect 90823 108065 90916 108151
rect 90476 106639 90916 108065
rect 90476 106553 90569 106639
rect 90655 106553 90737 106639
rect 90823 106553 90916 106639
rect 90476 106210 90916 106553
rect 90476 105830 90506 106210
rect 90886 105830 90916 106210
rect 90476 105127 90916 105830
rect 90476 105041 90569 105127
rect 90655 105041 90737 105127
rect 90823 105041 90916 105127
rect 90476 103615 90916 105041
rect 90476 103529 90569 103615
rect 90655 103529 90737 103615
rect 90823 103529 90916 103615
rect 90476 102103 90916 103529
rect 90476 102017 90569 102103
rect 90655 102017 90737 102103
rect 90823 102017 90916 102103
rect 90476 100591 90916 102017
rect 90476 100505 90569 100591
rect 90655 100505 90737 100591
rect 90823 100505 90916 100591
rect 90476 99079 90916 100505
rect 90476 98993 90569 99079
rect 90655 98993 90737 99079
rect 90823 98993 90916 99079
rect 90476 97567 90916 98993
rect 90476 97481 90569 97567
rect 90655 97481 90737 97567
rect 90823 97481 90916 97567
rect 90476 96055 90916 97481
rect 90476 95969 90569 96055
rect 90655 95969 90737 96055
rect 90823 95969 90916 96055
rect 90476 94543 90916 95969
rect 90476 94457 90569 94543
rect 90655 94457 90737 94543
rect 90823 94457 90916 94543
rect 90476 93031 90916 94457
rect 90476 92945 90569 93031
rect 90655 92945 90737 93031
rect 90823 92945 90916 93031
rect 90476 91519 90916 92945
rect 90476 91433 90569 91519
rect 90655 91433 90737 91519
rect 90823 91433 90916 91519
rect 90476 91090 90916 91433
rect 90476 90710 90506 91090
rect 90886 90710 90916 91090
rect 90476 90007 90916 90710
rect 90476 89921 90569 90007
rect 90655 89921 90737 90007
rect 90823 89921 90916 90007
rect 90476 88495 90916 89921
rect 90476 88409 90569 88495
rect 90655 88409 90737 88495
rect 90823 88409 90916 88495
rect 90476 86983 90916 88409
rect 90476 86897 90569 86983
rect 90655 86897 90737 86983
rect 90823 86897 90916 86983
rect 90476 85471 90916 86897
rect 90476 85385 90569 85471
rect 90655 85385 90737 85471
rect 90823 85385 90916 85471
rect 90476 83959 90916 85385
rect 90476 83873 90569 83959
rect 90655 83873 90737 83959
rect 90823 83873 90916 83959
rect 90476 82447 90916 83873
rect 90476 82361 90569 82447
rect 90655 82361 90737 82447
rect 90823 82361 90916 82447
rect 90476 80935 90916 82361
rect 90476 80849 90569 80935
rect 90655 80849 90737 80935
rect 90823 80849 90916 80935
rect 90476 79423 90916 80849
rect 90476 79337 90569 79423
rect 90655 79337 90737 79423
rect 90823 79337 90916 79423
rect 90476 77911 90916 79337
rect 90476 77825 90569 77911
rect 90655 77825 90737 77911
rect 90823 77825 90916 77911
rect 90476 76399 90916 77825
rect 90476 76313 90569 76399
rect 90655 76313 90737 76399
rect 90823 76313 90916 76399
rect 90476 75970 90916 76313
rect 90476 75590 90506 75970
rect 90886 75590 90916 75970
rect 90476 74887 90916 75590
rect 90476 74801 90569 74887
rect 90655 74801 90737 74887
rect 90823 74801 90916 74887
rect 90476 73375 90916 74801
rect 90476 73289 90569 73375
rect 90655 73289 90737 73375
rect 90823 73289 90916 73375
rect 90476 71863 90916 73289
rect 90476 71777 90569 71863
rect 90655 71777 90737 71863
rect 90823 71777 90916 71863
rect 90476 69406 90916 71777
rect 90476 69026 90506 69406
rect 90886 69026 90916 69406
rect 90476 69014 90916 69026
rect 90476 68634 90506 69014
rect 90886 68634 90916 69014
rect 90476 68520 90916 68634
rect 104356 153742 104796 155256
rect 104356 153362 104386 153742
rect 104766 153362 104796 153742
rect 104356 153350 104796 153362
rect 104356 152970 104386 153350
rect 104766 152970 104796 153350
rect 104356 151243 104796 152970
rect 104356 151157 104449 151243
rect 104535 151157 104617 151243
rect 104703 151157 104796 151243
rect 104356 150330 104796 151157
rect 104356 149950 104386 150330
rect 104766 149950 104796 150330
rect 104356 149731 104796 149950
rect 104356 149645 104449 149731
rect 104535 149645 104617 149731
rect 104703 149645 104796 149731
rect 104356 148219 104796 149645
rect 104356 148133 104449 148219
rect 104535 148133 104617 148219
rect 104703 148133 104796 148219
rect 104356 146707 104796 148133
rect 104356 146621 104449 146707
rect 104535 146621 104617 146707
rect 104703 146621 104796 146707
rect 104356 145195 104796 146621
rect 104356 145109 104449 145195
rect 104535 145109 104617 145195
rect 104703 145109 104796 145195
rect 104356 143683 104796 145109
rect 104356 143597 104449 143683
rect 104535 143597 104617 143683
rect 104703 143597 104796 143683
rect 104356 142171 104796 143597
rect 104356 142085 104449 142171
rect 104535 142085 104617 142171
rect 104703 142085 104796 142171
rect 104356 140659 104796 142085
rect 104356 140573 104449 140659
rect 104535 140573 104617 140659
rect 104703 140573 104796 140659
rect 104356 139147 104796 140573
rect 104356 139061 104449 139147
rect 104535 139061 104617 139147
rect 104703 139061 104796 139147
rect 104356 137635 104796 139061
rect 104356 137549 104449 137635
rect 104535 137549 104617 137635
rect 104703 137549 104796 137635
rect 104356 136123 104796 137549
rect 104356 136037 104449 136123
rect 104535 136037 104617 136123
rect 104703 136037 104796 136123
rect 104356 135210 104796 136037
rect 104356 134830 104386 135210
rect 104766 134830 104796 135210
rect 104356 134611 104796 134830
rect 104356 134525 104449 134611
rect 104535 134525 104617 134611
rect 104703 134525 104796 134611
rect 104356 133099 104796 134525
rect 104356 133013 104449 133099
rect 104535 133013 104617 133099
rect 104703 133013 104796 133099
rect 104356 131587 104796 133013
rect 104356 131501 104449 131587
rect 104535 131501 104617 131587
rect 104703 131501 104796 131587
rect 104356 130075 104796 131501
rect 104356 129989 104449 130075
rect 104535 129989 104617 130075
rect 104703 129989 104796 130075
rect 104356 128563 104796 129989
rect 104356 128477 104449 128563
rect 104535 128477 104617 128563
rect 104703 128477 104796 128563
rect 104356 127051 104796 128477
rect 104356 126965 104449 127051
rect 104535 126965 104617 127051
rect 104703 126965 104796 127051
rect 104356 125539 104796 126965
rect 104356 125453 104449 125539
rect 104535 125453 104617 125539
rect 104703 125453 104796 125539
rect 104356 124027 104796 125453
rect 104356 123941 104449 124027
rect 104535 123941 104617 124027
rect 104703 123941 104796 124027
rect 104356 122515 104796 123941
rect 104356 122429 104449 122515
rect 104535 122429 104617 122515
rect 104703 122429 104796 122515
rect 104356 121003 104796 122429
rect 104356 120917 104449 121003
rect 104535 120917 104617 121003
rect 104703 120917 104796 121003
rect 104356 120090 104796 120917
rect 104356 119710 104386 120090
rect 104766 119710 104796 120090
rect 104356 119491 104796 119710
rect 104356 119405 104449 119491
rect 104535 119405 104617 119491
rect 104703 119405 104796 119491
rect 104356 117979 104796 119405
rect 104356 117893 104449 117979
rect 104535 117893 104617 117979
rect 104703 117893 104796 117979
rect 104356 116467 104796 117893
rect 104356 116381 104449 116467
rect 104535 116381 104617 116467
rect 104703 116381 104796 116467
rect 104356 114955 104796 116381
rect 104356 114869 104449 114955
rect 104535 114869 104617 114955
rect 104703 114869 104796 114955
rect 104356 113443 104796 114869
rect 104356 113357 104449 113443
rect 104535 113357 104617 113443
rect 104703 113357 104796 113443
rect 104356 111931 104796 113357
rect 104356 111845 104449 111931
rect 104535 111845 104617 111931
rect 104703 111845 104796 111931
rect 104356 110419 104796 111845
rect 104356 110333 104449 110419
rect 104535 110333 104617 110419
rect 104703 110333 104796 110419
rect 104356 108907 104796 110333
rect 104356 108821 104449 108907
rect 104535 108821 104617 108907
rect 104703 108821 104796 108907
rect 104356 107395 104796 108821
rect 104356 107309 104449 107395
rect 104535 107309 104617 107395
rect 104703 107309 104796 107395
rect 104356 105883 104796 107309
rect 104356 105797 104449 105883
rect 104535 105797 104617 105883
rect 104703 105797 104796 105883
rect 104356 104970 104796 105797
rect 104356 104590 104386 104970
rect 104766 104590 104796 104970
rect 104356 104371 104796 104590
rect 104356 104285 104449 104371
rect 104535 104285 104617 104371
rect 104703 104285 104796 104371
rect 104356 102859 104796 104285
rect 104356 102773 104449 102859
rect 104535 102773 104617 102859
rect 104703 102773 104796 102859
rect 104356 101347 104796 102773
rect 104356 101261 104449 101347
rect 104535 101261 104617 101347
rect 104703 101261 104796 101347
rect 104356 99835 104796 101261
rect 104356 99749 104449 99835
rect 104535 99749 104617 99835
rect 104703 99749 104796 99835
rect 104356 98323 104796 99749
rect 104356 98237 104449 98323
rect 104535 98237 104617 98323
rect 104703 98237 104796 98323
rect 104356 96811 104796 98237
rect 104356 96725 104449 96811
rect 104535 96725 104617 96811
rect 104703 96725 104796 96811
rect 104356 95299 104796 96725
rect 104356 95213 104449 95299
rect 104535 95213 104617 95299
rect 104703 95213 104796 95299
rect 104356 93787 104796 95213
rect 104356 93701 104449 93787
rect 104535 93701 104617 93787
rect 104703 93701 104796 93787
rect 104356 92275 104796 93701
rect 104356 92189 104449 92275
rect 104535 92189 104617 92275
rect 104703 92189 104796 92275
rect 104356 90763 104796 92189
rect 104356 90677 104449 90763
rect 104535 90677 104617 90763
rect 104703 90677 104796 90763
rect 104356 89850 104796 90677
rect 104356 89470 104386 89850
rect 104766 89470 104796 89850
rect 104356 89251 104796 89470
rect 104356 89165 104449 89251
rect 104535 89165 104617 89251
rect 104703 89165 104796 89251
rect 104356 87739 104796 89165
rect 104356 87653 104449 87739
rect 104535 87653 104617 87739
rect 104703 87653 104796 87739
rect 104356 86227 104796 87653
rect 104356 86141 104449 86227
rect 104535 86141 104617 86227
rect 104703 86141 104796 86227
rect 104356 84715 104796 86141
rect 104356 84629 104449 84715
rect 104535 84629 104617 84715
rect 104703 84629 104796 84715
rect 104356 83203 104796 84629
rect 104356 83117 104449 83203
rect 104535 83117 104617 83203
rect 104703 83117 104796 83203
rect 104356 81691 104796 83117
rect 104356 81605 104449 81691
rect 104535 81605 104617 81691
rect 104703 81605 104796 81691
rect 104356 80179 104796 81605
rect 104356 80093 104449 80179
rect 104535 80093 104617 80179
rect 104703 80093 104796 80179
rect 104356 78667 104796 80093
rect 104356 78581 104449 78667
rect 104535 78581 104617 78667
rect 104703 78581 104796 78667
rect 104356 77155 104796 78581
rect 104356 77069 104449 77155
rect 104535 77069 104617 77155
rect 104703 77069 104796 77155
rect 104356 75643 104796 77069
rect 104356 75557 104449 75643
rect 104535 75557 104617 75643
rect 104703 75557 104796 75643
rect 104356 74730 104796 75557
rect 104356 74350 104386 74730
rect 104766 74350 104796 74730
rect 104356 74131 104796 74350
rect 104356 74045 104449 74131
rect 104535 74045 104617 74131
rect 104703 74045 104796 74131
rect 104356 72619 104796 74045
rect 104356 72533 104449 72619
rect 104535 72533 104617 72619
rect 104703 72533 104796 72619
rect 104356 70806 104796 72533
rect 104356 70426 104386 70806
rect 104766 70426 104796 70806
rect 104356 70414 104796 70426
rect 104356 70034 104386 70414
rect 104766 70034 104796 70414
rect 104356 68520 104796 70034
rect 105596 155142 106036 155256
rect 105596 154762 105626 155142
rect 106006 154762 106036 155142
rect 105596 154750 106036 154762
rect 105596 154370 105626 154750
rect 106006 154370 106036 154750
rect 105596 151999 106036 154370
rect 105596 151913 105689 151999
rect 105775 151913 105857 151999
rect 105943 151913 106036 151999
rect 105596 151570 106036 151913
rect 105596 151190 105626 151570
rect 106006 151190 106036 151570
rect 105596 150487 106036 151190
rect 105596 150401 105689 150487
rect 105775 150401 105857 150487
rect 105943 150401 106036 150487
rect 105596 148975 106036 150401
rect 105596 148889 105689 148975
rect 105775 148889 105857 148975
rect 105943 148889 106036 148975
rect 105596 147463 106036 148889
rect 105596 147377 105689 147463
rect 105775 147377 105857 147463
rect 105943 147377 106036 147463
rect 105596 145951 106036 147377
rect 105596 145865 105689 145951
rect 105775 145865 105857 145951
rect 105943 145865 106036 145951
rect 105596 144439 106036 145865
rect 105596 144353 105689 144439
rect 105775 144353 105857 144439
rect 105943 144353 106036 144439
rect 105596 142927 106036 144353
rect 105596 142841 105689 142927
rect 105775 142841 105857 142927
rect 105943 142841 106036 142927
rect 105596 141415 106036 142841
rect 105596 141329 105689 141415
rect 105775 141329 105857 141415
rect 105943 141329 106036 141415
rect 105596 139903 106036 141329
rect 105596 139817 105689 139903
rect 105775 139817 105857 139903
rect 105943 139817 106036 139903
rect 105596 138391 106036 139817
rect 105596 138305 105689 138391
rect 105775 138305 105857 138391
rect 105943 138305 106036 138391
rect 105596 136879 106036 138305
rect 105596 136793 105689 136879
rect 105775 136793 105857 136879
rect 105943 136793 106036 136879
rect 105596 136450 106036 136793
rect 105596 136070 105626 136450
rect 106006 136070 106036 136450
rect 105596 135367 106036 136070
rect 105596 135281 105689 135367
rect 105775 135281 105857 135367
rect 105943 135281 106036 135367
rect 105596 133855 106036 135281
rect 105596 133769 105689 133855
rect 105775 133769 105857 133855
rect 105943 133769 106036 133855
rect 105596 132343 106036 133769
rect 105596 132257 105689 132343
rect 105775 132257 105857 132343
rect 105943 132257 106036 132343
rect 105596 130831 106036 132257
rect 105596 130745 105689 130831
rect 105775 130745 105857 130831
rect 105943 130745 106036 130831
rect 105596 129319 106036 130745
rect 105596 129233 105689 129319
rect 105775 129233 105857 129319
rect 105943 129233 106036 129319
rect 105596 127807 106036 129233
rect 105596 127721 105689 127807
rect 105775 127721 105857 127807
rect 105943 127721 106036 127807
rect 105596 126295 106036 127721
rect 105596 126209 105689 126295
rect 105775 126209 105857 126295
rect 105943 126209 106036 126295
rect 105596 124783 106036 126209
rect 105596 124697 105689 124783
rect 105775 124697 105857 124783
rect 105943 124697 106036 124783
rect 105596 123271 106036 124697
rect 105596 123185 105689 123271
rect 105775 123185 105857 123271
rect 105943 123185 106036 123271
rect 105596 121759 106036 123185
rect 105596 121673 105689 121759
rect 105775 121673 105857 121759
rect 105943 121673 106036 121759
rect 105596 121330 106036 121673
rect 105596 120950 105626 121330
rect 106006 120950 106036 121330
rect 105596 120247 106036 120950
rect 105596 120161 105689 120247
rect 105775 120161 105857 120247
rect 105943 120161 106036 120247
rect 105596 118735 106036 120161
rect 105596 118649 105689 118735
rect 105775 118649 105857 118735
rect 105943 118649 106036 118735
rect 105596 117223 106036 118649
rect 105596 117137 105689 117223
rect 105775 117137 105857 117223
rect 105943 117137 106036 117223
rect 105596 115711 106036 117137
rect 105596 115625 105689 115711
rect 105775 115625 105857 115711
rect 105943 115625 106036 115711
rect 105596 114199 106036 115625
rect 105596 114113 105689 114199
rect 105775 114113 105857 114199
rect 105943 114113 106036 114199
rect 105596 112687 106036 114113
rect 105596 112601 105689 112687
rect 105775 112601 105857 112687
rect 105943 112601 106036 112687
rect 105596 111175 106036 112601
rect 105596 111089 105689 111175
rect 105775 111089 105857 111175
rect 105943 111089 106036 111175
rect 105596 109663 106036 111089
rect 105596 109577 105689 109663
rect 105775 109577 105857 109663
rect 105943 109577 106036 109663
rect 105596 108151 106036 109577
rect 105596 108065 105689 108151
rect 105775 108065 105857 108151
rect 105943 108065 106036 108151
rect 105596 106639 106036 108065
rect 105596 106553 105689 106639
rect 105775 106553 105857 106639
rect 105943 106553 106036 106639
rect 105596 106210 106036 106553
rect 105596 105830 105626 106210
rect 106006 105830 106036 106210
rect 105596 105127 106036 105830
rect 105596 105041 105689 105127
rect 105775 105041 105857 105127
rect 105943 105041 106036 105127
rect 105596 103615 106036 105041
rect 105596 103529 105689 103615
rect 105775 103529 105857 103615
rect 105943 103529 106036 103615
rect 105596 102103 106036 103529
rect 105596 102017 105689 102103
rect 105775 102017 105857 102103
rect 105943 102017 106036 102103
rect 105596 100591 106036 102017
rect 105596 100505 105689 100591
rect 105775 100505 105857 100591
rect 105943 100505 106036 100591
rect 105596 99079 106036 100505
rect 105596 98993 105689 99079
rect 105775 98993 105857 99079
rect 105943 98993 106036 99079
rect 105596 97567 106036 98993
rect 105596 97481 105689 97567
rect 105775 97481 105857 97567
rect 105943 97481 106036 97567
rect 105596 96055 106036 97481
rect 105596 95969 105689 96055
rect 105775 95969 105857 96055
rect 105943 95969 106036 96055
rect 105596 94543 106036 95969
rect 105596 94457 105689 94543
rect 105775 94457 105857 94543
rect 105943 94457 106036 94543
rect 105596 93031 106036 94457
rect 105596 92945 105689 93031
rect 105775 92945 105857 93031
rect 105943 92945 106036 93031
rect 105596 91519 106036 92945
rect 105596 91433 105689 91519
rect 105775 91433 105857 91519
rect 105943 91433 106036 91519
rect 105596 91090 106036 91433
rect 105596 90710 105626 91090
rect 106006 90710 106036 91090
rect 105596 90007 106036 90710
rect 105596 89921 105689 90007
rect 105775 89921 105857 90007
rect 105943 89921 106036 90007
rect 105596 88495 106036 89921
rect 105596 88409 105689 88495
rect 105775 88409 105857 88495
rect 105943 88409 106036 88495
rect 105596 86983 106036 88409
rect 105596 86897 105689 86983
rect 105775 86897 105857 86983
rect 105943 86897 106036 86983
rect 105596 85471 106036 86897
rect 105596 85385 105689 85471
rect 105775 85385 105857 85471
rect 105943 85385 106036 85471
rect 105596 83959 106036 85385
rect 105596 83873 105689 83959
rect 105775 83873 105857 83959
rect 105943 83873 106036 83959
rect 105596 82447 106036 83873
rect 105596 82361 105689 82447
rect 105775 82361 105857 82447
rect 105943 82361 106036 82447
rect 105596 80935 106036 82361
rect 105596 80849 105689 80935
rect 105775 80849 105857 80935
rect 105943 80849 106036 80935
rect 105596 79423 106036 80849
rect 105596 79337 105689 79423
rect 105775 79337 105857 79423
rect 105943 79337 106036 79423
rect 105596 77911 106036 79337
rect 105596 77825 105689 77911
rect 105775 77825 105857 77911
rect 105943 77825 106036 77911
rect 105596 76399 106036 77825
rect 105596 76313 105689 76399
rect 105775 76313 105857 76399
rect 105943 76313 106036 76399
rect 105596 75970 106036 76313
rect 105596 75590 105626 75970
rect 106006 75590 106036 75970
rect 105596 74887 106036 75590
rect 105596 74801 105689 74887
rect 105775 74801 105857 74887
rect 105943 74801 106036 74887
rect 105596 73375 106036 74801
rect 105596 73289 105689 73375
rect 105775 73289 105857 73375
rect 105943 73289 106036 73375
rect 105596 71863 106036 73289
rect 105596 71777 105689 71863
rect 105775 71777 105857 71863
rect 105943 71777 106036 71863
rect 105596 69406 106036 71777
rect 105596 69026 105626 69406
rect 106006 69026 106036 69406
rect 105596 69014 106036 69026
rect 105596 68634 105626 69014
rect 106006 68634 106036 69014
rect 105596 68520 106036 68634
rect 119476 153742 119916 155256
rect 119476 153362 119506 153742
rect 119886 153362 119916 153742
rect 119476 153350 119916 153362
rect 119476 152970 119506 153350
rect 119886 152970 119916 153350
rect 119476 151243 119916 152970
rect 119476 151157 119569 151243
rect 119655 151157 119737 151243
rect 119823 151157 119916 151243
rect 119476 150330 119916 151157
rect 119476 149950 119506 150330
rect 119886 149950 119916 150330
rect 119476 149731 119916 149950
rect 119476 149645 119569 149731
rect 119655 149645 119737 149731
rect 119823 149645 119916 149731
rect 119476 148219 119916 149645
rect 119476 148133 119569 148219
rect 119655 148133 119737 148219
rect 119823 148133 119916 148219
rect 119476 146707 119916 148133
rect 119476 146621 119569 146707
rect 119655 146621 119737 146707
rect 119823 146621 119916 146707
rect 119476 145195 119916 146621
rect 119476 145109 119569 145195
rect 119655 145109 119737 145195
rect 119823 145109 119916 145195
rect 119476 143683 119916 145109
rect 119476 143597 119569 143683
rect 119655 143597 119737 143683
rect 119823 143597 119916 143683
rect 119476 142171 119916 143597
rect 119476 142085 119569 142171
rect 119655 142085 119737 142171
rect 119823 142085 119916 142171
rect 119476 140659 119916 142085
rect 119476 140573 119569 140659
rect 119655 140573 119737 140659
rect 119823 140573 119916 140659
rect 119476 139147 119916 140573
rect 119476 139061 119569 139147
rect 119655 139061 119737 139147
rect 119823 139061 119916 139147
rect 119476 137635 119916 139061
rect 119476 137549 119569 137635
rect 119655 137549 119737 137635
rect 119823 137549 119916 137635
rect 119476 136123 119916 137549
rect 119476 136037 119569 136123
rect 119655 136037 119737 136123
rect 119823 136037 119916 136123
rect 119476 135210 119916 136037
rect 119476 134830 119506 135210
rect 119886 134830 119916 135210
rect 119476 134611 119916 134830
rect 119476 134525 119569 134611
rect 119655 134525 119737 134611
rect 119823 134525 119916 134611
rect 119476 133099 119916 134525
rect 119476 133013 119569 133099
rect 119655 133013 119737 133099
rect 119823 133013 119916 133099
rect 119476 131587 119916 133013
rect 119476 131501 119569 131587
rect 119655 131501 119737 131587
rect 119823 131501 119916 131587
rect 119476 130075 119916 131501
rect 119476 129989 119569 130075
rect 119655 129989 119737 130075
rect 119823 129989 119916 130075
rect 119476 128563 119916 129989
rect 119476 128477 119569 128563
rect 119655 128477 119737 128563
rect 119823 128477 119916 128563
rect 119476 127051 119916 128477
rect 119476 126965 119569 127051
rect 119655 126965 119737 127051
rect 119823 126965 119916 127051
rect 119476 125539 119916 126965
rect 119476 125453 119569 125539
rect 119655 125453 119737 125539
rect 119823 125453 119916 125539
rect 119476 124027 119916 125453
rect 119476 123941 119569 124027
rect 119655 123941 119737 124027
rect 119823 123941 119916 124027
rect 119476 122515 119916 123941
rect 119476 122429 119569 122515
rect 119655 122429 119737 122515
rect 119823 122429 119916 122515
rect 119476 121003 119916 122429
rect 119476 120917 119569 121003
rect 119655 120917 119737 121003
rect 119823 120917 119916 121003
rect 119476 120090 119916 120917
rect 119476 119710 119506 120090
rect 119886 119710 119916 120090
rect 119476 119491 119916 119710
rect 119476 119405 119569 119491
rect 119655 119405 119737 119491
rect 119823 119405 119916 119491
rect 119476 117979 119916 119405
rect 119476 117893 119569 117979
rect 119655 117893 119737 117979
rect 119823 117893 119916 117979
rect 119476 116467 119916 117893
rect 119476 116381 119569 116467
rect 119655 116381 119737 116467
rect 119823 116381 119916 116467
rect 119476 114955 119916 116381
rect 119476 114869 119569 114955
rect 119655 114869 119737 114955
rect 119823 114869 119916 114955
rect 119476 113443 119916 114869
rect 119476 113357 119569 113443
rect 119655 113357 119737 113443
rect 119823 113357 119916 113443
rect 119476 111931 119916 113357
rect 119476 111845 119569 111931
rect 119655 111845 119737 111931
rect 119823 111845 119916 111931
rect 119476 110419 119916 111845
rect 119476 110333 119569 110419
rect 119655 110333 119737 110419
rect 119823 110333 119916 110419
rect 119476 108907 119916 110333
rect 119476 108821 119569 108907
rect 119655 108821 119737 108907
rect 119823 108821 119916 108907
rect 119476 107395 119916 108821
rect 119476 107309 119569 107395
rect 119655 107309 119737 107395
rect 119823 107309 119916 107395
rect 119476 105883 119916 107309
rect 119476 105797 119569 105883
rect 119655 105797 119737 105883
rect 119823 105797 119916 105883
rect 119476 104970 119916 105797
rect 119476 104590 119506 104970
rect 119886 104590 119916 104970
rect 119476 104371 119916 104590
rect 119476 104285 119569 104371
rect 119655 104285 119737 104371
rect 119823 104285 119916 104371
rect 119476 102859 119916 104285
rect 119476 102773 119569 102859
rect 119655 102773 119737 102859
rect 119823 102773 119916 102859
rect 119476 101347 119916 102773
rect 119476 101261 119569 101347
rect 119655 101261 119737 101347
rect 119823 101261 119916 101347
rect 119476 99835 119916 101261
rect 119476 99749 119569 99835
rect 119655 99749 119737 99835
rect 119823 99749 119916 99835
rect 119476 98323 119916 99749
rect 119476 98237 119569 98323
rect 119655 98237 119737 98323
rect 119823 98237 119916 98323
rect 119476 96811 119916 98237
rect 119476 96725 119569 96811
rect 119655 96725 119737 96811
rect 119823 96725 119916 96811
rect 119476 95299 119916 96725
rect 119476 95213 119569 95299
rect 119655 95213 119737 95299
rect 119823 95213 119916 95299
rect 119476 93787 119916 95213
rect 119476 93701 119569 93787
rect 119655 93701 119737 93787
rect 119823 93701 119916 93787
rect 119476 92275 119916 93701
rect 119476 92189 119569 92275
rect 119655 92189 119737 92275
rect 119823 92189 119916 92275
rect 119476 90763 119916 92189
rect 119476 90677 119569 90763
rect 119655 90677 119737 90763
rect 119823 90677 119916 90763
rect 119476 89850 119916 90677
rect 119476 89470 119506 89850
rect 119886 89470 119916 89850
rect 119476 89251 119916 89470
rect 119476 89165 119569 89251
rect 119655 89165 119737 89251
rect 119823 89165 119916 89251
rect 119476 87739 119916 89165
rect 119476 87653 119569 87739
rect 119655 87653 119737 87739
rect 119823 87653 119916 87739
rect 119476 86227 119916 87653
rect 119476 86141 119569 86227
rect 119655 86141 119737 86227
rect 119823 86141 119916 86227
rect 119476 84715 119916 86141
rect 119476 84629 119569 84715
rect 119655 84629 119737 84715
rect 119823 84629 119916 84715
rect 119476 83203 119916 84629
rect 119476 83117 119569 83203
rect 119655 83117 119737 83203
rect 119823 83117 119916 83203
rect 119476 81691 119916 83117
rect 119476 81605 119569 81691
rect 119655 81605 119737 81691
rect 119823 81605 119916 81691
rect 119476 80179 119916 81605
rect 119476 80093 119569 80179
rect 119655 80093 119737 80179
rect 119823 80093 119916 80179
rect 119476 78667 119916 80093
rect 119476 78581 119569 78667
rect 119655 78581 119737 78667
rect 119823 78581 119916 78667
rect 119476 77155 119916 78581
rect 119476 77069 119569 77155
rect 119655 77069 119737 77155
rect 119823 77069 119916 77155
rect 119476 75643 119916 77069
rect 119476 75557 119569 75643
rect 119655 75557 119737 75643
rect 119823 75557 119916 75643
rect 119476 74730 119916 75557
rect 119476 74350 119506 74730
rect 119886 74350 119916 74730
rect 119476 74131 119916 74350
rect 119476 74045 119569 74131
rect 119655 74045 119737 74131
rect 119823 74045 119916 74131
rect 119476 72619 119916 74045
rect 119476 72533 119569 72619
rect 119655 72533 119737 72619
rect 119823 72533 119916 72619
rect 119476 70806 119916 72533
rect 119476 70426 119506 70806
rect 119886 70426 119916 70806
rect 119476 70414 119916 70426
rect 119476 70034 119506 70414
rect 119886 70034 119916 70414
rect 119476 68520 119916 70034
rect 120716 155142 121156 155256
rect 120716 154762 120746 155142
rect 121126 154762 121156 155142
rect 120716 154750 121156 154762
rect 120716 154370 120746 154750
rect 121126 154370 121156 154750
rect 120716 151999 121156 154370
rect 120716 151913 120809 151999
rect 120895 151913 120977 151999
rect 121063 151913 121156 151999
rect 120716 151570 121156 151913
rect 120716 151190 120746 151570
rect 121126 151190 121156 151570
rect 120716 150487 121156 151190
rect 120716 150401 120809 150487
rect 120895 150401 120977 150487
rect 121063 150401 121156 150487
rect 120716 148975 121156 150401
rect 120716 148889 120809 148975
rect 120895 148889 120977 148975
rect 121063 148889 121156 148975
rect 120716 147463 121156 148889
rect 120716 147377 120809 147463
rect 120895 147377 120977 147463
rect 121063 147377 121156 147463
rect 120716 145951 121156 147377
rect 120716 145865 120809 145951
rect 120895 145865 120977 145951
rect 121063 145865 121156 145951
rect 120716 144439 121156 145865
rect 120716 144353 120809 144439
rect 120895 144353 120977 144439
rect 121063 144353 121156 144439
rect 120716 142927 121156 144353
rect 120716 142841 120809 142927
rect 120895 142841 120977 142927
rect 121063 142841 121156 142927
rect 120716 141415 121156 142841
rect 120716 141329 120809 141415
rect 120895 141329 120977 141415
rect 121063 141329 121156 141415
rect 120716 139903 121156 141329
rect 120716 139817 120809 139903
rect 120895 139817 120977 139903
rect 121063 139817 121156 139903
rect 120716 138391 121156 139817
rect 120716 138305 120809 138391
rect 120895 138305 120977 138391
rect 121063 138305 121156 138391
rect 120716 136879 121156 138305
rect 120716 136793 120809 136879
rect 120895 136793 120977 136879
rect 121063 136793 121156 136879
rect 120716 136450 121156 136793
rect 120716 136070 120746 136450
rect 121126 136070 121156 136450
rect 120716 135367 121156 136070
rect 120716 135281 120809 135367
rect 120895 135281 120977 135367
rect 121063 135281 121156 135367
rect 120716 133855 121156 135281
rect 120716 133769 120809 133855
rect 120895 133769 120977 133855
rect 121063 133769 121156 133855
rect 120716 132343 121156 133769
rect 120716 132257 120809 132343
rect 120895 132257 120977 132343
rect 121063 132257 121156 132343
rect 120716 130831 121156 132257
rect 120716 130745 120809 130831
rect 120895 130745 120977 130831
rect 121063 130745 121156 130831
rect 120716 129319 121156 130745
rect 120716 129233 120809 129319
rect 120895 129233 120977 129319
rect 121063 129233 121156 129319
rect 120716 127807 121156 129233
rect 120716 127721 120809 127807
rect 120895 127721 120977 127807
rect 121063 127721 121156 127807
rect 120716 126295 121156 127721
rect 120716 126209 120809 126295
rect 120895 126209 120977 126295
rect 121063 126209 121156 126295
rect 120716 124783 121156 126209
rect 120716 124697 120809 124783
rect 120895 124697 120977 124783
rect 121063 124697 121156 124783
rect 120716 123271 121156 124697
rect 120716 123185 120809 123271
rect 120895 123185 120977 123271
rect 121063 123185 121156 123271
rect 120716 121759 121156 123185
rect 120716 121673 120809 121759
rect 120895 121673 120977 121759
rect 121063 121673 121156 121759
rect 120716 121330 121156 121673
rect 120716 120950 120746 121330
rect 121126 120950 121156 121330
rect 120716 120247 121156 120950
rect 120716 120161 120809 120247
rect 120895 120161 120977 120247
rect 121063 120161 121156 120247
rect 120716 118735 121156 120161
rect 120716 118649 120809 118735
rect 120895 118649 120977 118735
rect 121063 118649 121156 118735
rect 120716 117223 121156 118649
rect 120716 117137 120809 117223
rect 120895 117137 120977 117223
rect 121063 117137 121156 117223
rect 120716 115711 121156 117137
rect 120716 115625 120809 115711
rect 120895 115625 120977 115711
rect 121063 115625 121156 115711
rect 120716 114199 121156 115625
rect 120716 114113 120809 114199
rect 120895 114113 120977 114199
rect 121063 114113 121156 114199
rect 120716 112687 121156 114113
rect 120716 112601 120809 112687
rect 120895 112601 120977 112687
rect 121063 112601 121156 112687
rect 120716 111175 121156 112601
rect 120716 111089 120809 111175
rect 120895 111089 120977 111175
rect 121063 111089 121156 111175
rect 120716 109663 121156 111089
rect 120716 109577 120809 109663
rect 120895 109577 120977 109663
rect 121063 109577 121156 109663
rect 120716 108151 121156 109577
rect 120716 108065 120809 108151
rect 120895 108065 120977 108151
rect 121063 108065 121156 108151
rect 120716 106639 121156 108065
rect 120716 106553 120809 106639
rect 120895 106553 120977 106639
rect 121063 106553 121156 106639
rect 120716 106210 121156 106553
rect 120716 105830 120746 106210
rect 121126 105830 121156 106210
rect 120716 105127 121156 105830
rect 120716 105041 120809 105127
rect 120895 105041 120977 105127
rect 121063 105041 121156 105127
rect 120716 103615 121156 105041
rect 120716 103529 120809 103615
rect 120895 103529 120977 103615
rect 121063 103529 121156 103615
rect 120716 102103 121156 103529
rect 120716 102017 120809 102103
rect 120895 102017 120977 102103
rect 121063 102017 121156 102103
rect 120716 100591 121156 102017
rect 120716 100505 120809 100591
rect 120895 100505 120977 100591
rect 121063 100505 121156 100591
rect 120716 99079 121156 100505
rect 120716 98993 120809 99079
rect 120895 98993 120977 99079
rect 121063 98993 121156 99079
rect 120716 97567 121156 98993
rect 120716 97481 120809 97567
rect 120895 97481 120977 97567
rect 121063 97481 121156 97567
rect 120716 96055 121156 97481
rect 120716 95969 120809 96055
rect 120895 95969 120977 96055
rect 121063 95969 121156 96055
rect 120716 94543 121156 95969
rect 120716 94457 120809 94543
rect 120895 94457 120977 94543
rect 121063 94457 121156 94543
rect 120716 93031 121156 94457
rect 120716 92945 120809 93031
rect 120895 92945 120977 93031
rect 121063 92945 121156 93031
rect 120716 91519 121156 92945
rect 120716 91433 120809 91519
rect 120895 91433 120977 91519
rect 121063 91433 121156 91519
rect 120716 91090 121156 91433
rect 120716 90710 120746 91090
rect 121126 90710 121156 91090
rect 120716 90007 121156 90710
rect 120716 89921 120809 90007
rect 120895 89921 120977 90007
rect 121063 89921 121156 90007
rect 120716 88495 121156 89921
rect 120716 88409 120809 88495
rect 120895 88409 120977 88495
rect 121063 88409 121156 88495
rect 120716 86983 121156 88409
rect 120716 86897 120809 86983
rect 120895 86897 120977 86983
rect 121063 86897 121156 86983
rect 120716 85471 121156 86897
rect 120716 85385 120809 85471
rect 120895 85385 120977 85471
rect 121063 85385 121156 85471
rect 120716 83959 121156 85385
rect 120716 83873 120809 83959
rect 120895 83873 120977 83959
rect 121063 83873 121156 83959
rect 120716 82447 121156 83873
rect 120716 82361 120809 82447
rect 120895 82361 120977 82447
rect 121063 82361 121156 82447
rect 120716 80935 121156 82361
rect 120716 80849 120809 80935
rect 120895 80849 120977 80935
rect 121063 80849 121156 80935
rect 120716 79423 121156 80849
rect 120716 79337 120809 79423
rect 120895 79337 120977 79423
rect 121063 79337 121156 79423
rect 120716 77911 121156 79337
rect 120716 77825 120809 77911
rect 120895 77825 120977 77911
rect 121063 77825 121156 77911
rect 120716 76399 121156 77825
rect 120716 76313 120809 76399
rect 120895 76313 120977 76399
rect 121063 76313 121156 76399
rect 120716 75970 121156 76313
rect 120716 75590 120746 75970
rect 121126 75590 121156 75970
rect 120716 74887 121156 75590
rect 120716 74801 120809 74887
rect 120895 74801 120977 74887
rect 121063 74801 121156 74887
rect 120716 73375 121156 74801
rect 120716 73289 120809 73375
rect 120895 73289 120977 73375
rect 121063 73289 121156 73375
rect 120716 71863 121156 73289
rect 120716 71777 120809 71863
rect 120895 71777 120977 71863
rect 121063 71777 121156 71863
rect 120716 69406 121156 71777
rect 120716 69026 120746 69406
rect 121126 69026 121156 69406
rect 120716 69014 121156 69026
rect 120716 68634 120746 69014
rect 121126 68634 121156 69014
rect 120716 68520 121156 68634
rect 134596 153742 135036 155256
rect 134596 153362 134626 153742
rect 135006 153362 135036 153742
rect 134596 153350 135036 153362
rect 134596 152970 134626 153350
rect 135006 152970 135036 153350
rect 134596 151243 135036 152970
rect 134596 151157 134689 151243
rect 134775 151157 134857 151243
rect 134943 151157 135036 151243
rect 134596 150330 135036 151157
rect 134596 149950 134626 150330
rect 135006 149950 135036 150330
rect 134596 149731 135036 149950
rect 134596 149645 134689 149731
rect 134775 149645 134857 149731
rect 134943 149645 135036 149731
rect 134596 148219 135036 149645
rect 134596 148133 134689 148219
rect 134775 148133 134857 148219
rect 134943 148133 135036 148219
rect 134596 146707 135036 148133
rect 134596 146621 134689 146707
rect 134775 146621 134857 146707
rect 134943 146621 135036 146707
rect 134596 145195 135036 146621
rect 134596 145109 134689 145195
rect 134775 145109 134857 145195
rect 134943 145109 135036 145195
rect 134596 143683 135036 145109
rect 134596 143597 134689 143683
rect 134775 143597 134857 143683
rect 134943 143597 135036 143683
rect 134596 142171 135036 143597
rect 134596 142085 134689 142171
rect 134775 142085 134857 142171
rect 134943 142085 135036 142171
rect 134596 140659 135036 142085
rect 134596 140573 134689 140659
rect 134775 140573 134857 140659
rect 134943 140573 135036 140659
rect 134596 139147 135036 140573
rect 134596 139061 134689 139147
rect 134775 139061 134857 139147
rect 134943 139061 135036 139147
rect 134596 137635 135036 139061
rect 134596 137549 134689 137635
rect 134775 137549 134857 137635
rect 134943 137549 135036 137635
rect 134596 136123 135036 137549
rect 134596 136037 134689 136123
rect 134775 136037 134857 136123
rect 134943 136037 135036 136123
rect 134596 135210 135036 136037
rect 134596 134830 134626 135210
rect 135006 134830 135036 135210
rect 134596 134611 135036 134830
rect 134596 134525 134689 134611
rect 134775 134525 134857 134611
rect 134943 134525 135036 134611
rect 134596 133099 135036 134525
rect 134596 133013 134689 133099
rect 134775 133013 134857 133099
rect 134943 133013 135036 133099
rect 134596 131587 135036 133013
rect 134596 131501 134689 131587
rect 134775 131501 134857 131587
rect 134943 131501 135036 131587
rect 134596 130075 135036 131501
rect 134596 129989 134689 130075
rect 134775 129989 134857 130075
rect 134943 129989 135036 130075
rect 134596 128563 135036 129989
rect 134596 128477 134689 128563
rect 134775 128477 134857 128563
rect 134943 128477 135036 128563
rect 134596 127051 135036 128477
rect 134596 126965 134689 127051
rect 134775 126965 134857 127051
rect 134943 126965 135036 127051
rect 134596 125539 135036 126965
rect 134596 125453 134689 125539
rect 134775 125453 134857 125539
rect 134943 125453 135036 125539
rect 134596 124027 135036 125453
rect 134596 123941 134689 124027
rect 134775 123941 134857 124027
rect 134943 123941 135036 124027
rect 134596 122515 135036 123941
rect 134596 122429 134689 122515
rect 134775 122429 134857 122515
rect 134943 122429 135036 122515
rect 134596 121003 135036 122429
rect 134596 120917 134689 121003
rect 134775 120917 134857 121003
rect 134943 120917 135036 121003
rect 134596 120090 135036 120917
rect 134596 119710 134626 120090
rect 135006 119710 135036 120090
rect 134596 119491 135036 119710
rect 134596 119405 134689 119491
rect 134775 119405 134857 119491
rect 134943 119405 135036 119491
rect 134596 117979 135036 119405
rect 134596 117893 134689 117979
rect 134775 117893 134857 117979
rect 134943 117893 135036 117979
rect 134596 116467 135036 117893
rect 134596 116381 134689 116467
rect 134775 116381 134857 116467
rect 134943 116381 135036 116467
rect 134596 114955 135036 116381
rect 134596 114869 134689 114955
rect 134775 114869 134857 114955
rect 134943 114869 135036 114955
rect 134596 113443 135036 114869
rect 134596 113357 134689 113443
rect 134775 113357 134857 113443
rect 134943 113357 135036 113443
rect 134596 111931 135036 113357
rect 134596 111845 134689 111931
rect 134775 111845 134857 111931
rect 134943 111845 135036 111931
rect 134596 110419 135036 111845
rect 134596 110333 134689 110419
rect 134775 110333 134857 110419
rect 134943 110333 135036 110419
rect 134596 108907 135036 110333
rect 134596 108821 134689 108907
rect 134775 108821 134857 108907
rect 134943 108821 135036 108907
rect 134596 107395 135036 108821
rect 134596 107309 134689 107395
rect 134775 107309 134857 107395
rect 134943 107309 135036 107395
rect 134596 105883 135036 107309
rect 134596 105797 134689 105883
rect 134775 105797 134857 105883
rect 134943 105797 135036 105883
rect 134596 104970 135036 105797
rect 134596 104590 134626 104970
rect 135006 104590 135036 104970
rect 134596 104371 135036 104590
rect 134596 104285 134689 104371
rect 134775 104285 134857 104371
rect 134943 104285 135036 104371
rect 134596 102859 135036 104285
rect 134596 102773 134689 102859
rect 134775 102773 134857 102859
rect 134943 102773 135036 102859
rect 134596 101347 135036 102773
rect 134596 101261 134689 101347
rect 134775 101261 134857 101347
rect 134943 101261 135036 101347
rect 134596 99835 135036 101261
rect 134596 99749 134689 99835
rect 134775 99749 134857 99835
rect 134943 99749 135036 99835
rect 134596 98323 135036 99749
rect 134596 98237 134689 98323
rect 134775 98237 134857 98323
rect 134943 98237 135036 98323
rect 134596 96811 135036 98237
rect 134596 96725 134689 96811
rect 134775 96725 134857 96811
rect 134943 96725 135036 96811
rect 134596 95299 135036 96725
rect 134596 95213 134689 95299
rect 134775 95213 134857 95299
rect 134943 95213 135036 95299
rect 134596 93787 135036 95213
rect 134596 93701 134689 93787
rect 134775 93701 134857 93787
rect 134943 93701 135036 93787
rect 134596 92275 135036 93701
rect 134596 92189 134689 92275
rect 134775 92189 134857 92275
rect 134943 92189 135036 92275
rect 134596 90763 135036 92189
rect 134596 90677 134689 90763
rect 134775 90677 134857 90763
rect 134943 90677 135036 90763
rect 134596 89850 135036 90677
rect 134596 89470 134626 89850
rect 135006 89470 135036 89850
rect 134596 89251 135036 89470
rect 134596 89165 134689 89251
rect 134775 89165 134857 89251
rect 134943 89165 135036 89251
rect 134596 87739 135036 89165
rect 134596 87653 134689 87739
rect 134775 87653 134857 87739
rect 134943 87653 135036 87739
rect 134596 86227 135036 87653
rect 134596 86141 134689 86227
rect 134775 86141 134857 86227
rect 134943 86141 135036 86227
rect 134596 84715 135036 86141
rect 134596 84629 134689 84715
rect 134775 84629 134857 84715
rect 134943 84629 135036 84715
rect 134596 83203 135036 84629
rect 134596 83117 134689 83203
rect 134775 83117 134857 83203
rect 134943 83117 135036 83203
rect 134596 81691 135036 83117
rect 134596 81605 134689 81691
rect 134775 81605 134857 81691
rect 134943 81605 135036 81691
rect 134596 80179 135036 81605
rect 134596 80093 134689 80179
rect 134775 80093 134857 80179
rect 134943 80093 135036 80179
rect 134596 78667 135036 80093
rect 134596 78581 134689 78667
rect 134775 78581 134857 78667
rect 134943 78581 135036 78667
rect 134596 77155 135036 78581
rect 134596 77069 134689 77155
rect 134775 77069 134857 77155
rect 134943 77069 135036 77155
rect 134596 75643 135036 77069
rect 134596 75557 134689 75643
rect 134775 75557 134857 75643
rect 134943 75557 135036 75643
rect 134596 74730 135036 75557
rect 134596 74350 134626 74730
rect 135006 74350 135036 74730
rect 134596 74131 135036 74350
rect 134596 74045 134689 74131
rect 134775 74045 134857 74131
rect 134943 74045 135036 74131
rect 134596 72619 135036 74045
rect 134596 72533 134689 72619
rect 134775 72533 134857 72619
rect 134943 72533 135036 72619
rect 134596 70806 135036 72533
rect 134596 70426 134626 70806
rect 135006 70426 135036 70806
rect 134596 70414 135036 70426
rect 134596 70034 134626 70414
rect 135006 70034 135036 70414
rect 134596 68520 135036 70034
rect 135836 155142 136276 155256
rect 135836 154762 135866 155142
rect 136246 154762 136276 155142
rect 135836 154750 136276 154762
rect 135836 154370 135866 154750
rect 136246 154370 136276 154750
rect 135836 151999 136276 154370
rect 135836 151913 135929 151999
rect 136015 151913 136097 151999
rect 136183 151913 136276 151999
rect 135836 151570 136276 151913
rect 135836 151190 135866 151570
rect 136246 151190 136276 151570
rect 135836 150487 136276 151190
rect 135836 150401 135929 150487
rect 136015 150401 136097 150487
rect 136183 150401 136276 150487
rect 135836 148975 136276 150401
rect 135836 148889 135929 148975
rect 136015 148889 136097 148975
rect 136183 148889 136276 148975
rect 135836 147463 136276 148889
rect 135836 147377 135929 147463
rect 136015 147377 136097 147463
rect 136183 147377 136276 147463
rect 135836 145951 136276 147377
rect 135836 145865 135929 145951
rect 136015 145865 136097 145951
rect 136183 145865 136276 145951
rect 135836 144439 136276 145865
rect 135836 144353 135929 144439
rect 136015 144353 136097 144439
rect 136183 144353 136276 144439
rect 135836 142927 136276 144353
rect 135836 142841 135929 142927
rect 136015 142841 136097 142927
rect 136183 142841 136276 142927
rect 135836 141415 136276 142841
rect 135836 141329 135929 141415
rect 136015 141329 136097 141415
rect 136183 141329 136276 141415
rect 135836 139903 136276 141329
rect 135836 139817 135929 139903
rect 136015 139817 136097 139903
rect 136183 139817 136276 139903
rect 135836 138391 136276 139817
rect 135836 138305 135929 138391
rect 136015 138305 136097 138391
rect 136183 138305 136276 138391
rect 135836 136879 136276 138305
rect 135836 136793 135929 136879
rect 136015 136793 136097 136879
rect 136183 136793 136276 136879
rect 135836 136450 136276 136793
rect 135836 136070 135866 136450
rect 136246 136070 136276 136450
rect 135836 135367 136276 136070
rect 135836 135281 135929 135367
rect 136015 135281 136097 135367
rect 136183 135281 136276 135367
rect 135836 133855 136276 135281
rect 135836 133769 135929 133855
rect 136015 133769 136097 133855
rect 136183 133769 136276 133855
rect 135836 132343 136276 133769
rect 135836 132257 135929 132343
rect 136015 132257 136097 132343
rect 136183 132257 136276 132343
rect 135836 130831 136276 132257
rect 135836 130745 135929 130831
rect 136015 130745 136097 130831
rect 136183 130745 136276 130831
rect 135836 129319 136276 130745
rect 135836 129233 135929 129319
rect 136015 129233 136097 129319
rect 136183 129233 136276 129319
rect 135836 127807 136276 129233
rect 135836 127721 135929 127807
rect 136015 127721 136097 127807
rect 136183 127721 136276 127807
rect 135836 126295 136276 127721
rect 135836 126209 135929 126295
rect 136015 126209 136097 126295
rect 136183 126209 136276 126295
rect 135836 124783 136276 126209
rect 135836 124697 135929 124783
rect 136015 124697 136097 124783
rect 136183 124697 136276 124783
rect 135836 123271 136276 124697
rect 135836 123185 135929 123271
rect 136015 123185 136097 123271
rect 136183 123185 136276 123271
rect 135836 121759 136276 123185
rect 135836 121673 135929 121759
rect 136015 121673 136097 121759
rect 136183 121673 136276 121759
rect 135836 121330 136276 121673
rect 135836 120950 135866 121330
rect 136246 120950 136276 121330
rect 135836 120247 136276 120950
rect 135836 120161 135929 120247
rect 136015 120161 136097 120247
rect 136183 120161 136276 120247
rect 135836 118735 136276 120161
rect 135836 118649 135929 118735
rect 136015 118649 136097 118735
rect 136183 118649 136276 118735
rect 135836 117223 136276 118649
rect 135836 117137 135929 117223
rect 136015 117137 136097 117223
rect 136183 117137 136276 117223
rect 135836 115711 136276 117137
rect 135836 115625 135929 115711
rect 136015 115625 136097 115711
rect 136183 115625 136276 115711
rect 135836 114199 136276 115625
rect 135836 114113 135929 114199
rect 136015 114113 136097 114199
rect 136183 114113 136276 114199
rect 135836 112687 136276 114113
rect 135836 112601 135929 112687
rect 136015 112601 136097 112687
rect 136183 112601 136276 112687
rect 135836 111175 136276 112601
rect 135836 111089 135929 111175
rect 136015 111089 136097 111175
rect 136183 111089 136276 111175
rect 135836 109663 136276 111089
rect 135836 109577 135929 109663
rect 136015 109577 136097 109663
rect 136183 109577 136276 109663
rect 135836 108151 136276 109577
rect 135836 108065 135929 108151
rect 136015 108065 136097 108151
rect 136183 108065 136276 108151
rect 135836 106639 136276 108065
rect 135836 106553 135929 106639
rect 136015 106553 136097 106639
rect 136183 106553 136276 106639
rect 135836 106210 136276 106553
rect 135836 105830 135866 106210
rect 136246 105830 136276 106210
rect 135836 105127 136276 105830
rect 135836 105041 135929 105127
rect 136015 105041 136097 105127
rect 136183 105041 136276 105127
rect 135836 103615 136276 105041
rect 135836 103529 135929 103615
rect 136015 103529 136097 103615
rect 136183 103529 136276 103615
rect 135836 102103 136276 103529
rect 135836 102017 135929 102103
rect 136015 102017 136097 102103
rect 136183 102017 136276 102103
rect 135836 100591 136276 102017
rect 135836 100505 135929 100591
rect 136015 100505 136097 100591
rect 136183 100505 136276 100591
rect 135836 99079 136276 100505
rect 135836 98993 135929 99079
rect 136015 98993 136097 99079
rect 136183 98993 136276 99079
rect 135836 97567 136276 98993
rect 135836 97481 135929 97567
rect 136015 97481 136097 97567
rect 136183 97481 136276 97567
rect 135836 96055 136276 97481
rect 135836 95969 135929 96055
rect 136015 95969 136097 96055
rect 136183 95969 136276 96055
rect 135836 94543 136276 95969
rect 135836 94457 135929 94543
rect 136015 94457 136097 94543
rect 136183 94457 136276 94543
rect 135836 93031 136276 94457
rect 135836 92945 135929 93031
rect 136015 92945 136097 93031
rect 136183 92945 136276 93031
rect 135836 91519 136276 92945
rect 135836 91433 135929 91519
rect 136015 91433 136097 91519
rect 136183 91433 136276 91519
rect 135836 91090 136276 91433
rect 135836 90710 135866 91090
rect 136246 90710 136276 91090
rect 135836 90007 136276 90710
rect 135836 89921 135929 90007
rect 136015 89921 136097 90007
rect 136183 89921 136276 90007
rect 135836 88495 136276 89921
rect 135836 88409 135929 88495
rect 136015 88409 136097 88495
rect 136183 88409 136276 88495
rect 135836 86983 136276 88409
rect 135836 86897 135929 86983
rect 136015 86897 136097 86983
rect 136183 86897 136276 86983
rect 135836 85471 136276 86897
rect 135836 85385 135929 85471
rect 136015 85385 136097 85471
rect 136183 85385 136276 85471
rect 135836 83959 136276 85385
rect 135836 83873 135929 83959
rect 136015 83873 136097 83959
rect 136183 83873 136276 83959
rect 135836 82447 136276 83873
rect 135836 82361 135929 82447
rect 136015 82361 136097 82447
rect 136183 82361 136276 82447
rect 135836 80935 136276 82361
rect 135836 80849 135929 80935
rect 136015 80849 136097 80935
rect 136183 80849 136276 80935
rect 135836 79423 136276 80849
rect 135836 79337 135929 79423
rect 136015 79337 136097 79423
rect 136183 79337 136276 79423
rect 135836 77911 136276 79337
rect 135836 77825 135929 77911
rect 136015 77825 136097 77911
rect 136183 77825 136276 77911
rect 135836 76399 136276 77825
rect 135836 76313 135929 76399
rect 136015 76313 136097 76399
rect 136183 76313 136276 76399
rect 135836 75970 136276 76313
rect 135836 75590 135866 75970
rect 136246 75590 136276 75970
rect 135836 74887 136276 75590
rect 135836 74801 135929 74887
rect 136015 74801 136097 74887
rect 136183 74801 136276 74887
rect 135836 73375 136276 74801
rect 135836 73289 135929 73375
rect 136015 73289 136097 73375
rect 136183 73289 136276 73375
rect 135836 71863 136276 73289
rect 135836 71777 135929 71863
rect 136015 71777 136097 71863
rect 136183 71777 136276 71863
rect 135836 69406 136276 71777
rect 135836 69026 135866 69406
rect 136246 69026 136276 69406
rect 135836 69014 136276 69026
rect 135836 68634 135866 69014
rect 136246 68634 136276 69014
rect 135836 68520 136276 68634
rect 149716 153742 150156 155256
rect 149716 153362 149746 153742
rect 150126 153362 150156 153742
rect 149716 153350 150156 153362
rect 149716 152970 149746 153350
rect 150126 152970 150156 153350
rect 149716 151243 150156 152970
rect 149716 151157 149809 151243
rect 149895 151157 149977 151243
rect 150063 151157 150156 151243
rect 149716 150330 150156 151157
rect 149716 149950 149746 150330
rect 150126 149950 150156 150330
rect 149716 149731 150156 149950
rect 149716 149645 149809 149731
rect 149895 149645 149977 149731
rect 150063 149645 150156 149731
rect 149716 148219 150156 149645
rect 149716 148133 149809 148219
rect 149895 148133 149977 148219
rect 150063 148133 150156 148219
rect 149716 146707 150156 148133
rect 149716 146621 149809 146707
rect 149895 146621 149977 146707
rect 150063 146621 150156 146707
rect 149716 145195 150156 146621
rect 149716 145109 149809 145195
rect 149895 145109 149977 145195
rect 150063 145109 150156 145195
rect 149716 143683 150156 145109
rect 149716 143597 149809 143683
rect 149895 143597 149977 143683
rect 150063 143597 150156 143683
rect 149716 142171 150156 143597
rect 149716 142085 149809 142171
rect 149895 142085 149977 142171
rect 150063 142085 150156 142171
rect 149716 140659 150156 142085
rect 149716 140573 149809 140659
rect 149895 140573 149977 140659
rect 150063 140573 150156 140659
rect 149716 139147 150156 140573
rect 149716 139061 149809 139147
rect 149895 139061 149977 139147
rect 150063 139061 150156 139147
rect 149716 137635 150156 139061
rect 149716 137549 149809 137635
rect 149895 137549 149977 137635
rect 150063 137549 150156 137635
rect 149716 136123 150156 137549
rect 149716 136037 149809 136123
rect 149895 136037 149977 136123
rect 150063 136037 150156 136123
rect 149716 135210 150156 136037
rect 149716 134830 149746 135210
rect 150126 134830 150156 135210
rect 149716 134611 150156 134830
rect 149716 134525 149809 134611
rect 149895 134525 149977 134611
rect 150063 134525 150156 134611
rect 149716 133099 150156 134525
rect 149716 133013 149809 133099
rect 149895 133013 149977 133099
rect 150063 133013 150156 133099
rect 149716 131587 150156 133013
rect 149716 131501 149809 131587
rect 149895 131501 149977 131587
rect 150063 131501 150156 131587
rect 149716 130075 150156 131501
rect 149716 129989 149809 130075
rect 149895 129989 149977 130075
rect 150063 129989 150156 130075
rect 149716 128563 150156 129989
rect 149716 128477 149809 128563
rect 149895 128477 149977 128563
rect 150063 128477 150156 128563
rect 149716 127051 150156 128477
rect 149716 126965 149809 127051
rect 149895 126965 149977 127051
rect 150063 126965 150156 127051
rect 149716 125539 150156 126965
rect 149716 125453 149809 125539
rect 149895 125453 149977 125539
rect 150063 125453 150156 125539
rect 149716 124027 150156 125453
rect 149716 123941 149809 124027
rect 149895 123941 149977 124027
rect 150063 123941 150156 124027
rect 149716 122515 150156 123941
rect 149716 122429 149809 122515
rect 149895 122429 149977 122515
rect 150063 122429 150156 122515
rect 149716 121003 150156 122429
rect 149716 120917 149809 121003
rect 149895 120917 149977 121003
rect 150063 120917 150156 121003
rect 149716 120090 150156 120917
rect 149716 119710 149746 120090
rect 150126 119710 150156 120090
rect 149716 119491 150156 119710
rect 149716 119405 149809 119491
rect 149895 119405 149977 119491
rect 150063 119405 150156 119491
rect 149716 117979 150156 119405
rect 149716 117893 149809 117979
rect 149895 117893 149977 117979
rect 150063 117893 150156 117979
rect 149716 116467 150156 117893
rect 149716 116381 149809 116467
rect 149895 116381 149977 116467
rect 150063 116381 150156 116467
rect 149716 114955 150156 116381
rect 149716 114869 149809 114955
rect 149895 114869 149977 114955
rect 150063 114869 150156 114955
rect 149716 113443 150156 114869
rect 149716 113357 149809 113443
rect 149895 113357 149977 113443
rect 150063 113357 150156 113443
rect 149716 111931 150156 113357
rect 149716 111845 149809 111931
rect 149895 111845 149977 111931
rect 150063 111845 150156 111931
rect 149716 110419 150156 111845
rect 149716 110333 149809 110419
rect 149895 110333 149977 110419
rect 150063 110333 150156 110419
rect 149716 108907 150156 110333
rect 149716 108821 149809 108907
rect 149895 108821 149977 108907
rect 150063 108821 150156 108907
rect 149716 107395 150156 108821
rect 149716 107309 149809 107395
rect 149895 107309 149977 107395
rect 150063 107309 150156 107395
rect 149716 105883 150156 107309
rect 149716 105797 149809 105883
rect 149895 105797 149977 105883
rect 150063 105797 150156 105883
rect 149716 104970 150156 105797
rect 149716 104590 149746 104970
rect 150126 104590 150156 104970
rect 149716 104371 150156 104590
rect 149716 104285 149809 104371
rect 149895 104285 149977 104371
rect 150063 104285 150156 104371
rect 149716 102859 150156 104285
rect 149716 102773 149809 102859
rect 149895 102773 149977 102859
rect 150063 102773 150156 102859
rect 149716 101347 150156 102773
rect 149716 101261 149809 101347
rect 149895 101261 149977 101347
rect 150063 101261 150156 101347
rect 149716 99835 150156 101261
rect 149716 99749 149809 99835
rect 149895 99749 149977 99835
rect 150063 99749 150156 99835
rect 149716 98323 150156 99749
rect 149716 98237 149809 98323
rect 149895 98237 149977 98323
rect 150063 98237 150156 98323
rect 149716 96811 150156 98237
rect 149716 96725 149809 96811
rect 149895 96725 149977 96811
rect 150063 96725 150156 96811
rect 149716 95299 150156 96725
rect 149716 95213 149809 95299
rect 149895 95213 149977 95299
rect 150063 95213 150156 95299
rect 149716 93787 150156 95213
rect 149716 93701 149809 93787
rect 149895 93701 149977 93787
rect 150063 93701 150156 93787
rect 149716 92275 150156 93701
rect 149716 92189 149809 92275
rect 149895 92189 149977 92275
rect 150063 92189 150156 92275
rect 149716 90763 150156 92189
rect 149716 90677 149809 90763
rect 149895 90677 149977 90763
rect 150063 90677 150156 90763
rect 149716 89850 150156 90677
rect 149716 89470 149746 89850
rect 150126 89470 150156 89850
rect 149716 89251 150156 89470
rect 149716 89165 149809 89251
rect 149895 89165 149977 89251
rect 150063 89165 150156 89251
rect 149716 87739 150156 89165
rect 149716 87653 149809 87739
rect 149895 87653 149977 87739
rect 150063 87653 150156 87739
rect 149716 86227 150156 87653
rect 149716 86141 149809 86227
rect 149895 86141 149977 86227
rect 150063 86141 150156 86227
rect 149716 84715 150156 86141
rect 149716 84629 149809 84715
rect 149895 84629 149977 84715
rect 150063 84629 150156 84715
rect 149716 83203 150156 84629
rect 149716 83117 149809 83203
rect 149895 83117 149977 83203
rect 150063 83117 150156 83203
rect 149716 81691 150156 83117
rect 149716 81605 149809 81691
rect 149895 81605 149977 81691
rect 150063 81605 150156 81691
rect 149716 80179 150156 81605
rect 149716 80093 149809 80179
rect 149895 80093 149977 80179
rect 150063 80093 150156 80179
rect 149716 78667 150156 80093
rect 149716 78581 149809 78667
rect 149895 78581 149977 78667
rect 150063 78581 150156 78667
rect 149716 77155 150156 78581
rect 149716 77069 149809 77155
rect 149895 77069 149977 77155
rect 150063 77069 150156 77155
rect 149716 75643 150156 77069
rect 149716 75557 149809 75643
rect 149895 75557 149977 75643
rect 150063 75557 150156 75643
rect 149716 74730 150156 75557
rect 149716 74350 149746 74730
rect 150126 74350 150156 74730
rect 149716 74131 150156 74350
rect 149716 74045 149809 74131
rect 149895 74045 149977 74131
rect 150063 74045 150156 74131
rect 149716 72619 150156 74045
rect 149716 72533 149809 72619
rect 149895 72533 149977 72619
rect 150063 72533 150156 72619
rect 149716 70806 150156 72533
rect 149716 70426 149746 70806
rect 150126 70426 150156 70806
rect 149716 70414 150156 70426
rect 149716 70034 149746 70414
rect 150126 70034 150156 70414
rect 149716 68520 150156 70034
rect 150956 155142 151396 155256
rect 150956 154762 150986 155142
rect 151366 154762 151396 155142
rect 150956 154750 151396 154762
rect 150956 154370 150986 154750
rect 151366 154370 151396 154750
rect 150956 151999 151396 154370
rect 154652 155142 155652 155256
rect 154652 154762 154766 155142
rect 155146 154762 155158 155142
rect 155538 154762 155652 155142
rect 154652 154750 155652 154762
rect 154652 154370 154766 154750
rect 155146 154370 155158 154750
rect 155538 154370 155652 154750
rect 150956 151913 151049 151999
rect 151135 151913 151217 151999
rect 151303 151913 151396 151999
rect 150956 151570 151396 151913
rect 150956 151190 150986 151570
rect 151366 151190 151396 151570
rect 150956 150487 151396 151190
rect 150956 150401 151049 150487
rect 151135 150401 151217 150487
rect 151303 150401 151396 150487
rect 150956 148975 151396 150401
rect 150956 148889 151049 148975
rect 151135 148889 151217 148975
rect 151303 148889 151396 148975
rect 150956 147463 151396 148889
rect 150956 147377 151049 147463
rect 151135 147377 151217 147463
rect 151303 147377 151396 147463
rect 150956 145951 151396 147377
rect 150956 145865 151049 145951
rect 151135 145865 151217 145951
rect 151303 145865 151396 145951
rect 150956 144439 151396 145865
rect 150956 144353 151049 144439
rect 151135 144353 151217 144439
rect 151303 144353 151396 144439
rect 150956 142927 151396 144353
rect 150956 142841 151049 142927
rect 151135 142841 151217 142927
rect 151303 142841 151396 142927
rect 150956 141415 151396 142841
rect 150956 141329 151049 141415
rect 151135 141329 151217 141415
rect 151303 141329 151396 141415
rect 150956 139903 151396 141329
rect 150956 139817 151049 139903
rect 151135 139817 151217 139903
rect 151303 139817 151396 139903
rect 150956 138391 151396 139817
rect 150956 138305 151049 138391
rect 151135 138305 151217 138391
rect 151303 138305 151396 138391
rect 150956 136879 151396 138305
rect 150956 136793 151049 136879
rect 151135 136793 151217 136879
rect 151303 136793 151396 136879
rect 150956 136450 151396 136793
rect 150956 136070 150986 136450
rect 151366 136070 151396 136450
rect 150956 135367 151396 136070
rect 150956 135281 151049 135367
rect 151135 135281 151217 135367
rect 151303 135281 151396 135367
rect 150956 133855 151396 135281
rect 150956 133769 151049 133855
rect 151135 133769 151217 133855
rect 151303 133769 151396 133855
rect 150956 132343 151396 133769
rect 150956 132257 151049 132343
rect 151135 132257 151217 132343
rect 151303 132257 151396 132343
rect 150956 130831 151396 132257
rect 150956 130745 151049 130831
rect 151135 130745 151217 130831
rect 151303 130745 151396 130831
rect 150956 129319 151396 130745
rect 150956 129233 151049 129319
rect 151135 129233 151217 129319
rect 151303 129233 151396 129319
rect 150956 127807 151396 129233
rect 150956 127721 151049 127807
rect 151135 127721 151217 127807
rect 151303 127721 151396 127807
rect 150956 126295 151396 127721
rect 150956 126209 151049 126295
rect 151135 126209 151217 126295
rect 151303 126209 151396 126295
rect 150956 124783 151396 126209
rect 150956 124697 151049 124783
rect 151135 124697 151217 124783
rect 151303 124697 151396 124783
rect 150956 123271 151396 124697
rect 150956 123185 151049 123271
rect 151135 123185 151217 123271
rect 151303 123185 151396 123271
rect 150956 121759 151396 123185
rect 150956 121673 151049 121759
rect 151135 121673 151217 121759
rect 151303 121673 151396 121759
rect 150956 121330 151396 121673
rect 150956 120950 150986 121330
rect 151366 120950 151396 121330
rect 150956 120247 151396 120950
rect 150956 120161 151049 120247
rect 151135 120161 151217 120247
rect 151303 120161 151396 120247
rect 150956 118735 151396 120161
rect 150956 118649 151049 118735
rect 151135 118649 151217 118735
rect 151303 118649 151396 118735
rect 150956 117223 151396 118649
rect 150956 117137 151049 117223
rect 151135 117137 151217 117223
rect 151303 117137 151396 117223
rect 150956 115711 151396 117137
rect 150956 115625 151049 115711
rect 151135 115625 151217 115711
rect 151303 115625 151396 115711
rect 150956 114199 151396 115625
rect 150956 114113 151049 114199
rect 151135 114113 151217 114199
rect 151303 114113 151396 114199
rect 150956 112687 151396 114113
rect 150956 112601 151049 112687
rect 151135 112601 151217 112687
rect 151303 112601 151396 112687
rect 150956 111175 151396 112601
rect 150956 111089 151049 111175
rect 151135 111089 151217 111175
rect 151303 111089 151396 111175
rect 150956 109663 151396 111089
rect 150956 109577 151049 109663
rect 151135 109577 151217 109663
rect 151303 109577 151396 109663
rect 150956 108151 151396 109577
rect 150956 108065 151049 108151
rect 151135 108065 151217 108151
rect 151303 108065 151396 108151
rect 150956 106639 151396 108065
rect 150956 106553 151049 106639
rect 151135 106553 151217 106639
rect 151303 106553 151396 106639
rect 150956 106210 151396 106553
rect 150956 105830 150986 106210
rect 151366 105830 151396 106210
rect 150956 105127 151396 105830
rect 150956 105041 151049 105127
rect 151135 105041 151217 105127
rect 151303 105041 151396 105127
rect 150956 103615 151396 105041
rect 150956 103529 151049 103615
rect 151135 103529 151217 103615
rect 151303 103529 151396 103615
rect 150956 102103 151396 103529
rect 150956 102017 151049 102103
rect 151135 102017 151217 102103
rect 151303 102017 151396 102103
rect 150956 100591 151396 102017
rect 150956 100505 151049 100591
rect 151135 100505 151217 100591
rect 151303 100505 151396 100591
rect 150956 99079 151396 100505
rect 150956 98993 151049 99079
rect 151135 98993 151217 99079
rect 151303 98993 151396 99079
rect 150956 97567 151396 98993
rect 150956 97481 151049 97567
rect 151135 97481 151217 97567
rect 151303 97481 151396 97567
rect 150956 96055 151396 97481
rect 150956 95969 151049 96055
rect 151135 95969 151217 96055
rect 151303 95969 151396 96055
rect 150956 94543 151396 95969
rect 150956 94457 151049 94543
rect 151135 94457 151217 94543
rect 151303 94457 151396 94543
rect 150956 93031 151396 94457
rect 150956 92945 151049 93031
rect 151135 92945 151217 93031
rect 151303 92945 151396 93031
rect 150956 91519 151396 92945
rect 150956 91433 151049 91519
rect 151135 91433 151217 91519
rect 151303 91433 151396 91519
rect 150956 91090 151396 91433
rect 150956 90710 150986 91090
rect 151366 90710 151396 91090
rect 150956 90007 151396 90710
rect 150956 89921 151049 90007
rect 151135 89921 151217 90007
rect 151303 89921 151396 90007
rect 150956 88495 151396 89921
rect 150956 88409 151049 88495
rect 151135 88409 151217 88495
rect 151303 88409 151396 88495
rect 150956 86983 151396 88409
rect 150956 86897 151049 86983
rect 151135 86897 151217 86983
rect 151303 86897 151396 86983
rect 150956 85471 151396 86897
rect 150956 85385 151049 85471
rect 151135 85385 151217 85471
rect 151303 85385 151396 85471
rect 150956 83959 151396 85385
rect 150956 83873 151049 83959
rect 151135 83873 151217 83959
rect 151303 83873 151396 83959
rect 150956 82447 151396 83873
rect 150956 82361 151049 82447
rect 151135 82361 151217 82447
rect 151303 82361 151396 82447
rect 150956 80935 151396 82361
rect 150956 80849 151049 80935
rect 151135 80849 151217 80935
rect 151303 80849 151396 80935
rect 150956 79423 151396 80849
rect 150956 79337 151049 79423
rect 151135 79337 151217 79423
rect 151303 79337 151396 79423
rect 150956 77911 151396 79337
rect 150956 77825 151049 77911
rect 151135 77825 151217 77911
rect 151303 77825 151396 77911
rect 150956 76399 151396 77825
rect 150956 76313 151049 76399
rect 151135 76313 151217 76399
rect 151303 76313 151396 76399
rect 150956 75970 151396 76313
rect 150956 75590 150986 75970
rect 151366 75590 151396 75970
rect 150956 74887 151396 75590
rect 150956 74801 151049 74887
rect 151135 74801 151217 74887
rect 151303 74801 151396 74887
rect 150956 73375 151396 74801
rect 150956 73289 151049 73375
rect 151135 73289 151217 73375
rect 151303 73289 151396 73375
rect 150956 71863 151396 73289
rect 150956 71777 151049 71863
rect 151135 71777 151217 71863
rect 151303 71777 151396 71863
rect 150956 69406 151396 71777
rect 153252 153742 154252 153856
rect 153252 153362 153366 153742
rect 153746 153362 153758 153742
rect 154138 153362 154252 153742
rect 153252 153350 154252 153362
rect 153252 152970 153366 153350
rect 153746 152970 153758 153350
rect 154138 152970 154252 153350
rect 153252 149169 154252 152970
rect 153252 148789 153366 149169
rect 153746 148789 153758 149169
rect 154138 148789 154252 149169
rect 153252 148777 154252 148789
rect 153252 148397 153366 148777
rect 153746 148397 153758 148777
rect 154138 148397 154252 148777
rect 153252 148385 154252 148397
rect 153252 148005 153366 148385
rect 153746 148005 153758 148385
rect 154138 148005 154252 148385
rect 153252 147993 154252 148005
rect 153252 147613 153366 147993
rect 153746 147613 153758 147993
rect 154138 147613 154252 147993
rect 153252 147601 154252 147613
rect 153252 147221 153366 147601
rect 153746 147221 153758 147601
rect 154138 147221 154252 147601
rect 153252 147209 154252 147221
rect 153252 146829 153366 147209
rect 153746 146829 153758 147209
rect 154138 146829 154252 147209
rect 153252 135210 154252 146829
rect 153252 134830 153366 135210
rect 153746 134830 153758 135210
rect 154138 134830 154252 135210
rect 153252 133169 154252 134830
rect 153252 132789 153366 133169
rect 153746 132789 153758 133169
rect 154138 132789 154252 133169
rect 153252 132777 154252 132789
rect 153252 132397 153366 132777
rect 153746 132397 153758 132777
rect 154138 132397 154252 132777
rect 153252 132385 154252 132397
rect 153252 132005 153366 132385
rect 153746 132005 153758 132385
rect 154138 132005 154252 132385
rect 153252 131993 154252 132005
rect 153252 131613 153366 131993
rect 153746 131613 153758 131993
rect 154138 131613 154252 131993
rect 153252 131601 154252 131613
rect 153252 131221 153366 131601
rect 153746 131221 153758 131601
rect 154138 131221 154252 131601
rect 153252 131209 154252 131221
rect 153252 130829 153366 131209
rect 153746 130829 153758 131209
rect 154138 130829 154252 131209
rect 153252 120090 154252 130829
rect 153252 119710 153366 120090
rect 153746 119710 153758 120090
rect 154138 119710 154252 120090
rect 153252 117169 154252 119710
rect 153252 116789 153366 117169
rect 153746 116789 153758 117169
rect 154138 116789 154252 117169
rect 153252 116777 154252 116789
rect 153252 116397 153366 116777
rect 153746 116397 153758 116777
rect 154138 116397 154252 116777
rect 153252 116385 154252 116397
rect 153252 116005 153366 116385
rect 153746 116005 153758 116385
rect 154138 116005 154252 116385
rect 153252 115993 154252 116005
rect 153252 115613 153366 115993
rect 153746 115613 153758 115993
rect 154138 115613 154252 115993
rect 153252 115601 154252 115613
rect 153252 115221 153366 115601
rect 153746 115221 153758 115601
rect 154138 115221 154252 115601
rect 153252 115209 154252 115221
rect 153252 114829 153366 115209
rect 153746 114829 153758 115209
rect 154138 114829 154252 115209
rect 153252 104970 154252 114829
rect 153252 104590 153366 104970
rect 153746 104590 153758 104970
rect 154138 104590 154252 104970
rect 153252 101169 154252 104590
rect 153252 100789 153366 101169
rect 153746 100789 153758 101169
rect 154138 100789 154252 101169
rect 153252 100777 154252 100789
rect 153252 100397 153366 100777
rect 153746 100397 153758 100777
rect 154138 100397 154252 100777
rect 153252 100385 154252 100397
rect 153252 100005 153366 100385
rect 153746 100005 153758 100385
rect 154138 100005 154252 100385
rect 153252 99993 154252 100005
rect 153252 99613 153366 99993
rect 153746 99613 153758 99993
rect 154138 99613 154252 99993
rect 153252 99601 154252 99613
rect 153252 99221 153366 99601
rect 153746 99221 153758 99601
rect 154138 99221 154252 99601
rect 153252 99209 154252 99221
rect 153252 98829 153366 99209
rect 153746 98829 153758 99209
rect 154138 98829 154252 99209
rect 153252 89850 154252 98829
rect 153252 89470 153366 89850
rect 153746 89470 153758 89850
rect 154138 89470 154252 89850
rect 153252 85169 154252 89470
rect 153252 84789 153366 85169
rect 153746 84789 153758 85169
rect 154138 84789 154252 85169
rect 153252 84777 154252 84789
rect 153252 84397 153366 84777
rect 153746 84397 153758 84777
rect 154138 84397 154252 84777
rect 153252 84385 154252 84397
rect 153252 84005 153366 84385
rect 153746 84005 153758 84385
rect 154138 84005 154252 84385
rect 153252 83993 154252 84005
rect 153252 83613 153366 83993
rect 153746 83613 153758 83993
rect 154138 83613 154252 83993
rect 153252 83601 154252 83613
rect 153252 83221 153366 83601
rect 153746 83221 153758 83601
rect 154138 83221 154252 83601
rect 153252 83209 154252 83221
rect 153252 82829 153366 83209
rect 153746 82829 153758 83209
rect 154138 82829 154252 83209
rect 153252 74730 154252 82829
rect 153252 74350 153366 74730
rect 153746 74350 153758 74730
rect 154138 74350 154252 74730
rect 153252 70806 154252 74350
rect 153252 70426 153366 70806
rect 153746 70426 153758 70806
rect 154138 70426 154252 70806
rect 153252 70414 154252 70426
rect 153252 70034 153366 70414
rect 153746 70034 153758 70414
rect 154138 70034 154252 70414
rect 153252 69920 154252 70034
rect 154652 151570 155652 154370
rect 160400 154501 164000 154664
rect 160400 154121 160442 154501
rect 160822 154121 160834 154501
rect 161214 154121 161226 154501
rect 161606 154121 161618 154501
rect 161998 154121 162010 154501
rect 162390 154121 162402 154501
rect 162782 154121 162794 154501
rect 163174 154121 163186 154501
rect 163566 154121 163578 154501
rect 163958 154121 164000 154501
rect 160400 154109 164000 154121
rect 160400 153729 160442 154109
rect 160822 153729 160834 154109
rect 161214 153729 161226 154109
rect 161606 153729 161618 154109
rect 161998 153729 162010 154109
rect 162390 153729 162402 154109
rect 162782 153729 162794 154109
rect 163174 153729 163186 154109
rect 163566 153729 163578 154109
rect 163958 153729 164000 154109
rect 160400 153717 164000 153729
rect 160400 153337 160442 153717
rect 160822 153337 160834 153717
rect 161214 153337 161226 153717
rect 161606 153337 161618 153717
rect 161998 153337 162010 153717
rect 162390 153337 162402 153717
rect 162782 153337 162794 153717
rect 163174 153337 163186 153717
rect 163566 153337 163578 153717
rect 163958 153337 164000 153717
rect 160400 153325 164000 153337
rect 160400 152945 160442 153325
rect 160822 152945 160834 153325
rect 161214 152945 161226 153325
rect 161606 152945 161618 153325
rect 161998 152945 162010 153325
rect 162390 152945 162402 153325
rect 162782 152945 162794 153325
rect 163174 152945 163186 153325
rect 163566 152945 163578 153325
rect 163958 152945 164000 153325
rect 160400 152933 164000 152945
rect 160400 152553 160442 152933
rect 160822 152553 160834 152933
rect 161214 152553 161226 152933
rect 161606 152553 161618 152933
rect 161998 152553 162010 152933
rect 162390 152553 162402 152933
rect 162782 152553 162794 152933
rect 163174 152553 163186 152933
rect 163566 152553 163578 152933
rect 163958 152553 164000 152933
rect 160400 152541 164000 152553
rect 160400 152161 160442 152541
rect 160822 152161 160834 152541
rect 161214 152161 161226 152541
rect 161606 152161 161618 152541
rect 161998 152161 162010 152541
rect 162390 152161 162402 152541
rect 162782 152161 162794 152541
rect 163174 152161 163186 152541
rect 163566 152161 163578 152541
rect 163958 152161 164000 152541
rect 160400 151998 164000 152161
rect 154652 151190 154766 151570
rect 155146 151190 155158 151570
rect 155538 151190 155652 151570
rect 154652 138501 155652 151190
rect 164400 149169 168000 149332
rect 164400 148789 164442 149169
rect 164822 148789 164834 149169
rect 165214 148789 165226 149169
rect 165606 148789 165618 149169
rect 165998 148789 166010 149169
rect 166390 148789 166402 149169
rect 166782 148789 166794 149169
rect 167174 148789 167186 149169
rect 167566 148789 167578 149169
rect 167958 148789 168000 149169
rect 164400 148777 168000 148789
rect 164400 148397 164442 148777
rect 164822 148397 164834 148777
rect 165214 148397 165226 148777
rect 165606 148397 165618 148777
rect 165998 148397 166010 148777
rect 166390 148397 166402 148777
rect 166782 148397 166794 148777
rect 167174 148397 167186 148777
rect 167566 148397 167578 148777
rect 167958 148397 168000 148777
rect 164400 148385 168000 148397
rect 164400 148005 164442 148385
rect 164822 148005 164834 148385
rect 165214 148005 165226 148385
rect 165606 148005 165618 148385
rect 165998 148005 166010 148385
rect 166390 148005 166402 148385
rect 166782 148005 166794 148385
rect 167174 148005 167186 148385
rect 167566 148005 167578 148385
rect 167958 148005 168000 148385
rect 164400 147993 168000 148005
rect 164400 147613 164442 147993
rect 164822 147613 164834 147993
rect 165214 147613 165226 147993
rect 165606 147613 165618 147993
rect 165998 147613 166010 147993
rect 166390 147613 166402 147993
rect 166782 147613 166794 147993
rect 167174 147613 167186 147993
rect 167566 147613 167578 147993
rect 167958 147613 168000 147993
rect 164400 147601 168000 147613
rect 164400 147221 164442 147601
rect 164822 147221 164834 147601
rect 165214 147221 165226 147601
rect 165606 147221 165618 147601
rect 165998 147221 166010 147601
rect 166390 147221 166402 147601
rect 166782 147221 166794 147601
rect 167174 147221 167186 147601
rect 167566 147221 167578 147601
rect 167958 147221 168000 147601
rect 164400 147209 168000 147221
rect 164400 146829 164442 147209
rect 164822 146829 164834 147209
rect 165214 146829 165226 147209
rect 165606 146829 165618 147209
rect 165998 146829 166010 147209
rect 166390 146829 166402 147209
rect 166782 146829 166794 147209
rect 167174 146829 167186 147209
rect 167566 146829 167578 147209
rect 167958 146829 168000 147209
rect 164400 146666 168000 146829
rect 154652 138121 154766 138501
rect 155146 138121 155158 138501
rect 155538 138121 155652 138501
rect 154652 138109 155652 138121
rect 154652 137729 154766 138109
rect 155146 137729 155158 138109
rect 155538 137729 155652 138109
rect 154652 137717 155652 137729
rect 154652 137337 154766 137717
rect 155146 137337 155158 137717
rect 155538 137337 155652 137717
rect 154652 137325 155652 137337
rect 154652 136945 154766 137325
rect 155146 136945 155158 137325
rect 155538 136945 155652 137325
rect 154652 136933 155652 136945
rect 154652 136553 154766 136933
rect 155146 136553 155158 136933
rect 155538 136553 155652 136933
rect 154652 136541 155652 136553
rect 154652 136161 154766 136541
rect 155146 136161 155158 136541
rect 155538 136161 155652 136541
rect 154652 122501 155652 136161
rect 160400 138501 164000 138664
rect 160400 138121 160442 138501
rect 160822 138121 160834 138501
rect 161214 138121 161226 138501
rect 161606 138121 161618 138501
rect 161998 138121 162010 138501
rect 162390 138121 162402 138501
rect 162782 138121 162794 138501
rect 163174 138121 163186 138501
rect 163566 138121 163578 138501
rect 163958 138121 164000 138501
rect 160400 138109 164000 138121
rect 160400 137729 160442 138109
rect 160822 137729 160834 138109
rect 161214 137729 161226 138109
rect 161606 137729 161618 138109
rect 161998 137729 162010 138109
rect 162390 137729 162402 138109
rect 162782 137729 162794 138109
rect 163174 137729 163186 138109
rect 163566 137729 163578 138109
rect 163958 137729 164000 138109
rect 160400 137717 164000 137729
rect 160400 137337 160442 137717
rect 160822 137337 160834 137717
rect 161214 137337 161226 137717
rect 161606 137337 161618 137717
rect 161998 137337 162010 137717
rect 162390 137337 162402 137717
rect 162782 137337 162794 137717
rect 163174 137337 163186 137717
rect 163566 137337 163578 137717
rect 163958 137337 164000 137717
rect 160400 137325 164000 137337
rect 160400 136945 160442 137325
rect 160822 136945 160834 137325
rect 161214 136945 161226 137325
rect 161606 136945 161618 137325
rect 161998 136945 162010 137325
rect 162390 136945 162402 137325
rect 162782 136945 162794 137325
rect 163174 136945 163186 137325
rect 163566 136945 163578 137325
rect 163958 136945 164000 137325
rect 160400 136933 164000 136945
rect 160400 136553 160442 136933
rect 160822 136553 160834 136933
rect 161214 136553 161226 136933
rect 161606 136553 161618 136933
rect 161998 136553 162010 136933
rect 162390 136553 162402 136933
rect 162782 136553 162794 136933
rect 163174 136553 163186 136933
rect 163566 136553 163578 136933
rect 163958 136553 164000 136933
rect 160400 136541 164000 136553
rect 160400 136161 160442 136541
rect 160822 136161 160834 136541
rect 161214 136161 161226 136541
rect 161606 136161 161618 136541
rect 161998 136161 162010 136541
rect 162390 136161 162402 136541
rect 162782 136161 162794 136541
rect 163174 136161 163186 136541
rect 163566 136161 163578 136541
rect 163958 136161 164000 136541
rect 160400 135998 164000 136161
rect 164400 133169 168000 133332
rect 164400 132789 164442 133169
rect 164822 132789 164834 133169
rect 165214 132789 165226 133169
rect 165606 132789 165618 133169
rect 165998 132789 166010 133169
rect 166390 132789 166402 133169
rect 166782 132789 166794 133169
rect 167174 132789 167186 133169
rect 167566 132789 167578 133169
rect 167958 132789 168000 133169
rect 164400 132777 168000 132789
rect 164400 132397 164442 132777
rect 164822 132397 164834 132777
rect 165214 132397 165226 132777
rect 165606 132397 165618 132777
rect 165998 132397 166010 132777
rect 166390 132397 166402 132777
rect 166782 132397 166794 132777
rect 167174 132397 167186 132777
rect 167566 132397 167578 132777
rect 167958 132397 168000 132777
rect 164400 132385 168000 132397
rect 164400 132005 164442 132385
rect 164822 132005 164834 132385
rect 165214 132005 165226 132385
rect 165606 132005 165618 132385
rect 165998 132005 166010 132385
rect 166390 132005 166402 132385
rect 166782 132005 166794 132385
rect 167174 132005 167186 132385
rect 167566 132005 167578 132385
rect 167958 132005 168000 132385
rect 164400 131993 168000 132005
rect 164400 131613 164442 131993
rect 164822 131613 164834 131993
rect 165214 131613 165226 131993
rect 165606 131613 165618 131993
rect 165998 131613 166010 131993
rect 166390 131613 166402 131993
rect 166782 131613 166794 131993
rect 167174 131613 167186 131993
rect 167566 131613 167578 131993
rect 167958 131613 168000 131993
rect 164400 131601 168000 131613
rect 164400 131221 164442 131601
rect 164822 131221 164834 131601
rect 165214 131221 165226 131601
rect 165606 131221 165618 131601
rect 165998 131221 166010 131601
rect 166390 131221 166402 131601
rect 166782 131221 166794 131601
rect 167174 131221 167186 131601
rect 167566 131221 167578 131601
rect 167958 131221 168000 131601
rect 164400 131209 168000 131221
rect 164400 130829 164442 131209
rect 164822 130829 164834 131209
rect 165214 130829 165226 131209
rect 165606 130829 165618 131209
rect 165998 130829 166010 131209
rect 166390 130829 166402 131209
rect 166782 130829 166794 131209
rect 167174 130829 167186 131209
rect 167566 130829 167578 131209
rect 167958 130829 168000 131209
rect 164400 130666 168000 130829
rect 154652 122121 154766 122501
rect 155146 122121 155158 122501
rect 155538 122121 155652 122501
rect 154652 122109 155652 122121
rect 154652 121729 154766 122109
rect 155146 121729 155158 122109
rect 155538 121729 155652 122109
rect 154652 121717 155652 121729
rect 154652 121337 154766 121717
rect 155146 121337 155158 121717
rect 155538 121337 155652 121717
rect 154652 121325 155652 121337
rect 154652 120945 154766 121325
rect 155146 120945 155158 121325
rect 155538 120945 155652 121325
rect 154652 120933 155652 120945
rect 154652 120553 154766 120933
rect 155146 120553 155158 120933
rect 155538 120553 155652 120933
rect 154652 120541 155652 120553
rect 154652 120161 154766 120541
rect 155146 120161 155158 120541
rect 155538 120161 155652 120541
rect 154652 106501 155652 120161
rect 160400 122501 164000 122664
rect 160400 122121 160442 122501
rect 160822 122121 160834 122501
rect 161214 122121 161226 122501
rect 161606 122121 161618 122501
rect 161998 122121 162010 122501
rect 162390 122121 162402 122501
rect 162782 122121 162794 122501
rect 163174 122121 163186 122501
rect 163566 122121 163578 122501
rect 163958 122121 164000 122501
rect 160400 122109 164000 122121
rect 160400 121729 160442 122109
rect 160822 121729 160834 122109
rect 161214 121729 161226 122109
rect 161606 121729 161618 122109
rect 161998 121729 162010 122109
rect 162390 121729 162402 122109
rect 162782 121729 162794 122109
rect 163174 121729 163186 122109
rect 163566 121729 163578 122109
rect 163958 121729 164000 122109
rect 160400 121717 164000 121729
rect 160400 121337 160442 121717
rect 160822 121337 160834 121717
rect 161214 121337 161226 121717
rect 161606 121337 161618 121717
rect 161998 121337 162010 121717
rect 162390 121337 162402 121717
rect 162782 121337 162794 121717
rect 163174 121337 163186 121717
rect 163566 121337 163578 121717
rect 163958 121337 164000 121717
rect 160400 121325 164000 121337
rect 160400 120945 160442 121325
rect 160822 120945 160834 121325
rect 161214 120945 161226 121325
rect 161606 120945 161618 121325
rect 161998 120945 162010 121325
rect 162390 120945 162402 121325
rect 162782 120945 162794 121325
rect 163174 120945 163186 121325
rect 163566 120945 163578 121325
rect 163958 120945 164000 121325
rect 160400 120933 164000 120945
rect 160400 120553 160442 120933
rect 160822 120553 160834 120933
rect 161214 120553 161226 120933
rect 161606 120553 161618 120933
rect 161998 120553 162010 120933
rect 162390 120553 162402 120933
rect 162782 120553 162794 120933
rect 163174 120553 163186 120933
rect 163566 120553 163578 120933
rect 163958 120553 164000 120933
rect 160400 120541 164000 120553
rect 160400 120161 160442 120541
rect 160822 120161 160834 120541
rect 161214 120161 161226 120541
rect 161606 120161 161618 120541
rect 161998 120161 162010 120541
rect 162390 120161 162402 120541
rect 162782 120161 162794 120541
rect 163174 120161 163186 120541
rect 163566 120161 163578 120541
rect 163958 120161 164000 120541
rect 160400 119998 164000 120161
rect 164400 117169 168000 117332
rect 164400 116789 164442 117169
rect 164822 116789 164834 117169
rect 165214 116789 165226 117169
rect 165606 116789 165618 117169
rect 165998 116789 166010 117169
rect 166390 116789 166402 117169
rect 166782 116789 166794 117169
rect 167174 116789 167186 117169
rect 167566 116789 167578 117169
rect 167958 116789 168000 117169
rect 164400 116777 168000 116789
rect 164400 116397 164442 116777
rect 164822 116397 164834 116777
rect 165214 116397 165226 116777
rect 165606 116397 165618 116777
rect 165998 116397 166010 116777
rect 166390 116397 166402 116777
rect 166782 116397 166794 116777
rect 167174 116397 167186 116777
rect 167566 116397 167578 116777
rect 167958 116397 168000 116777
rect 164400 116385 168000 116397
rect 164400 116005 164442 116385
rect 164822 116005 164834 116385
rect 165214 116005 165226 116385
rect 165606 116005 165618 116385
rect 165998 116005 166010 116385
rect 166390 116005 166402 116385
rect 166782 116005 166794 116385
rect 167174 116005 167186 116385
rect 167566 116005 167578 116385
rect 167958 116005 168000 116385
rect 164400 115993 168000 116005
rect 164400 115613 164442 115993
rect 164822 115613 164834 115993
rect 165214 115613 165226 115993
rect 165606 115613 165618 115993
rect 165998 115613 166010 115993
rect 166390 115613 166402 115993
rect 166782 115613 166794 115993
rect 167174 115613 167186 115993
rect 167566 115613 167578 115993
rect 167958 115613 168000 115993
rect 164400 115601 168000 115613
rect 164400 115221 164442 115601
rect 164822 115221 164834 115601
rect 165214 115221 165226 115601
rect 165606 115221 165618 115601
rect 165998 115221 166010 115601
rect 166390 115221 166402 115601
rect 166782 115221 166794 115601
rect 167174 115221 167186 115601
rect 167566 115221 167578 115601
rect 167958 115221 168000 115601
rect 164400 115209 168000 115221
rect 164400 114829 164442 115209
rect 164822 114829 164834 115209
rect 165214 114829 165226 115209
rect 165606 114829 165618 115209
rect 165998 114829 166010 115209
rect 166390 114829 166402 115209
rect 166782 114829 166794 115209
rect 167174 114829 167186 115209
rect 167566 114829 167578 115209
rect 167958 114829 168000 115209
rect 164400 114666 168000 114829
rect 154652 106121 154766 106501
rect 155146 106121 155158 106501
rect 155538 106121 155652 106501
rect 154652 106109 155652 106121
rect 154652 105729 154766 106109
rect 155146 105729 155158 106109
rect 155538 105729 155652 106109
rect 154652 105717 155652 105729
rect 154652 105337 154766 105717
rect 155146 105337 155158 105717
rect 155538 105337 155652 105717
rect 154652 105325 155652 105337
rect 154652 104945 154766 105325
rect 155146 104945 155158 105325
rect 155538 104945 155652 105325
rect 154652 104933 155652 104945
rect 154652 104553 154766 104933
rect 155146 104553 155158 104933
rect 155538 104553 155652 104933
rect 154652 104541 155652 104553
rect 154652 104161 154766 104541
rect 155146 104161 155158 104541
rect 155538 104161 155652 104541
rect 154652 90501 155652 104161
rect 160400 106501 164000 106664
rect 160400 106121 160442 106501
rect 160822 106121 160834 106501
rect 161214 106121 161226 106501
rect 161606 106121 161618 106501
rect 161998 106121 162010 106501
rect 162390 106121 162402 106501
rect 162782 106121 162794 106501
rect 163174 106121 163186 106501
rect 163566 106121 163578 106501
rect 163958 106121 164000 106501
rect 160400 106109 164000 106121
rect 160400 105729 160442 106109
rect 160822 105729 160834 106109
rect 161214 105729 161226 106109
rect 161606 105729 161618 106109
rect 161998 105729 162010 106109
rect 162390 105729 162402 106109
rect 162782 105729 162794 106109
rect 163174 105729 163186 106109
rect 163566 105729 163578 106109
rect 163958 105729 164000 106109
rect 160400 105717 164000 105729
rect 160400 105337 160442 105717
rect 160822 105337 160834 105717
rect 161214 105337 161226 105717
rect 161606 105337 161618 105717
rect 161998 105337 162010 105717
rect 162390 105337 162402 105717
rect 162782 105337 162794 105717
rect 163174 105337 163186 105717
rect 163566 105337 163578 105717
rect 163958 105337 164000 105717
rect 160400 105325 164000 105337
rect 160400 104945 160442 105325
rect 160822 104945 160834 105325
rect 161214 104945 161226 105325
rect 161606 104945 161618 105325
rect 161998 104945 162010 105325
rect 162390 104945 162402 105325
rect 162782 104945 162794 105325
rect 163174 104945 163186 105325
rect 163566 104945 163578 105325
rect 163958 104945 164000 105325
rect 160400 104933 164000 104945
rect 160400 104553 160442 104933
rect 160822 104553 160834 104933
rect 161214 104553 161226 104933
rect 161606 104553 161618 104933
rect 161998 104553 162010 104933
rect 162390 104553 162402 104933
rect 162782 104553 162794 104933
rect 163174 104553 163186 104933
rect 163566 104553 163578 104933
rect 163958 104553 164000 104933
rect 160400 104541 164000 104553
rect 160400 104161 160442 104541
rect 160822 104161 160834 104541
rect 161214 104161 161226 104541
rect 161606 104161 161618 104541
rect 161998 104161 162010 104541
rect 162390 104161 162402 104541
rect 162782 104161 162794 104541
rect 163174 104161 163186 104541
rect 163566 104161 163578 104541
rect 163958 104161 164000 104541
rect 160400 103998 164000 104161
rect 164400 101169 168000 101332
rect 164400 100789 164442 101169
rect 164822 100789 164834 101169
rect 165214 100789 165226 101169
rect 165606 100789 165618 101169
rect 165998 100789 166010 101169
rect 166390 100789 166402 101169
rect 166782 100789 166794 101169
rect 167174 100789 167186 101169
rect 167566 100789 167578 101169
rect 167958 100789 168000 101169
rect 164400 100777 168000 100789
rect 164400 100397 164442 100777
rect 164822 100397 164834 100777
rect 165214 100397 165226 100777
rect 165606 100397 165618 100777
rect 165998 100397 166010 100777
rect 166390 100397 166402 100777
rect 166782 100397 166794 100777
rect 167174 100397 167186 100777
rect 167566 100397 167578 100777
rect 167958 100397 168000 100777
rect 164400 100385 168000 100397
rect 164400 100005 164442 100385
rect 164822 100005 164834 100385
rect 165214 100005 165226 100385
rect 165606 100005 165618 100385
rect 165998 100005 166010 100385
rect 166390 100005 166402 100385
rect 166782 100005 166794 100385
rect 167174 100005 167186 100385
rect 167566 100005 167578 100385
rect 167958 100005 168000 100385
rect 164400 99993 168000 100005
rect 164400 99613 164442 99993
rect 164822 99613 164834 99993
rect 165214 99613 165226 99993
rect 165606 99613 165618 99993
rect 165998 99613 166010 99993
rect 166390 99613 166402 99993
rect 166782 99613 166794 99993
rect 167174 99613 167186 99993
rect 167566 99613 167578 99993
rect 167958 99613 168000 99993
rect 164400 99601 168000 99613
rect 164400 99221 164442 99601
rect 164822 99221 164834 99601
rect 165214 99221 165226 99601
rect 165606 99221 165618 99601
rect 165998 99221 166010 99601
rect 166390 99221 166402 99601
rect 166782 99221 166794 99601
rect 167174 99221 167186 99601
rect 167566 99221 167578 99601
rect 167958 99221 168000 99601
rect 164400 99209 168000 99221
rect 164400 98829 164442 99209
rect 164822 98829 164834 99209
rect 165214 98829 165226 99209
rect 165606 98829 165618 99209
rect 165998 98829 166010 99209
rect 166390 98829 166402 99209
rect 166782 98829 166794 99209
rect 167174 98829 167186 99209
rect 167566 98829 167578 99209
rect 167958 98829 168000 99209
rect 164400 98666 168000 98829
rect 154652 90121 154766 90501
rect 155146 90121 155158 90501
rect 155538 90121 155652 90501
rect 154652 90109 155652 90121
rect 154652 89729 154766 90109
rect 155146 89729 155158 90109
rect 155538 89729 155652 90109
rect 154652 89717 155652 89729
rect 154652 89337 154766 89717
rect 155146 89337 155158 89717
rect 155538 89337 155652 89717
rect 154652 89325 155652 89337
rect 154652 88945 154766 89325
rect 155146 88945 155158 89325
rect 155538 88945 155652 89325
rect 154652 88933 155652 88945
rect 154652 88553 154766 88933
rect 155146 88553 155158 88933
rect 155538 88553 155652 88933
rect 154652 88541 155652 88553
rect 154652 88161 154766 88541
rect 155146 88161 155158 88541
rect 155538 88161 155652 88541
rect 154652 75970 155652 88161
rect 160400 90501 164000 90664
rect 160400 90121 160442 90501
rect 160822 90121 160834 90501
rect 161214 90121 161226 90501
rect 161606 90121 161618 90501
rect 161998 90121 162010 90501
rect 162390 90121 162402 90501
rect 162782 90121 162794 90501
rect 163174 90121 163186 90501
rect 163566 90121 163578 90501
rect 163958 90121 164000 90501
rect 160400 90109 164000 90121
rect 160400 89729 160442 90109
rect 160822 89729 160834 90109
rect 161214 89729 161226 90109
rect 161606 89729 161618 90109
rect 161998 89729 162010 90109
rect 162390 89729 162402 90109
rect 162782 89729 162794 90109
rect 163174 89729 163186 90109
rect 163566 89729 163578 90109
rect 163958 89729 164000 90109
rect 160400 89717 164000 89729
rect 160400 89337 160442 89717
rect 160822 89337 160834 89717
rect 161214 89337 161226 89717
rect 161606 89337 161618 89717
rect 161998 89337 162010 89717
rect 162390 89337 162402 89717
rect 162782 89337 162794 89717
rect 163174 89337 163186 89717
rect 163566 89337 163578 89717
rect 163958 89337 164000 89717
rect 160400 89325 164000 89337
rect 160400 88945 160442 89325
rect 160822 88945 160834 89325
rect 161214 88945 161226 89325
rect 161606 88945 161618 89325
rect 161998 88945 162010 89325
rect 162390 88945 162402 89325
rect 162782 88945 162794 89325
rect 163174 88945 163186 89325
rect 163566 88945 163578 89325
rect 163958 88945 164000 89325
rect 160400 88933 164000 88945
rect 160400 88553 160442 88933
rect 160822 88553 160834 88933
rect 161214 88553 161226 88933
rect 161606 88553 161618 88933
rect 161998 88553 162010 88933
rect 162390 88553 162402 88933
rect 162782 88553 162794 88933
rect 163174 88553 163186 88933
rect 163566 88553 163578 88933
rect 163958 88553 164000 88933
rect 160400 88541 164000 88553
rect 160400 88161 160442 88541
rect 160822 88161 160834 88541
rect 161214 88161 161226 88541
rect 161606 88161 161618 88541
rect 161998 88161 162010 88541
rect 162390 88161 162402 88541
rect 162782 88161 162794 88541
rect 163174 88161 163186 88541
rect 163566 88161 163578 88541
rect 163958 88161 164000 88541
rect 160400 87998 164000 88161
rect 164400 85169 168000 85332
rect 164400 84789 164442 85169
rect 164822 84789 164834 85169
rect 165214 84789 165226 85169
rect 165606 84789 165618 85169
rect 165998 84789 166010 85169
rect 166390 84789 166402 85169
rect 166782 84789 166794 85169
rect 167174 84789 167186 85169
rect 167566 84789 167578 85169
rect 167958 84789 168000 85169
rect 164400 84777 168000 84789
rect 164400 84397 164442 84777
rect 164822 84397 164834 84777
rect 165214 84397 165226 84777
rect 165606 84397 165618 84777
rect 165998 84397 166010 84777
rect 166390 84397 166402 84777
rect 166782 84397 166794 84777
rect 167174 84397 167186 84777
rect 167566 84397 167578 84777
rect 167958 84397 168000 84777
rect 164400 84385 168000 84397
rect 164400 84005 164442 84385
rect 164822 84005 164834 84385
rect 165214 84005 165226 84385
rect 165606 84005 165618 84385
rect 165998 84005 166010 84385
rect 166390 84005 166402 84385
rect 166782 84005 166794 84385
rect 167174 84005 167186 84385
rect 167566 84005 167578 84385
rect 167958 84005 168000 84385
rect 164400 83993 168000 84005
rect 164400 83613 164442 83993
rect 164822 83613 164834 83993
rect 165214 83613 165226 83993
rect 165606 83613 165618 83993
rect 165998 83613 166010 83993
rect 166390 83613 166402 83993
rect 166782 83613 166794 83993
rect 167174 83613 167186 83993
rect 167566 83613 167578 83993
rect 167958 83613 168000 83993
rect 164400 83601 168000 83613
rect 164400 83221 164442 83601
rect 164822 83221 164834 83601
rect 165214 83221 165226 83601
rect 165606 83221 165618 83601
rect 165998 83221 166010 83601
rect 166390 83221 166402 83601
rect 166782 83221 166794 83601
rect 167174 83221 167186 83601
rect 167566 83221 167578 83601
rect 167958 83221 168000 83601
rect 164400 83209 168000 83221
rect 164400 82829 164442 83209
rect 164822 82829 164834 83209
rect 165214 82829 165226 83209
rect 165606 82829 165618 83209
rect 165998 82829 166010 83209
rect 166390 82829 166402 83209
rect 166782 82829 166794 83209
rect 167174 82829 167186 83209
rect 167566 82829 167578 83209
rect 167958 82829 168000 83209
rect 164400 82666 168000 82829
rect 154652 75590 154766 75970
rect 155146 75590 155158 75970
rect 155538 75590 155652 75970
rect 154652 74501 155652 75590
rect 154652 74121 154766 74501
rect 155146 74121 155158 74501
rect 155538 74121 155652 74501
rect 154652 74109 155652 74121
rect 154652 73729 154766 74109
rect 155146 73729 155158 74109
rect 155538 73729 155652 74109
rect 154652 73717 155652 73729
rect 154652 73337 154766 73717
rect 155146 73337 155158 73717
rect 155538 73337 155652 73717
rect 154652 73325 155652 73337
rect 154652 72945 154766 73325
rect 155146 72945 155158 73325
rect 155538 72945 155652 73325
rect 154652 72933 155652 72945
rect 154652 72553 154766 72933
rect 155146 72553 155158 72933
rect 155538 72553 155652 72933
rect 154652 72541 155652 72553
rect 154652 72161 154766 72541
rect 155146 72161 155158 72541
rect 155538 72161 155652 72541
rect 150956 69026 150986 69406
rect 151366 69026 151396 69406
rect 150956 69014 151396 69026
rect 150956 68634 150986 69014
rect 151366 68634 151396 69014
rect 150956 68520 151396 68634
rect 154652 69406 155652 72161
rect 160400 74501 164000 74664
rect 160400 74121 160442 74501
rect 160822 74121 160834 74501
rect 161214 74121 161226 74501
rect 161606 74121 161618 74501
rect 161998 74121 162010 74501
rect 162390 74121 162402 74501
rect 162782 74121 162794 74501
rect 163174 74121 163186 74501
rect 163566 74121 163578 74501
rect 163958 74121 164000 74501
rect 160400 74109 164000 74121
rect 160400 73729 160442 74109
rect 160822 73729 160834 74109
rect 161214 73729 161226 74109
rect 161606 73729 161618 74109
rect 161998 73729 162010 74109
rect 162390 73729 162402 74109
rect 162782 73729 162794 74109
rect 163174 73729 163186 74109
rect 163566 73729 163578 74109
rect 163958 73729 164000 74109
rect 160400 73717 164000 73729
rect 160400 73337 160442 73717
rect 160822 73337 160834 73717
rect 161214 73337 161226 73717
rect 161606 73337 161618 73717
rect 161998 73337 162010 73717
rect 162390 73337 162402 73717
rect 162782 73337 162794 73717
rect 163174 73337 163186 73717
rect 163566 73337 163578 73717
rect 163958 73337 164000 73717
rect 160400 73325 164000 73337
rect 160400 72945 160442 73325
rect 160822 72945 160834 73325
rect 161214 72945 161226 73325
rect 161606 72945 161618 73325
rect 161998 72945 162010 73325
rect 162390 72945 162402 73325
rect 162782 72945 162794 73325
rect 163174 72945 163186 73325
rect 163566 72945 163578 73325
rect 163958 72945 164000 73325
rect 160400 72933 164000 72945
rect 160400 72553 160442 72933
rect 160822 72553 160834 72933
rect 161214 72553 161226 72933
rect 161606 72553 161618 72933
rect 161998 72553 162010 72933
rect 162390 72553 162402 72933
rect 162782 72553 162794 72933
rect 163174 72553 163186 72933
rect 163566 72553 163578 72933
rect 163958 72553 164000 72933
rect 160400 72541 164000 72553
rect 160400 72161 160442 72541
rect 160822 72161 160834 72541
rect 161214 72161 161226 72541
rect 161606 72161 161618 72541
rect 161998 72161 162010 72541
rect 162390 72161 162402 72541
rect 162782 72161 162794 72541
rect 163174 72161 163186 72541
rect 163566 72161 163578 72541
rect 163958 72161 164000 72541
rect 160400 71998 164000 72161
rect 154652 69026 154766 69406
rect 155146 69026 155158 69406
rect 155538 69026 155652 69406
rect 154652 69014 155652 69026
rect 154652 68634 154766 69014
rect 155146 68634 155158 69014
rect 155538 68634 155652 69014
rect 154652 68520 155652 68634
rect 71998 63558 74664 63600
rect 71998 63178 72161 63558
rect 72541 63178 72553 63558
rect 72933 63178 72945 63558
rect 73325 63178 73337 63558
rect 73717 63178 73729 63558
rect 74109 63178 74121 63558
rect 74501 63178 74664 63558
rect 71998 63166 74664 63178
rect 71998 62786 72161 63166
rect 72541 62786 72553 63166
rect 72933 62786 72945 63166
rect 73325 62786 73337 63166
rect 73717 62786 73729 63166
rect 74109 62786 74121 63166
rect 74501 62786 74664 63166
rect 71998 62774 74664 62786
rect 71998 62394 72161 62774
rect 72541 62394 72553 62774
rect 72933 62394 72945 62774
rect 73325 62394 73337 62774
rect 73717 62394 73729 62774
rect 74109 62394 74121 62774
rect 74501 62394 74664 62774
rect 71998 62382 74664 62394
rect 71998 62002 72161 62382
rect 72541 62002 72553 62382
rect 72933 62002 72945 62382
rect 73325 62002 73337 62382
rect 73717 62002 73729 62382
rect 74109 62002 74121 62382
rect 74501 62002 74664 62382
rect 71998 61990 74664 62002
rect 71998 61610 72161 61990
rect 72541 61610 72553 61990
rect 72933 61610 72945 61990
rect 73325 61610 73337 61990
rect 73717 61610 73729 61990
rect 74109 61610 74121 61990
rect 74501 61610 74664 61990
rect 71998 61598 74664 61610
rect 71998 61218 72161 61598
rect 72541 61218 72553 61598
rect 72933 61218 72945 61598
rect 73325 61218 73337 61598
rect 73717 61218 73729 61598
rect 74109 61218 74121 61598
rect 74501 61218 74664 61598
rect 71998 61206 74664 61218
rect 71998 60826 72161 61206
rect 72541 60826 72553 61206
rect 72933 60826 72945 61206
rect 73325 60826 73337 61206
rect 73717 60826 73729 61206
rect 74109 60826 74121 61206
rect 74501 60826 74664 61206
rect 71998 60814 74664 60826
rect 71998 60434 72161 60814
rect 72541 60434 72553 60814
rect 72933 60434 72945 60814
rect 73325 60434 73337 60814
rect 73717 60434 73729 60814
rect 74109 60434 74121 60814
rect 74501 60434 74664 60814
rect 71998 60422 74664 60434
rect 71998 60042 72161 60422
rect 72541 60042 72553 60422
rect 72933 60042 72945 60422
rect 73325 60042 73337 60422
rect 73717 60042 73729 60422
rect 74109 60042 74121 60422
rect 74501 60042 74664 60422
rect 71998 60000 74664 60042
rect 87998 63558 90664 63600
rect 87998 63178 88161 63558
rect 88541 63178 88553 63558
rect 88933 63178 88945 63558
rect 89325 63178 89337 63558
rect 89717 63178 89729 63558
rect 90109 63178 90121 63558
rect 90501 63178 90664 63558
rect 87998 63166 90664 63178
rect 87998 62786 88161 63166
rect 88541 62786 88553 63166
rect 88933 62786 88945 63166
rect 89325 62786 89337 63166
rect 89717 62786 89729 63166
rect 90109 62786 90121 63166
rect 90501 62786 90664 63166
rect 87998 62774 90664 62786
rect 87998 62394 88161 62774
rect 88541 62394 88553 62774
rect 88933 62394 88945 62774
rect 89325 62394 89337 62774
rect 89717 62394 89729 62774
rect 90109 62394 90121 62774
rect 90501 62394 90664 62774
rect 87998 62382 90664 62394
rect 87998 62002 88161 62382
rect 88541 62002 88553 62382
rect 88933 62002 88945 62382
rect 89325 62002 89337 62382
rect 89717 62002 89729 62382
rect 90109 62002 90121 62382
rect 90501 62002 90664 62382
rect 87998 61990 90664 62002
rect 87998 61610 88161 61990
rect 88541 61610 88553 61990
rect 88933 61610 88945 61990
rect 89325 61610 89337 61990
rect 89717 61610 89729 61990
rect 90109 61610 90121 61990
rect 90501 61610 90664 61990
rect 87998 61598 90664 61610
rect 87998 61218 88161 61598
rect 88541 61218 88553 61598
rect 88933 61218 88945 61598
rect 89325 61218 89337 61598
rect 89717 61218 89729 61598
rect 90109 61218 90121 61598
rect 90501 61218 90664 61598
rect 87998 61206 90664 61218
rect 87998 60826 88161 61206
rect 88541 60826 88553 61206
rect 88933 60826 88945 61206
rect 89325 60826 89337 61206
rect 89717 60826 89729 61206
rect 90109 60826 90121 61206
rect 90501 60826 90664 61206
rect 87998 60814 90664 60826
rect 87998 60434 88161 60814
rect 88541 60434 88553 60814
rect 88933 60434 88945 60814
rect 89325 60434 89337 60814
rect 89717 60434 89729 60814
rect 90109 60434 90121 60814
rect 90501 60434 90664 60814
rect 87998 60422 90664 60434
rect 87998 60042 88161 60422
rect 88541 60042 88553 60422
rect 88933 60042 88945 60422
rect 89325 60042 89337 60422
rect 89717 60042 89729 60422
rect 90109 60042 90121 60422
rect 90501 60042 90664 60422
rect 87998 60000 90664 60042
rect 103998 63558 106664 63600
rect 103998 63178 104161 63558
rect 104541 63178 104553 63558
rect 104933 63178 104945 63558
rect 105325 63178 105337 63558
rect 105717 63178 105729 63558
rect 106109 63178 106121 63558
rect 106501 63178 106664 63558
rect 103998 63166 106664 63178
rect 103998 62786 104161 63166
rect 104541 62786 104553 63166
rect 104933 62786 104945 63166
rect 105325 62786 105337 63166
rect 105717 62786 105729 63166
rect 106109 62786 106121 63166
rect 106501 62786 106664 63166
rect 103998 62774 106664 62786
rect 103998 62394 104161 62774
rect 104541 62394 104553 62774
rect 104933 62394 104945 62774
rect 105325 62394 105337 62774
rect 105717 62394 105729 62774
rect 106109 62394 106121 62774
rect 106501 62394 106664 62774
rect 103998 62382 106664 62394
rect 103998 62002 104161 62382
rect 104541 62002 104553 62382
rect 104933 62002 104945 62382
rect 105325 62002 105337 62382
rect 105717 62002 105729 62382
rect 106109 62002 106121 62382
rect 106501 62002 106664 62382
rect 103998 61990 106664 62002
rect 103998 61610 104161 61990
rect 104541 61610 104553 61990
rect 104933 61610 104945 61990
rect 105325 61610 105337 61990
rect 105717 61610 105729 61990
rect 106109 61610 106121 61990
rect 106501 61610 106664 61990
rect 103998 61598 106664 61610
rect 103998 61218 104161 61598
rect 104541 61218 104553 61598
rect 104933 61218 104945 61598
rect 105325 61218 105337 61598
rect 105717 61218 105729 61598
rect 106109 61218 106121 61598
rect 106501 61218 106664 61598
rect 103998 61206 106664 61218
rect 103998 60826 104161 61206
rect 104541 60826 104553 61206
rect 104933 60826 104945 61206
rect 105325 60826 105337 61206
rect 105717 60826 105729 61206
rect 106109 60826 106121 61206
rect 106501 60826 106664 61206
rect 103998 60814 106664 60826
rect 103998 60434 104161 60814
rect 104541 60434 104553 60814
rect 104933 60434 104945 60814
rect 105325 60434 105337 60814
rect 105717 60434 105729 60814
rect 106109 60434 106121 60814
rect 106501 60434 106664 60814
rect 103998 60422 106664 60434
rect 103998 60042 104161 60422
rect 104541 60042 104553 60422
rect 104933 60042 104945 60422
rect 105325 60042 105337 60422
rect 105717 60042 105729 60422
rect 106109 60042 106121 60422
rect 106501 60042 106664 60422
rect 103998 60000 106664 60042
rect 119998 63558 122664 63600
rect 119998 63178 120161 63558
rect 120541 63178 120553 63558
rect 120933 63178 120945 63558
rect 121325 63178 121337 63558
rect 121717 63178 121729 63558
rect 122109 63178 122121 63558
rect 122501 63178 122664 63558
rect 119998 63166 122664 63178
rect 119998 62786 120161 63166
rect 120541 62786 120553 63166
rect 120933 62786 120945 63166
rect 121325 62786 121337 63166
rect 121717 62786 121729 63166
rect 122109 62786 122121 63166
rect 122501 62786 122664 63166
rect 119998 62774 122664 62786
rect 119998 62394 120161 62774
rect 120541 62394 120553 62774
rect 120933 62394 120945 62774
rect 121325 62394 121337 62774
rect 121717 62394 121729 62774
rect 122109 62394 122121 62774
rect 122501 62394 122664 62774
rect 119998 62382 122664 62394
rect 119998 62002 120161 62382
rect 120541 62002 120553 62382
rect 120933 62002 120945 62382
rect 121325 62002 121337 62382
rect 121717 62002 121729 62382
rect 122109 62002 122121 62382
rect 122501 62002 122664 62382
rect 119998 61990 122664 62002
rect 119998 61610 120161 61990
rect 120541 61610 120553 61990
rect 120933 61610 120945 61990
rect 121325 61610 121337 61990
rect 121717 61610 121729 61990
rect 122109 61610 122121 61990
rect 122501 61610 122664 61990
rect 119998 61598 122664 61610
rect 119998 61218 120161 61598
rect 120541 61218 120553 61598
rect 120933 61218 120945 61598
rect 121325 61218 121337 61598
rect 121717 61218 121729 61598
rect 122109 61218 122121 61598
rect 122501 61218 122664 61598
rect 119998 61206 122664 61218
rect 119998 60826 120161 61206
rect 120541 60826 120553 61206
rect 120933 60826 120945 61206
rect 121325 60826 121337 61206
rect 121717 60826 121729 61206
rect 122109 60826 122121 61206
rect 122501 60826 122664 61206
rect 119998 60814 122664 60826
rect 119998 60434 120161 60814
rect 120541 60434 120553 60814
rect 120933 60434 120945 60814
rect 121325 60434 121337 60814
rect 121717 60434 121729 60814
rect 122109 60434 122121 60814
rect 122501 60434 122664 60814
rect 119998 60422 122664 60434
rect 119998 60042 120161 60422
rect 120541 60042 120553 60422
rect 120933 60042 120945 60422
rect 121325 60042 121337 60422
rect 121717 60042 121729 60422
rect 122109 60042 122121 60422
rect 122501 60042 122664 60422
rect 119998 60000 122664 60042
rect 132000 63558 136000 63600
rect 132000 63178 132046 63558
rect 132426 63178 132438 63558
rect 132818 63178 132830 63558
rect 133210 63178 133222 63558
rect 133602 63178 133614 63558
rect 133994 63178 134006 63558
rect 134386 63178 134398 63558
rect 134778 63178 134790 63558
rect 135170 63178 135182 63558
rect 135562 63178 135574 63558
rect 135954 63178 136000 63558
rect 132000 63166 136000 63178
rect 132000 62786 132046 63166
rect 132426 62786 132438 63166
rect 132818 62786 132830 63166
rect 133210 62786 133222 63166
rect 133602 62786 133614 63166
rect 133994 62786 134006 63166
rect 134386 62786 134398 63166
rect 134778 62786 134790 63166
rect 135170 62786 135182 63166
rect 135562 62786 135574 63166
rect 135954 62786 136000 63166
rect 132000 62774 136000 62786
rect 132000 62394 132046 62774
rect 132426 62394 132438 62774
rect 132818 62394 132830 62774
rect 133210 62394 133222 62774
rect 133602 62394 133614 62774
rect 133994 62394 134006 62774
rect 134386 62394 134398 62774
rect 134778 62394 134790 62774
rect 135170 62394 135182 62774
rect 135562 62394 135574 62774
rect 135954 62394 136000 62774
rect 132000 62382 136000 62394
rect 132000 62002 132046 62382
rect 132426 62002 132438 62382
rect 132818 62002 132830 62382
rect 133210 62002 133222 62382
rect 133602 62002 133614 62382
rect 133994 62002 134006 62382
rect 134386 62002 134398 62382
rect 134778 62002 134790 62382
rect 135170 62002 135182 62382
rect 135562 62002 135574 62382
rect 135954 62002 136000 62382
rect 132000 61990 136000 62002
rect 132000 61610 132046 61990
rect 132426 61610 132438 61990
rect 132818 61610 132830 61990
rect 133210 61610 133222 61990
rect 133602 61610 133614 61990
rect 133994 61610 134006 61990
rect 134386 61610 134398 61990
rect 134778 61610 134790 61990
rect 135170 61610 135182 61990
rect 135562 61610 135574 61990
rect 135954 61610 136000 61990
rect 132000 61598 136000 61610
rect 132000 61218 132046 61598
rect 132426 61218 132438 61598
rect 132818 61218 132830 61598
rect 133210 61218 133222 61598
rect 133602 61218 133614 61598
rect 133994 61218 134006 61598
rect 134386 61218 134398 61598
rect 134778 61218 134790 61598
rect 135170 61218 135182 61598
rect 135562 61218 135574 61598
rect 135954 61218 136000 61598
rect 132000 61206 136000 61218
rect 132000 60826 132046 61206
rect 132426 60826 132438 61206
rect 132818 60826 132830 61206
rect 133210 60826 133222 61206
rect 133602 60826 133614 61206
rect 133994 60826 134006 61206
rect 134386 60826 134398 61206
rect 134778 60826 134790 61206
rect 135170 60826 135182 61206
rect 135562 60826 135574 61206
rect 135954 60826 136000 61206
rect 132000 60814 136000 60826
rect 132000 60434 132046 60814
rect 132426 60434 132438 60814
rect 132818 60434 132830 60814
rect 133210 60434 133222 60814
rect 133602 60434 133614 60814
rect 133994 60434 134006 60814
rect 134386 60434 134398 60814
rect 134778 60434 134790 60814
rect 135170 60434 135182 60814
rect 135562 60434 135574 60814
rect 135954 60434 136000 60814
rect 132000 60422 136000 60434
rect 132000 60042 132046 60422
rect 132426 60042 132438 60422
rect 132818 60042 132830 60422
rect 133210 60042 133222 60422
rect 133602 60042 133614 60422
rect 133994 60042 134006 60422
rect 134386 60042 134398 60422
rect 134778 60042 134790 60422
rect 135170 60042 135182 60422
rect 135562 60042 135574 60422
rect 135954 60042 136000 60422
rect 132000 60000 136000 60042
rect 151998 63558 154664 63600
rect 151998 63178 152161 63558
rect 152541 63178 152553 63558
rect 152933 63178 152945 63558
rect 153325 63178 153337 63558
rect 153717 63178 153729 63558
rect 154109 63178 154121 63558
rect 154501 63178 154664 63558
rect 151998 63166 154664 63178
rect 151998 62786 152161 63166
rect 152541 62786 152553 63166
rect 152933 62786 152945 63166
rect 153325 62786 153337 63166
rect 153717 62786 153729 63166
rect 154109 62786 154121 63166
rect 154501 62786 154664 63166
rect 151998 62774 154664 62786
rect 151998 62394 152161 62774
rect 152541 62394 152553 62774
rect 152933 62394 152945 62774
rect 153325 62394 153337 62774
rect 153717 62394 153729 62774
rect 154109 62394 154121 62774
rect 154501 62394 154664 62774
rect 151998 62382 154664 62394
rect 151998 62002 152161 62382
rect 152541 62002 152553 62382
rect 152933 62002 152945 62382
rect 153325 62002 153337 62382
rect 153717 62002 153729 62382
rect 154109 62002 154121 62382
rect 154501 62002 154664 62382
rect 151998 61990 154664 62002
rect 151998 61610 152161 61990
rect 152541 61610 152553 61990
rect 152933 61610 152945 61990
rect 153325 61610 153337 61990
rect 153717 61610 153729 61990
rect 154109 61610 154121 61990
rect 154501 61610 154664 61990
rect 151998 61598 154664 61610
rect 151998 61218 152161 61598
rect 152541 61218 152553 61598
rect 152933 61218 152945 61598
rect 153325 61218 153337 61598
rect 153717 61218 153729 61598
rect 154109 61218 154121 61598
rect 154501 61218 154664 61598
rect 151998 61206 154664 61218
rect 151998 60826 152161 61206
rect 152541 60826 152553 61206
rect 152933 60826 152945 61206
rect 153325 60826 153337 61206
rect 153717 60826 153729 61206
rect 154109 60826 154121 61206
rect 154501 60826 154664 61206
rect 151998 60814 154664 60826
rect 151998 60434 152161 60814
rect 152541 60434 152553 60814
rect 152933 60434 152945 60814
rect 153325 60434 153337 60814
rect 153717 60434 153729 60814
rect 154109 60434 154121 60814
rect 154501 60434 154664 60814
rect 151998 60422 154664 60434
rect 151998 60042 152161 60422
rect 152541 60042 152553 60422
rect 152933 60042 152945 60422
rect 153325 60042 153337 60422
rect 153717 60042 153729 60422
rect 154109 60042 154121 60422
rect 154501 60042 154664 60422
rect 151998 60000 154664 60042
rect 82666 59558 85332 59600
rect 82666 59178 82829 59558
rect 83209 59178 83221 59558
rect 83601 59178 83613 59558
rect 83993 59178 84005 59558
rect 84385 59178 84397 59558
rect 84777 59178 84789 59558
rect 85169 59178 85332 59558
rect 82666 59166 85332 59178
rect 82666 58786 82829 59166
rect 83209 58786 83221 59166
rect 83601 58786 83613 59166
rect 83993 58786 84005 59166
rect 84385 58786 84397 59166
rect 84777 58786 84789 59166
rect 85169 58786 85332 59166
rect 82666 58774 85332 58786
rect 82666 58394 82829 58774
rect 83209 58394 83221 58774
rect 83601 58394 83613 58774
rect 83993 58394 84005 58774
rect 84385 58394 84397 58774
rect 84777 58394 84789 58774
rect 85169 58394 85332 58774
rect 82666 58382 85332 58394
rect 82666 58002 82829 58382
rect 83209 58002 83221 58382
rect 83601 58002 83613 58382
rect 83993 58002 84005 58382
rect 84385 58002 84397 58382
rect 84777 58002 84789 58382
rect 85169 58002 85332 58382
rect 82666 57990 85332 58002
rect 82666 57610 82829 57990
rect 83209 57610 83221 57990
rect 83601 57610 83613 57990
rect 83993 57610 84005 57990
rect 84385 57610 84397 57990
rect 84777 57610 84789 57990
rect 85169 57610 85332 57990
rect 82666 57598 85332 57610
rect 82666 57218 82829 57598
rect 83209 57218 83221 57598
rect 83601 57218 83613 57598
rect 83993 57218 84005 57598
rect 84385 57218 84397 57598
rect 84777 57218 84789 57598
rect 85169 57218 85332 57598
rect 82666 57206 85332 57218
rect 82666 56826 82829 57206
rect 83209 56826 83221 57206
rect 83601 56826 83613 57206
rect 83993 56826 84005 57206
rect 84385 56826 84397 57206
rect 84777 56826 84789 57206
rect 85169 56826 85332 57206
rect 82666 56814 85332 56826
rect 82666 56434 82829 56814
rect 83209 56434 83221 56814
rect 83601 56434 83613 56814
rect 83993 56434 84005 56814
rect 84385 56434 84397 56814
rect 84777 56434 84789 56814
rect 85169 56434 85332 56814
rect 82666 56422 85332 56434
rect 82666 56042 82829 56422
rect 83209 56042 83221 56422
rect 83601 56042 83613 56422
rect 83993 56042 84005 56422
rect 84385 56042 84397 56422
rect 84777 56042 84789 56422
rect 85169 56042 85332 56422
rect 82666 56000 85332 56042
rect 98666 59558 101332 59600
rect 98666 59178 98829 59558
rect 99209 59178 99221 59558
rect 99601 59178 99613 59558
rect 99993 59178 100005 59558
rect 100385 59178 100397 59558
rect 100777 59178 100789 59558
rect 101169 59178 101332 59558
rect 98666 59166 101332 59178
rect 98666 58786 98829 59166
rect 99209 58786 99221 59166
rect 99601 58786 99613 59166
rect 99993 58786 100005 59166
rect 100385 58786 100397 59166
rect 100777 58786 100789 59166
rect 101169 58786 101332 59166
rect 98666 58774 101332 58786
rect 98666 58394 98829 58774
rect 99209 58394 99221 58774
rect 99601 58394 99613 58774
rect 99993 58394 100005 58774
rect 100385 58394 100397 58774
rect 100777 58394 100789 58774
rect 101169 58394 101332 58774
rect 98666 58382 101332 58394
rect 98666 58002 98829 58382
rect 99209 58002 99221 58382
rect 99601 58002 99613 58382
rect 99993 58002 100005 58382
rect 100385 58002 100397 58382
rect 100777 58002 100789 58382
rect 101169 58002 101332 58382
rect 98666 57990 101332 58002
rect 98666 57610 98829 57990
rect 99209 57610 99221 57990
rect 99601 57610 99613 57990
rect 99993 57610 100005 57990
rect 100385 57610 100397 57990
rect 100777 57610 100789 57990
rect 101169 57610 101332 57990
rect 98666 57598 101332 57610
rect 98666 57218 98829 57598
rect 99209 57218 99221 57598
rect 99601 57218 99613 57598
rect 99993 57218 100005 57598
rect 100385 57218 100397 57598
rect 100777 57218 100789 57598
rect 101169 57218 101332 57598
rect 98666 57206 101332 57218
rect 98666 56826 98829 57206
rect 99209 56826 99221 57206
rect 99601 56826 99613 57206
rect 99993 56826 100005 57206
rect 100385 56826 100397 57206
rect 100777 56826 100789 57206
rect 101169 56826 101332 57206
rect 98666 56814 101332 56826
rect 98666 56434 98829 56814
rect 99209 56434 99221 56814
rect 99601 56434 99613 56814
rect 99993 56434 100005 56814
rect 100385 56434 100397 56814
rect 100777 56434 100789 56814
rect 101169 56434 101332 56814
rect 98666 56422 101332 56434
rect 98666 56042 98829 56422
rect 99209 56042 99221 56422
rect 99601 56042 99613 56422
rect 99993 56042 100005 56422
rect 100385 56042 100397 56422
rect 100777 56042 100789 56422
rect 101169 56042 101332 56422
rect 98666 56000 101332 56042
rect 114666 59558 117332 59600
rect 114666 59178 114829 59558
rect 115209 59178 115221 59558
rect 115601 59178 115613 59558
rect 115993 59178 116005 59558
rect 116385 59178 116397 59558
rect 116777 59178 116789 59558
rect 117169 59178 117332 59558
rect 114666 59166 117332 59178
rect 114666 58786 114829 59166
rect 115209 58786 115221 59166
rect 115601 58786 115613 59166
rect 115993 58786 116005 59166
rect 116385 58786 116397 59166
rect 116777 58786 116789 59166
rect 117169 58786 117332 59166
rect 114666 58774 117332 58786
rect 114666 58394 114829 58774
rect 115209 58394 115221 58774
rect 115601 58394 115613 58774
rect 115993 58394 116005 58774
rect 116385 58394 116397 58774
rect 116777 58394 116789 58774
rect 117169 58394 117332 58774
rect 114666 58382 117332 58394
rect 114666 58002 114829 58382
rect 115209 58002 115221 58382
rect 115601 58002 115613 58382
rect 115993 58002 116005 58382
rect 116385 58002 116397 58382
rect 116777 58002 116789 58382
rect 117169 58002 117332 58382
rect 114666 57990 117332 58002
rect 114666 57610 114829 57990
rect 115209 57610 115221 57990
rect 115601 57610 115613 57990
rect 115993 57610 116005 57990
rect 116385 57610 116397 57990
rect 116777 57610 116789 57990
rect 117169 57610 117332 57990
rect 114666 57598 117332 57610
rect 114666 57218 114829 57598
rect 115209 57218 115221 57598
rect 115601 57218 115613 57598
rect 115993 57218 116005 57598
rect 116385 57218 116397 57598
rect 116777 57218 116789 57598
rect 117169 57218 117332 57598
rect 114666 57206 117332 57218
rect 114666 56826 114829 57206
rect 115209 56826 115221 57206
rect 115601 56826 115613 57206
rect 115993 56826 116005 57206
rect 116385 56826 116397 57206
rect 116777 56826 116789 57206
rect 117169 56826 117332 57206
rect 114666 56814 117332 56826
rect 114666 56434 114829 56814
rect 115209 56434 115221 56814
rect 115601 56434 115613 56814
rect 115993 56434 116005 56814
rect 116385 56434 116397 56814
rect 116777 56434 116789 56814
rect 117169 56434 117332 56814
rect 114666 56422 117332 56434
rect 114666 56042 114829 56422
rect 115209 56042 115221 56422
rect 115601 56042 115613 56422
rect 115993 56042 116005 56422
rect 116385 56042 116397 56422
rect 116777 56042 116789 56422
rect 117169 56042 117332 56422
rect 114666 56000 117332 56042
rect 146666 59558 149332 59600
rect 146666 59178 146829 59558
rect 147209 59178 147221 59558
rect 147601 59178 147613 59558
rect 147993 59178 148005 59558
rect 148385 59178 148397 59558
rect 148777 59178 148789 59558
rect 149169 59178 149332 59558
rect 146666 59166 149332 59178
rect 146666 58786 146829 59166
rect 147209 58786 147221 59166
rect 147601 58786 147613 59166
rect 147993 58786 148005 59166
rect 148385 58786 148397 59166
rect 148777 58786 148789 59166
rect 149169 58786 149332 59166
rect 146666 58774 149332 58786
rect 146666 58394 146829 58774
rect 147209 58394 147221 58774
rect 147601 58394 147613 58774
rect 147993 58394 148005 58774
rect 148385 58394 148397 58774
rect 148777 58394 148789 58774
rect 149169 58394 149332 58774
rect 146666 58382 149332 58394
rect 146666 58002 146829 58382
rect 147209 58002 147221 58382
rect 147601 58002 147613 58382
rect 147993 58002 148005 58382
rect 148385 58002 148397 58382
rect 148777 58002 148789 58382
rect 149169 58002 149332 58382
rect 146666 57990 149332 58002
rect 146666 57610 146829 57990
rect 147209 57610 147221 57990
rect 147601 57610 147613 57990
rect 147993 57610 148005 57990
rect 148385 57610 148397 57990
rect 148777 57610 148789 57990
rect 149169 57610 149332 57990
rect 146666 57598 149332 57610
rect 146666 57218 146829 57598
rect 147209 57218 147221 57598
rect 147601 57218 147613 57598
rect 147993 57218 148005 57598
rect 148385 57218 148397 57598
rect 148777 57218 148789 57598
rect 149169 57218 149332 57598
rect 146666 57206 149332 57218
rect 146666 56826 146829 57206
rect 147209 56826 147221 57206
rect 147601 56826 147613 57206
rect 147993 56826 148005 57206
rect 148385 56826 148397 57206
rect 148777 56826 148789 57206
rect 149169 56826 149332 57206
rect 146666 56814 149332 56826
rect 146666 56434 146829 56814
rect 147209 56434 147221 56814
rect 147601 56434 147613 56814
rect 147993 56434 148005 56814
rect 148385 56434 148397 56814
rect 148777 56434 148789 56814
rect 149169 56434 149332 56814
rect 146666 56422 149332 56434
rect 146666 56042 146829 56422
rect 147209 56042 147221 56422
rect 147601 56042 147613 56422
rect 147993 56042 148005 56422
rect 148385 56042 148397 56422
rect 148777 56042 148789 56422
rect 149169 56042 149332 56422
rect 146666 56000 149332 56042
<< via6 >>
rect 82829 167578 83209 167958
rect 83221 167578 83601 167958
rect 83613 167578 83993 167958
rect 84005 167578 84385 167958
rect 84397 167578 84777 167958
rect 84789 167578 85169 167958
rect 82829 167186 83209 167566
rect 83221 167186 83601 167566
rect 83613 167186 83993 167566
rect 84005 167186 84385 167566
rect 84397 167186 84777 167566
rect 84789 167186 85169 167566
rect 82829 166794 83209 167174
rect 83221 166794 83601 167174
rect 83613 166794 83993 167174
rect 84005 166794 84385 167174
rect 84397 166794 84777 167174
rect 84789 166794 85169 167174
rect 82829 166402 83209 166782
rect 83221 166402 83601 166782
rect 83613 166402 83993 166782
rect 84005 166402 84385 166782
rect 84397 166402 84777 166782
rect 84789 166402 85169 166782
rect 82829 166010 83209 166390
rect 83221 166010 83601 166390
rect 83613 166010 83993 166390
rect 84005 166010 84385 166390
rect 84397 166010 84777 166390
rect 84789 166010 85169 166390
rect 82829 165618 83209 165998
rect 83221 165618 83601 165998
rect 83613 165618 83993 165998
rect 84005 165618 84385 165998
rect 84397 165618 84777 165998
rect 84789 165618 85169 165998
rect 82829 165226 83209 165606
rect 83221 165226 83601 165606
rect 83613 165226 83993 165606
rect 84005 165226 84385 165606
rect 84397 165226 84777 165606
rect 84789 165226 85169 165606
rect 82829 164834 83209 165214
rect 83221 164834 83601 165214
rect 83613 164834 83993 165214
rect 84005 164834 84385 165214
rect 84397 164834 84777 165214
rect 84789 164834 85169 165214
rect 82829 164442 83209 164822
rect 83221 164442 83601 164822
rect 83613 164442 83993 164822
rect 84005 164442 84385 164822
rect 84397 164442 84777 164822
rect 84789 164442 85169 164822
rect 98829 167578 99209 167958
rect 99221 167578 99601 167958
rect 99613 167578 99993 167958
rect 100005 167578 100385 167958
rect 100397 167578 100777 167958
rect 100789 167578 101169 167958
rect 98829 167186 99209 167566
rect 99221 167186 99601 167566
rect 99613 167186 99993 167566
rect 100005 167186 100385 167566
rect 100397 167186 100777 167566
rect 100789 167186 101169 167566
rect 98829 166794 99209 167174
rect 99221 166794 99601 167174
rect 99613 166794 99993 167174
rect 100005 166794 100385 167174
rect 100397 166794 100777 167174
rect 100789 166794 101169 167174
rect 98829 166402 99209 166782
rect 99221 166402 99601 166782
rect 99613 166402 99993 166782
rect 100005 166402 100385 166782
rect 100397 166402 100777 166782
rect 100789 166402 101169 166782
rect 98829 166010 99209 166390
rect 99221 166010 99601 166390
rect 99613 166010 99993 166390
rect 100005 166010 100385 166390
rect 100397 166010 100777 166390
rect 100789 166010 101169 166390
rect 98829 165618 99209 165998
rect 99221 165618 99601 165998
rect 99613 165618 99993 165998
rect 100005 165618 100385 165998
rect 100397 165618 100777 165998
rect 100789 165618 101169 165998
rect 98829 165226 99209 165606
rect 99221 165226 99601 165606
rect 99613 165226 99993 165606
rect 100005 165226 100385 165606
rect 100397 165226 100777 165606
rect 100789 165226 101169 165606
rect 98829 164834 99209 165214
rect 99221 164834 99601 165214
rect 99613 164834 99993 165214
rect 100005 164834 100385 165214
rect 100397 164834 100777 165214
rect 100789 164834 101169 165214
rect 98829 164442 99209 164822
rect 99221 164442 99601 164822
rect 99613 164442 99993 164822
rect 100005 164442 100385 164822
rect 100397 164442 100777 164822
rect 100789 164442 101169 164822
rect 114829 167578 115209 167958
rect 115221 167578 115601 167958
rect 115613 167578 115993 167958
rect 116005 167578 116385 167958
rect 116397 167578 116777 167958
rect 116789 167578 117169 167958
rect 114829 167186 115209 167566
rect 115221 167186 115601 167566
rect 115613 167186 115993 167566
rect 116005 167186 116385 167566
rect 116397 167186 116777 167566
rect 116789 167186 117169 167566
rect 114829 166794 115209 167174
rect 115221 166794 115601 167174
rect 115613 166794 115993 167174
rect 116005 166794 116385 167174
rect 116397 166794 116777 167174
rect 116789 166794 117169 167174
rect 114829 166402 115209 166782
rect 115221 166402 115601 166782
rect 115613 166402 115993 166782
rect 116005 166402 116385 166782
rect 116397 166402 116777 166782
rect 116789 166402 117169 166782
rect 114829 166010 115209 166390
rect 115221 166010 115601 166390
rect 115613 166010 115993 166390
rect 116005 166010 116385 166390
rect 116397 166010 116777 166390
rect 116789 166010 117169 166390
rect 114829 165618 115209 165998
rect 115221 165618 115601 165998
rect 115613 165618 115993 165998
rect 116005 165618 116385 165998
rect 116397 165618 116777 165998
rect 116789 165618 117169 165998
rect 114829 165226 115209 165606
rect 115221 165226 115601 165606
rect 115613 165226 115993 165606
rect 116005 165226 116385 165606
rect 116397 165226 116777 165606
rect 116789 165226 117169 165606
rect 114829 164834 115209 165214
rect 115221 164834 115601 165214
rect 115613 164834 115993 165214
rect 116005 164834 116385 165214
rect 116397 164834 116777 165214
rect 116789 164834 117169 165214
rect 114829 164442 115209 164822
rect 115221 164442 115601 164822
rect 115613 164442 115993 164822
rect 116005 164442 116385 164822
rect 116397 164442 116777 164822
rect 116789 164442 117169 164822
rect 130829 167578 131209 167958
rect 131221 167578 131601 167958
rect 131613 167578 131993 167958
rect 132005 167578 132385 167958
rect 132397 167578 132777 167958
rect 132789 167578 133169 167958
rect 130829 167186 131209 167566
rect 131221 167186 131601 167566
rect 131613 167186 131993 167566
rect 132005 167186 132385 167566
rect 132397 167186 132777 167566
rect 132789 167186 133169 167566
rect 130829 166794 131209 167174
rect 131221 166794 131601 167174
rect 131613 166794 131993 167174
rect 132005 166794 132385 167174
rect 132397 166794 132777 167174
rect 132789 166794 133169 167174
rect 130829 166402 131209 166782
rect 131221 166402 131601 166782
rect 131613 166402 131993 166782
rect 132005 166402 132385 166782
rect 132397 166402 132777 166782
rect 132789 166402 133169 166782
rect 130829 166010 131209 166390
rect 131221 166010 131601 166390
rect 131613 166010 131993 166390
rect 132005 166010 132385 166390
rect 132397 166010 132777 166390
rect 132789 166010 133169 166390
rect 130829 165618 131209 165998
rect 131221 165618 131601 165998
rect 131613 165618 131993 165998
rect 132005 165618 132385 165998
rect 132397 165618 132777 165998
rect 132789 165618 133169 165998
rect 130829 165226 131209 165606
rect 131221 165226 131601 165606
rect 131613 165226 131993 165606
rect 132005 165226 132385 165606
rect 132397 165226 132777 165606
rect 132789 165226 133169 165606
rect 130829 164834 131209 165214
rect 131221 164834 131601 165214
rect 131613 164834 131993 165214
rect 132005 164834 132385 165214
rect 132397 164834 132777 165214
rect 132789 164834 133169 165214
rect 130829 164442 131209 164822
rect 131221 164442 131601 164822
rect 131613 164442 131993 164822
rect 132005 164442 132385 164822
rect 132397 164442 132777 164822
rect 132789 164442 133169 164822
rect 146829 167578 147209 167958
rect 147221 167578 147601 167958
rect 147613 167578 147993 167958
rect 148005 167578 148385 167958
rect 148397 167578 148777 167958
rect 148789 167578 149169 167958
rect 146829 167186 147209 167566
rect 147221 167186 147601 167566
rect 147613 167186 147993 167566
rect 148005 167186 148385 167566
rect 148397 167186 148777 167566
rect 148789 167186 149169 167566
rect 146829 166794 147209 167174
rect 147221 166794 147601 167174
rect 147613 166794 147993 167174
rect 148005 166794 148385 167174
rect 148397 166794 148777 167174
rect 148789 166794 149169 167174
rect 146829 166402 147209 166782
rect 147221 166402 147601 166782
rect 147613 166402 147993 166782
rect 148005 166402 148385 166782
rect 148397 166402 148777 166782
rect 148789 166402 149169 166782
rect 146829 166010 147209 166390
rect 147221 166010 147601 166390
rect 147613 166010 147993 166390
rect 148005 166010 148385 166390
rect 148397 166010 148777 166390
rect 148789 166010 149169 166390
rect 146829 165618 147209 165998
rect 147221 165618 147601 165998
rect 147613 165618 147993 165998
rect 148005 165618 148385 165998
rect 148397 165618 148777 165998
rect 148789 165618 149169 165998
rect 146829 165226 147209 165606
rect 147221 165226 147601 165606
rect 147613 165226 147993 165606
rect 148005 165226 148385 165606
rect 148397 165226 148777 165606
rect 148789 165226 149169 165606
rect 146829 164834 147209 165214
rect 147221 164834 147601 165214
rect 147613 164834 147993 165214
rect 148005 164834 148385 165214
rect 148397 164834 148777 165214
rect 148789 164834 149169 165214
rect 146829 164442 147209 164822
rect 147221 164442 147601 164822
rect 147613 164442 147993 164822
rect 148005 164442 148385 164822
rect 148397 164442 148777 164822
rect 148789 164442 149169 164822
rect 72161 163578 72541 163958
rect 72553 163578 72933 163958
rect 72945 163578 73325 163958
rect 73337 163578 73717 163958
rect 73729 163578 74109 163958
rect 74121 163578 74501 163958
rect 72161 163186 72541 163566
rect 72553 163186 72933 163566
rect 72945 163186 73325 163566
rect 73337 163186 73717 163566
rect 73729 163186 74109 163566
rect 74121 163186 74501 163566
rect 72161 162794 72541 163174
rect 72553 162794 72933 163174
rect 72945 162794 73325 163174
rect 73337 162794 73717 163174
rect 73729 162794 74109 163174
rect 74121 162794 74501 163174
rect 72161 162402 72541 162782
rect 72553 162402 72933 162782
rect 72945 162402 73325 162782
rect 73337 162402 73717 162782
rect 73729 162402 74109 162782
rect 74121 162402 74501 162782
rect 72161 162010 72541 162390
rect 72553 162010 72933 162390
rect 72945 162010 73325 162390
rect 73337 162010 73717 162390
rect 73729 162010 74109 162390
rect 74121 162010 74501 162390
rect 72161 161618 72541 161998
rect 72553 161618 72933 161998
rect 72945 161618 73325 161998
rect 73337 161618 73717 161998
rect 73729 161618 74109 161998
rect 74121 161618 74501 161998
rect 72161 161226 72541 161606
rect 72553 161226 72933 161606
rect 72945 161226 73325 161606
rect 73337 161226 73717 161606
rect 73729 161226 74109 161606
rect 74121 161226 74501 161606
rect 72161 160834 72541 161214
rect 72553 160834 72933 161214
rect 72945 160834 73325 161214
rect 73337 160834 73717 161214
rect 73729 160834 74109 161214
rect 74121 160834 74501 161214
rect 72161 160442 72541 160822
rect 72553 160442 72933 160822
rect 72945 160442 73325 160822
rect 73337 160442 73717 160822
rect 73729 160442 74109 160822
rect 74121 160442 74501 160822
rect 88161 163578 88541 163958
rect 88553 163578 88933 163958
rect 88945 163578 89325 163958
rect 89337 163578 89717 163958
rect 89729 163578 90109 163958
rect 90121 163578 90501 163958
rect 88161 163186 88541 163566
rect 88553 163186 88933 163566
rect 88945 163186 89325 163566
rect 89337 163186 89717 163566
rect 89729 163186 90109 163566
rect 90121 163186 90501 163566
rect 88161 162794 88541 163174
rect 88553 162794 88933 163174
rect 88945 162794 89325 163174
rect 89337 162794 89717 163174
rect 89729 162794 90109 163174
rect 90121 162794 90501 163174
rect 88161 162402 88541 162782
rect 88553 162402 88933 162782
rect 88945 162402 89325 162782
rect 89337 162402 89717 162782
rect 89729 162402 90109 162782
rect 90121 162402 90501 162782
rect 88161 162010 88541 162390
rect 88553 162010 88933 162390
rect 88945 162010 89325 162390
rect 89337 162010 89717 162390
rect 89729 162010 90109 162390
rect 90121 162010 90501 162390
rect 88161 161618 88541 161998
rect 88553 161618 88933 161998
rect 88945 161618 89325 161998
rect 89337 161618 89717 161998
rect 89729 161618 90109 161998
rect 90121 161618 90501 161998
rect 88161 161226 88541 161606
rect 88553 161226 88933 161606
rect 88945 161226 89325 161606
rect 89337 161226 89717 161606
rect 89729 161226 90109 161606
rect 90121 161226 90501 161606
rect 88161 160834 88541 161214
rect 88553 160834 88933 161214
rect 88945 160834 89325 161214
rect 89337 160834 89717 161214
rect 89729 160834 90109 161214
rect 90121 160834 90501 161214
rect 88161 160442 88541 160822
rect 88553 160442 88933 160822
rect 88945 160442 89325 160822
rect 89337 160442 89717 160822
rect 89729 160442 90109 160822
rect 90121 160442 90501 160822
rect 104161 163578 104541 163958
rect 104553 163578 104933 163958
rect 104945 163578 105325 163958
rect 105337 163578 105717 163958
rect 105729 163578 106109 163958
rect 106121 163578 106501 163958
rect 104161 163186 104541 163566
rect 104553 163186 104933 163566
rect 104945 163186 105325 163566
rect 105337 163186 105717 163566
rect 105729 163186 106109 163566
rect 106121 163186 106501 163566
rect 104161 162794 104541 163174
rect 104553 162794 104933 163174
rect 104945 162794 105325 163174
rect 105337 162794 105717 163174
rect 105729 162794 106109 163174
rect 106121 162794 106501 163174
rect 104161 162402 104541 162782
rect 104553 162402 104933 162782
rect 104945 162402 105325 162782
rect 105337 162402 105717 162782
rect 105729 162402 106109 162782
rect 106121 162402 106501 162782
rect 104161 162010 104541 162390
rect 104553 162010 104933 162390
rect 104945 162010 105325 162390
rect 105337 162010 105717 162390
rect 105729 162010 106109 162390
rect 106121 162010 106501 162390
rect 104161 161618 104541 161998
rect 104553 161618 104933 161998
rect 104945 161618 105325 161998
rect 105337 161618 105717 161998
rect 105729 161618 106109 161998
rect 106121 161618 106501 161998
rect 104161 161226 104541 161606
rect 104553 161226 104933 161606
rect 104945 161226 105325 161606
rect 105337 161226 105717 161606
rect 105729 161226 106109 161606
rect 106121 161226 106501 161606
rect 104161 160834 104541 161214
rect 104553 160834 104933 161214
rect 104945 160834 105325 161214
rect 105337 160834 105717 161214
rect 105729 160834 106109 161214
rect 106121 160834 106501 161214
rect 104161 160442 104541 160822
rect 104553 160442 104933 160822
rect 104945 160442 105325 160822
rect 105337 160442 105717 160822
rect 105729 160442 106109 160822
rect 106121 160442 106501 160822
rect 120161 163578 120541 163958
rect 120553 163578 120933 163958
rect 120945 163578 121325 163958
rect 121337 163578 121717 163958
rect 121729 163578 122109 163958
rect 122121 163578 122501 163958
rect 120161 163186 120541 163566
rect 120553 163186 120933 163566
rect 120945 163186 121325 163566
rect 121337 163186 121717 163566
rect 121729 163186 122109 163566
rect 122121 163186 122501 163566
rect 120161 162794 120541 163174
rect 120553 162794 120933 163174
rect 120945 162794 121325 163174
rect 121337 162794 121717 163174
rect 121729 162794 122109 163174
rect 122121 162794 122501 163174
rect 120161 162402 120541 162782
rect 120553 162402 120933 162782
rect 120945 162402 121325 162782
rect 121337 162402 121717 162782
rect 121729 162402 122109 162782
rect 122121 162402 122501 162782
rect 120161 162010 120541 162390
rect 120553 162010 120933 162390
rect 120945 162010 121325 162390
rect 121337 162010 121717 162390
rect 121729 162010 122109 162390
rect 122121 162010 122501 162390
rect 120161 161618 120541 161998
rect 120553 161618 120933 161998
rect 120945 161618 121325 161998
rect 121337 161618 121717 161998
rect 121729 161618 122109 161998
rect 122121 161618 122501 161998
rect 120161 161226 120541 161606
rect 120553 161226 120933 161606
rect 120945 161226 121325 161606
rect 121337 161226 121717 161606
rect 121729 161226 122109 161606
rect 122121 161226 122501 161606
rect 120161 160834 120541 161214
rect 120553 160834 120933 161214
rect 120945 160834 121325 161214
rect 121337 160834 121717 161214
rect 121729 160834 122109 161214
rect 122121 160834 122501 161214
rect 120161 160442 120541 160822
rect 120553 160442 120933 160822
rect 120945 160442 121325 160822
rect 121337 160442 121717 160822
rect 121729 160442 122109 160822
rect 122121 160442 122501 160822
rect 136161 163578 136541 163958
rect 136553 163578 136933 163958
rect 136945 163578 137325 163958
rect 137337 163578 137717 163958
rect 137729 163578 138109 163958
rect 138121 163578 138501 163958
rect 136161 163186 136541 163566
rect 136553 163186 136933 163566
rect 136945 163186 137325 163566
rect 137337 163186 137717 163566
rect 137729 163186 138109 163566
rect 138121 163186 138501 163566
rect 136161 162794 136541 163174
rect 136553 162794 136933 163174
rect 136945 162794 137325 163174
rect 137337 162794 137717 163174
rect 137729 162794 138109 163174
rect 138121 162794 138501 163174
rect 136161 162402 136541 162782
rect 136553 162402 136933 162782
rect 136945 162402 137325 162782
rect 137337 162402 137717 162782
rect 137729 162402 138109 162782
rect 138121 162402 138501 162782
rect 136161 162010 136541 162390
rect 136553 162010 136933 162390
rect 136945 162010 137325 162390
rect 137337 162010 137717 162390
rect 137729 162010 138109 162390
rect 138121 162010 138501 162390
rect 136161 161618 136541 161998
rect 136553 161618 136933 161998
rect 136945 161618 137325 161998
rect 137337 161618 137717 161998
rect 137729 161618 138109 161998
rect 138121 161618 138501 161998
rect 136161 161226 136541 161606
rect 136553 161226 136933 161606
rect 136945 161226 137325 161606
rect 137337 161226 137717 161606
rect 137729 161226 138109 161606
rect 138121 161226 138501 161606
rect 136161 160834 136541 161214
rect 136553 160834 136933 161214
rect 136945 160834 137325 161214
rect 137337 160834 137717 161214
rect 137729 160834 138109 161214
rect 138121 160834 138501 161214
rect 136161 160442 136541 160822
rect 136553 160442 136933 160822
rect 136945 160442 137325 160822
rect 137337 160442 137717 160822
rect 137729 160442 138109 160822
rect 138121 160442 138501 160822
rect 152161 163578 152541 163958
rect 152553 163578 152933 163958
rect 152945 163578 153325 163958
rect 153337 163578 153717 163958
rect 153729 163578 154109 163958
rect 154121 163578 154501 163958
rect 152161 163186 152541 163566
rect 152553 163186 152933 163566
rect 152945 163186 153325 163566
rect 153337 163186 153717 163566
rect 153729 163186 154109 163566
rect 154121 163186 154501 163566
rect 152161 162794 152541 163174
rect 152553 162794 152933 163174
rect 152945 162794 153325 163174
rect 153337 162794 153717 163174
rect 153729 162794 154109 163174
rect 154121 162794 154501 163174
rect 152161 162402 152541 162782
rect 152553 162402 152933 162782
rect 152945 162402 153325 162782
rect 153337 162402 153717 162782
rect 153729 162402 154109 162782
rect 154121 162402 154501 162782
rect 152161 162010 152541 162390
rect 152553 162010 152933 162390
rect 152945 162010 153325 162390
rect 153337 162010 153717 162390
rect 153729 162010 154109 162390
rect 154121 162010 154501 162390
rect 152161 161618 152541 161998
rect 152553 161618 152933 161998
rect 152945 161618 153325 161998
rect 153337 161618 153717 161998
rect 153729 161618 154109 161998
rect 154121 161618 154501 161998
rect 152161 161226 152541 161606
rect 152553 161226 152933 161606
rect 152945 161226 153325 161606
rect 153337 161226 153717 161606
rect 153729 161226 154109 161606
rect 154121 161226 154501 161606
rect 152161 160834 152541 161214
rect 152553 160834 152933 161214
rect 152945 160834 153325 161214
rect 153337 160834 153717 161214
rect 153729 160834 154109 161214
rect 154121 160834 154501 161214
rect 152161 160442 152541 160822
rect 152553 160442 152933 160822
rect 152945 160442 153325 160822
rect 153337 160442 153717 160822
rect 153729 160442 154109 160822
rect 154121 160442 154501 160822
rect 68430 154762 68810 155142
rect 68822 154762 69202 155142
rect 60042 154121 60422 154501
rect 60434 154121 60814 154501
rect 60826 154121 61206 154501
rect 61218 154121 61598 154501
rect 61610 154121 61990 154501
rect 62002 154121 62382 154501
rect 62394 154121 62774 154501
rect 62786 154121 63166 154501
rect 63178 154121 63558 154501
rect 60042 153729 60422 154109
rect 60434 153729 60814 154109
rect 60826 153729 61206 154109
rect 61218 153729 61598 154109
rect 61610 153729 61990 154109
rect 62002 153729 62382 154109
rect 62394 153729 62774 154109
rect 62786 153729 63166 154109
rect 63178 153729 63558 154109
rect 60042 153337 60422 153717
rect 60434 153337 60814 153717
rect 60826 153337 61206 153717
rect 61218 153337 61598 153717
rect 61610 153337 61990 153717
rect 62002 153337 62382 153717
rect 62394 153337 62774 153717
rect 62786 153337 63166 153717
rect 63178 153337 63558 153717
rect 60042 152945 60422 153325
rect 60434 152945 60814 153325
rect 60826 152945 61206 153325
rect 61218 152945 61598 153325
rect 61610 152945 61990 153325
rect 62002 152945 62382 153325
rect 62394 152945 62774 153325
rect 62786 152945 63166 153325
rect 63178 152945 63558 153325
rect 60042 152553 60422 152933
rect 60434 152553 60814 152933
rect 60826 152553 61206 152933
rect 61218 152553 61598 152933
rect 61610 152553 61990 152933
rect 62002 152553 62382 152933
rect 62394 152553 62774 152933
rect 62786 152553 63166 152933
rect 63178 152553 63558 152933
rect 60042 152161 60422 152541
rect 60434 152161 60814 152541
rect 60826 152161 61206 152541
rect 61218 152161 61598 152541
rect 61610 152161 61990 152541
rect 62002 152161 62382 152541
rect 62394 152161 62774 152541
rect 62786 152161 63166 152541
rect 63178 152161 63558 152541
rect 68430 154370 68810 154750
rect 68822 154370 69202 154750
rect 68430 151190 68810 151570
rect 68822 151190 69202 151570
rect 56042 148789 56422 149169
rect 56434 148789 56814 149169
rect 56826 148789 57206 149169
rect 57218 148789 57598 149169
rect 57610 148789 57990 149169
rect 58002 148789 58382 149169
rect 58394 148789 58774 149169
rect 58786 148789 59166 149169
rect 59178 148789 59558 149169
rect 56042 148397 56422 148777
rect 56434 148397 56814 148777
rect 56826 148397 57206 148777
rect 57218 148397 57598 148777
rect 57610 148397 57990 148777
rect 58002 148397 58382 148777
rect 58394 148397 58774 148777
rect 58786 148397 59166 148777
rect 59178 148397 59558 148777
rect 56042 148005 56422 148385
rect 56434 148005 56814 148385
rect 56826 148005 57206 148385
rect 57218 148005 57598 148385
rect 57610 148005 57990 148385
rect 58002 148005 58382 148385
rect 58394 148005 58774 148385
rect 58786 148005 59166 148385
rect 59178 148005 59558 148385
rect 56042 147613 56422 147993
rect 56434 147613 56814 147993
rect 56826 147613 57206 147993
rect 57218 147613 57598 147993
rect 57610 147613 57990 147993
rect 58002 147613 58382 147993
rect 58394 147613 58774 147993
rect 58786 147613 59166 147993
rect 59178 147613 59558 147993
rect 56042 147221 56422 147601
rect 56434 147221 56814 147601
rect 56826 147221 57206 147601
rect 57218 147221 57598 147601
rect 57610 147221 57990 147601
rect 58002 147221 58382 147601
rect 58394 147221 58774 147601
rect 58786 147221 59166 147601
rect 59178 147221 59558 147601
rect 56042 146829 56422 147209
rect 56434 146829 56814 147209
rect 56826 146829 57206 147209
rect 57218 146829 57598 147209
rect 57610 146829 57990 147209
rect 58002 146829 58382 147209
rect 58394 146829 58774 147209
rect 58786 146829 59166 147209
rect 59178 146829 59558 147209
rect 60042 138121 60422 138501
rect 60434 138121 60814 138501
rect 60826 138121 61206 138501
rect 61218 138121 61598 138501
rect 61610 138121 61990 138501
rect 62002 138121 62382 138501
rect 62394 138121 62774 138501
rect 62786 138121 63166 138501
rect 63178 138121 63558 138501
rect 60042 137729 60422 138109
rect 60434 137729 60814 138109
rect 60826 137729 61206 138109
rect 61218 137729 61598 138109
rect 61610 137729 61990 138109
rect 62002 137729 62382 138109
rect 62394 137729 62774 138109
rect 62786 137729 63166 138109
rect 63178 137729 63558 138109
rect 60042 137337 60422 137717
rect 60434 137337 60814 137717
rect 60826 137337 61206 137717
rect 61218 137337 61598 137717
rect 61610 137337 61990 137717
rect 62002 137337 62382 137717
rect 62394 137337 62774 137717
rect 62786 137337 63166 137717
rect 63178 137337 63558 137717
rect 60042 136945 60422 137325
rect 60434 136945 60814 137325
rect 60826 136945 61206 137325
rect 61218 136945 61598 137325
rect 61610 136945 61990 137325
rect 62002 136945 62382 137325
rect 62394 136945 62774 137325
rect 62786 136945 63166 137325
rect 63178 136945 63558 137325
rect 60042 136553 60422 136933
rect 60434 136553 60814 136933
rect 60826 136553 61206 136933
rect 61218 136553 61598 136933
rect 61610 136553 61990 136933
rect 62002 136553 62382 136933
rect 62394 136553 62774 136933
rect 62786 136553 63166 136933
rect 63178 136553 63558 136933
rect 60042 136161 60422 136541
rect 60434 136161 60814 136541
rect 60826 136161 61206 136541
rect 61218 136161 61598 136541
rect 61610 136161 61990 136541
rect 62002 136161 62382 136541
rect 62394 136161 62774 136541
rect 62786 136161 63166 136541
rect 63178 136161 63558 136541
rect 68430 138121 68810 138501
rect 68822 138121 69202 138501
rect 68430 137729 68810 138109
rect 68822 137729 69202 138109
rect 68430 137337 68810 137717
rect 68822 137337 69202 137717
rect 68430 136945 68810 137325
rect 68822 136945 69202 137325
rect 68430 136553 68810 136933
rect 68822 136553 69202 136933
rect 68430 136161 68810 136541
rect 68822 136161 69202 136541
rect 56042 132789 56422 133169
rect 56434 132789 56814 133169
rect 56826 132789 57206 133169
rect 57218 132789 57598 133169
rect 57610 132789 57990 133169
rect 58002 132789 58382 133169
rect 58394 132789 58774 133169
rect 58786 132789 59166 133169
rect 59178 132789 59558 133169
rect 56042 132397 56422 132777
rect 56434 132397 56814 132777
rect 56826 132397 57206 132777
rect 57218 132397 57598 132777
rect 57610 132397 57990 132777
rect 58002 132397 58382 132777
rect 58394 132397 58774 132777
rect 58786 132397 59166 132777
rect 59178 132397 59558 132777
rect 56042 132005 56422 132385
rect 56434 132005 56814 132385
rect 56826 132005 57206 132385
rect 57218 132005 57598 132385
rect 57610 132005 57990 132385
rect 58002 132005 58382 132385
rect 58394 132005 58774 132385
rect 58786 132005 59166 132385
rect 59178 132005 59558 132385
rect 56042 131613 56422 131993
rect 56434 131613 56814 131993
rect 56826 131613 57206 131993
rect 57218 131613 57598 131993
rect 57610 131613 57990 131993
rect 58002 131613 58382 131993
rect 58394 131613 58774 131993
rect 58786 131613 59166 131993
rect 59178 131613 59558 131993
rect 56042 131221 56422 131601
rect 56434 131221 56814 131601
rect 56826 131221 57206 131601
rect 57218 131221 57598 131601
rect 57610 131221 57990 131601
rect 58002 131221 58382 131601
rect 58394 131221 58774 131601
rect 58786 131221 59166 131601
rect 59178 131221 59558 131601
rect 56042 130829 56422 131209
rect 56434 130829 56814 131209
rect 56826 130829 57206 131209
rect 57218 130829 57598 131209
rect 57610 130829 57990 131209
rect 58002 130829 58382 131209
rect 58394 130829 58774 131209
rect 58786 130829 59166 131209
rect 59178 130829 59558 131209
rect 60042 122121 60422 122501
rect 60434 122121 60814 122501
rect 60826 122121 61206 122501
rect 61218 122121 61598 122501
rect 61610 122121 61990 122501
rect 62002 122121 62382 122501
rect 62394 122121 62774 122501
rect 62786 122121 63166 122501
rect 63178 122121 63558 122501
rect 60042 121729 60422 122109
rect 60434 121729 60814 122109
rect 60826 121729 61206 122109
rect 61218 121729 61598 122109
rect 61610 121729 61990 122109
rect 62002 121729 62382 122109
rect 62394 121729 62774 122109
rect 62786 121729 63166 122109
rect 63178 121729 63558 122109
rect 60042 121337 60422 121717
rect 60434 121337 60814 121717
rect 60826 121337 61206 121717
rect 61218 121337 61598 121717
rect 61610 121337 61990 121717
rect 62002 121337 62382 121717
rect 62394 121337 62774 121717
rect 62786 121337 63166 121717
rect 63178 121337 63558 121717
rect 60042 120945 60422 121325
rect 60434 120945 60814 121325
rect 60826 120945 61206 121325
rect 61218 120945 61598 121325
rect 61610 120945 61990 121325
rect 62002 120945 62382 121325
rect 62394 120945 62774 121325
rect 62786 120945 63166 121325
rect 63178 120945 63558 121325
rect 60042 120553 60422 120933
rect 60434 120553 60814 120933
rect 60826 120553 61206 120933
rect 61218 120553 61598 120933
rect 61610 120553 61990 120933
rect 62002 120553 62382 120933
rect 62394 120553 62774 120933
rect 62786 120553 63166 120933
rect 63178 120553 63558 120933
rect 60042 120161 60422 120541
rect 60434 120161 60814 120541
rect 60826 120161 61206 120541
rect 61218 120161 61598 120541
rect 61610 120161 61990 120541
rect 62002 120161 62382 120541
rect 62394 120161 62774 120541
rect 62786 120161 63166 120541
rect 63178 120161 63558 120541
rect 68430 122121 68810 122501
rect 68822 122121 69202 122501
rect 68430 121729 68810 122109
rect 68822 121729 69202 122109
rect 68430 121337 68810 121717
rect 68822 121337 69202 121717
rect 68430 120945 68810 121325
rect 68822 120945 69202 121325
rect 68430 120553 68810 120933
rect 68822 120553 69202 120933
rect 68430 120161 68810 120541
rect 68822 120161 69202 120541
rect 56042 116789 56422 117169
rect 56434 116789 56814 117169
rect 56826 116789 57206 117169
rect 57218 116789 57598 117169
rect 57610 116789 57990 117169
rect 58002 116789 58382 117169
rect 58394 116789 58774 117169
rect 58786 116789 59166 117169
rect 59178 116789 59558 117169
rect 56042 116397 56422 116777
rect 56434 116397 56814 116777
rect 56826 116397 57206 116777
rect 57218 116397 57598 116777
rect 57610 116397 57990 116777
rect 58002 116397 58382 116777
rect 58394 116397 58774 116777
rect 58786 116397 59166 116777
rect 59178 116397 59558 116777
rect 56042 116005 56422 116385
rect 56434 116005 56814 116385
rect 56826 116005 57206 116385
rect 57218 116005 57598 116385
rect 57610 116005 57990 116385
rect 58002 116005 58382 116385
rect 58394 116005 58774 116385
rect 58786 116005 59166 116385
rect 59178 116005 59558 116385
rect 56042 115613 56422 115993
rect 56434 115613 56814 115993
rect 56826 115613 57206 115993
rect 57218 115613 57598 115993
rect 57610 115613 57990 115993
rect 58002 115613 58382 115993
rect 58394 115613 58774 115993
rect 58786 115613 59166 115993
rect 59178 115613 59558 115993
rect 56042 115221 56422 115601
rect 56434 115221 56814 115601
rect 56826 115221 57206 115601
rect 57218 115221 57598 115601
rect 57610 115221 57990 115601
rect 58002 115221 58382 115601
rect 58394 115221 58774 115601
rect 58786 115221 59166 115601
rect 59178 115221 59558 115601
rect 56042 114829 56422 115209
rect 56434 114829 56814 115209
rect 56826 114829 57206 115209
rect 57218 114829 57598 115209
rect 57610 114829 57990 115209
rect 58002 114829 58382 115209
rect 58394 114829 58774 115209
rect 58786 114829 59166 115209
rect 59178 114829 59558 115209
rect 60042 106121 60422 106501
rect 60434 106121 60814 106501
rect 60826 106121 61206 106501
rect 61218 106121 61598 106501
rect 61610 106121 61990 106501
rect 62002 106121 62382 106501
rect 62394 106121 62774 106501
rect 62786 106121 63166 106501
rect 63178 106121 63558 106501
rect 60042 105729 60422 106109
rect 60434 105729 60814 106109
rect 60826 105729 61206 106109
rect 61218 105729 61598 106109
rect 61610 105729 61990 106109
rect 62002 105729 62382 106109
rect 62394 105729 62774 106109
rect 62786 105729 63166 106109
rect 63178 105729 63558 106109
rect 60042 105337 60422 105717
rect 60434 105337 60814 105717
rect 60826 105337 61206 105717
rect 61218 105337 61598 105717
rect 61610 105337 61990 105717
rect 62002 105337 62382 105717
rect 62394 105337 62774 105717
rect 62786 105337 63166 105717
rect 63178 105337 63558 105717
rect 60042 104945 60422 105325
rect 60434 104945 60814 105325
rect 60826 104945 61206 105325
rect 61218 104945 61598 105325
rect 61610 104945 61990 105325
rect 62002 104945 62382 105325
rect 62394 104945 62774 105325
rect 62786 104945 63166 105325
rect 63178 104945 63558 105325
rect 60042 104553 60422 104933
rect 60434 104553 60814 104933
rect 60826 104553 61206 104933
rect 61218 104553 61598 104933
rect 61610 104553 61990 104933
rect 62002 104553 62382 104933
rect 62394 104553 62774 104933
rect 62786 104553 63166 104933
rect 63178 104553 63558 104933
rect 60042 104161 60422 104541
rect 60434 104161 60814 104541
rect 60826 104161 61206 104541
rect 61218 104161 61598 104541
rect 61610 104161 61990 104541
rect 62002 104161 62382 104541
rect 62394 104161 62774 104541
rect 62786 104161 63166 104541
rect 63178 104161 63558 104541
rect 68430 106121 68810 106501
rect 68822 106121 69202 106501
rect 68430 105729 68810 106109
rect 68822 105729 69202 106109
rect 68430 105337 68810 105717
rect 68822 105337 69202 105717
rect 68430 104945 68810 105325
rect 68822 104945 69202 105325
rect 68430 104553 68810 104933
rect 68822 104553 69202 104933
rect 68430 104161 68810 104541
rect 68822 104161 69202 104541
rect 56042 100789 56422 101169
rect 56434 100789 56814 101169
rect 56826 100789 57206 101169
rect 57218 100789 57598 101169
rect 57610 100789 57990 101169
rect 58002 100789 58382 101169
rect 58394 100789 58774 101169
rect 58786 100789 59166 101169
rect 59178 100789 59558 101169
rect 56042 100397 56422 100777
rect 56434 100397 56814 100777
rect 56826 100397 57206 100777
rect 57218 100397 57598 100777
rect 57610 100397 57990 100777
rect 58002 100397 58382 100777
rect 58394 100397 58774 100777
rect 58786 100397 59166 100777
rect 59178 100397 59558 100777
rect 56042 100005 56422 100385
rect 56434 100005 56814 100385
rect 56826 100005 57206 100385
rect 57218 100005 57598 100385
rect 57610 100005 57990 100385
rect 58002 100005 58382 100385
rect 58394 100005 58774 100385
rect 58786 100005 59166 100385
rect 59178 100005 59558 100385
rect 56042 99613 56422 99993
rect 56434 99613 56814 99993
rect 56826 99613 57206 99993
rect 57218 99613 57598 99993
rect 57610 99613 57990 99993
rect 58002 99613 58382 99993
rect 58394 99613 58774 99993
rect 58786 99613 59166 99993
rect 59178 99613 59558 99993
rect 56042 99221 56422 99601
rect 56434 99221 56814 99601
rect 56826 99221 57206 99601
rect 57218 99221 57598 99601
rect 57610 99221 57990 99601
rect 58002 99221 58382 99601
rect 58394 99221 58774 99601
rect 58786 99221 59166 99601
rect 59178 99221 59558 99601
rect 56042 98829 56422 99209
rect 56434 98829 56814 99209
rect 56826 98829 57206 99209
rect 57218 98829 57598 99209
rect 57610 98829 57990 99209
rect 58002 98829 58382 99209
rect 58394 98829 58774 99209
rect 58786 98829 59166 99209
rect 59178 98829 59558 99209
rect 60042 90121 60422 90501
rect 60434 90121 60814 90501
rect 60826 90121 61206 90501
rect 61218 90121 61598 90501
rect 61610 90121 61990 90501
rect 62002 90121 62382 90501
rect 62394 90121 62774 90501
rect 62786 90121 63166 90501
rect 63178 90121 63558 90501
rect 60042 89729 60422 90109
rect 60434 89729 60814 90109
rect 60826 89729 61206 90109
rect 61218 89729 61598 90109
rect 61610 89729 61990 90109
rect 62002 89729 62382 90109
rect 62394 89729 62774 90109
rect 62786 89729 63166 90109
rect 63178 89729 63558 90109
rect 60042 89337 60422 89717
rect 60434 89337 60814 89717
rect 60826 89337 61206 89717
rect 61218 89337 61598 89717
rect 61610 89337 61990 89717
rect 62002 89337 62382 89717
rect 62394 89337 62774 89717
rect 62786 89337 63166 89717
rect 63178 89337 63558 89717
rect 60042 88945 60422 89325
rect 60434 88945 60814 89325
rect 60826 88945 61206 89325
rect 61218 88945 61598 89325
rect 61610 88945 61990 89325
rect 62002 88945 62382 89325
rect 62394 88945 62774 89325
rect 62786 88945 63166 89325
rect 63178 88945 63558 89325
rect 60042 88553 60422 88933
rect 60434 88553 60814 88933
rect 60826 88553 61206 88933
rect 61218 88553 61598 88933
rect 61610 88553 61990 88933
rect 62002 88553 62382 88933
rect 62394 88553 62774 88933
rect 62786 88553 63166 88933
rect 63178 88553 63558 88933
rect 60042 88161 60422 88541
rect 60434 88161 60814 88541
rect 60826 88161 61206 88541
rect 61218 88161 61598 88541
rect 61610 88161 61990 88541
rect 62002 88161 62382 88541
rect 62394 88161 62774 88541
rect 62786 88161 63166 88541
rect 63178 88161 63558 88541
rect 68430 90121 68810 90501
rect 68822 90121 69202 90501
rect 68430 89729 68810 90109
rect 68822 89729 69202 90109
rect 68430 89337 68810 89717
rect 68822 89337 69202 89717
rect 68430 88945 68810 89325
rect 68822 88945 69202 89325
rect 68430 88553 68810 88933
rect 68822 88553 69202 88933
rect 68430 88161 68810 88541
rect 68822 88161 69202 88541
rect 56042 84789 56422 85169
rect 56434 84789 56814 85169
rect 56826 84789 57206 85169
rect 57218 84789 57598 85169
rect 57610 84789 57990 85169
rect 58002 84789 58382 85169
rect 58394 84789 58774 85169
rect 58786 84789 59166 85169
rect 59178 84789 59558 85169
rect 56042 84397 56422 84777
rect 56434 84397 56814 84777
rect 56826 84397 57206 84777
rect 57218 84397 57598 84777
rect 57610 84397 57990 84777
rect 58002 84397 58382 84777
rect 58394 84397 58774 84777
rect 58786 84397 59166 84777
rect 59178 84397 59558 84777
rect 56042 84005 56422 84385
rect 56434 84005 56814 84385
rect 56826 84005 57206 84385
rect 57218 84005 57598 84385
rect 57610 84005 57990 84385
rect 58002 84005 58382 84385
rect 58394 84005 58774 84385
rect 58786 84005 59166 84385
rect 59178 84005 59558 84385
rect 56042 83613 56422 83993
rect 56434 83613 56814 83993
rect 56826 83613 57206 83993
rect 57218 83613 57598 83993
rect 57610 83613 57990 83993
rect 58002 83613 58382 83993
rect 58394 83613 58774 83993
rect 58786 83613 59166 83993
rect 59178 83613 59558 83993
rect 56042 83221 56422 83601
rect 56434 83221 56814 83601
rect 56826 83221 57206 83601
rect 57218 83221 57598 83601
rect 57610 83221 57990 83601
rect 58002 83221 58382 83601
rect 58394 83221 58774 83601
rect 58786 83221 59166 83601
rect 59178 83221 59558 83601
rect 56042 82829 56422 83209
rect 56434 82829 56814 83209
rect 56826 82829 57206 83209
rect 57218 82829 57598 83209
rect 57610 82829 57990 83209
rect 58002 82829 58382 83209
rect 58394 82829 58774 83209
rect 58786 82829 59166 83209
rect 59178 82829 59558 83209
rect 68430 75590 68810 75970
rect 68822 75590 69202 75970
rect 60042 74121 60422 74501
rect 60434 74121 60814 74501
rect 60826 74121 61206 74501
rect 61218 74121 61598 74501
rect 61610 74121 61990 74501
rect 62002 74121 62382 74501
rect 62394 74121 62774 74501
rect 62786 74121 63166 74501
rect 63178 74121 63558 74501
rect 60042 73729 60422 74109
rect 60434 73729 60814 74109
rect 60826 73729 61206 74109
rect 61218 73729 61598 74109
rect 61610 73729 61990 74109
rect 62002 73729 62382 74109
rect 62394 73729 62774 74109
rect 62786 73729 63166 74109
rect 63178 73729 63558 74109
rect 60042 73337 60422 73717
rect 60434 73337 60814 73717
rect 60826 73337 61206 73717
rect 61218 73337 61598 73717
rect 61610 73337 61990 73717
rect 62002 73337 62382 73717
rect 62394 73337 62774 73717
rect 62786 73337 63166 73717
rect 63178 73337 63558 73717
rect 60042 72945 60422 73325
rect 60434 72945 60814 73325
rect 60826 72945 61206 73325
rect 61218 72945 61598 73325
rect 61610 72945 61990 73325
rect 62002 72945 62382 73325
rect 62394 72945 62774 73325
rect 62786 72945 63166 73325
rect 63178 72945 63558 73325
rect 60042 72553 60422 72933
rect 60434 72553 60814 72933
rect 60826 72553 61206 72933
rect 61218 72553 61598 72933
rect 61610 72553 61990 72933
rect 62002 72553 62382 72933
rect 62394 72553 62774 72933
rect 62786 72553 63166 72933
rect 63178 72553 63558 72933
rect 60042 72161 60422 72541
rect 60434 72161 60814 72541
rect 60826 72161 61206 72541
rect 61218 72161 61598 72541
rect 61610 72161 61990 72541
rect 62002 72161 62382 72541
rect 62394 72161 62774 72541
rect 62786 72161 63166 72541
rect 63178 72161 63558 72541
rect 68430 74121 68810 74501
rect 68822 74121 69202 74501
rect 68430 73729 68810 74109
rect 68822 73729 69202 74109
rect 68430 73337 68810 73717
rect 68822 73337 69202 73717
rect 68430 72945 68810 73325
rect 68822 72945 69202 73325
rect 68430 72553 68810 72933
rect 68822 72553 69202 72933
rect 68430 72161 68810 72541
rect 68822 72161 69202 72541
rect 69830 153362 70210 153742
rect 70222 153362 70602 153742
rect 69830 152970 70210 153350
rect 70222 152970 70602 153350
rect 69830 148789 70210 149169
rect 70222 148789 70602 149169
rect 69830 148397 70210 148777
rect 70222 148397 70602 148777
rect 69830 148005 70210 148385
rect 70222 148005 70602 148385
rect 69830 147613 70210 147993
rect 70222 147613 70602 147993
rect 69830 147221 70210 147601
rect 70222 147221 70602 147601
rect 69830 146829 70210 147209
rect 70222 146829 70602 147209
rect 69830 134830 70210 135210
rect 70222 134830 70602 135210
rect 69830 132789 70210 133169
rect 70222 132789 70602 133169
rect 69830 132397 70210 132777
rect 70222 132397 70602 132777
rect 69830 132005 70210 132385
rect 70222 132005 70602 132385
rect 69830 131613 70210 131993
rect 70222 131613 70602 131993
rect 69830 131221 70210 131601
rect 70222 131221 70602 131601
rect 69830 130829 70210 131209
rect 70222 130829 70602 131209
rect 69830 119710 70210 120090
rect 70222 119710 70602 120090
rect 69830 116789 70210 117169
rect 70222 116789 70602 117169
rect 69830 116397 70210 116777
rect 70222 116397 70602 116777
rect 69830 116005 70210 116385
rect 70222 116005 70602 116385
rect 69830 115613 70210 115993
rect 70222 115613 70602 115993
rect 69830 115221 70210 115601
rect 70222 115221 70602 115601
rect 69830 114829 70210 115209
rect 70222 114829 70602 115209
rect 69830 104590 70210 104970
rect 70222 104590 70602 104970
rect 69830 100789 70210 101169
rect 70222 100789 70602 101169
rect 69830 100397 70210 100777
rect 70222 100397 70602 100777
rect 69830 100005 70210 100385
rect 70222 100005 70602 100385
rect 69830 99613 70210 99993
rect 70222 99613 70602 99993
rect 69830 99221 70210 99601
rect 70222 99221 70602 99601
rect 69830 98829 70210 99209
rect 70222 98829 70602 99209
rect 69830 89470 70210 89850
rect 70222 89470 70602 89850
rect 69830 84789 70210 85169
rect 70222 84789 70602 85169
rect 69830 84397 70210 84777
rect 70222 84397 70602 84777
rect 69830 84005 70210 84385
rect 70222 84005 70602 84385
rect 69830 83613 70210 83993
rect 70222 83613 70602 83993
rect 69830 83221 70210 83601
rect 70222 83221 70602 83601
rect 69830 82829 70210 83209
rect 70222 82829 70602 83209
rect 69830 74350 70210 74730
rect 70222 74350 70602 74730
rect 69830 70426 70210 70806
rect 70222 70426 70602 70806
rect 69830 70034 70210 70414
rect 70222 70034 70602 70414
rect 74146 153362 74526 153742
rect 74146 152970 74526 153350
rect 74146 149950 74526 150330
rect 74146 134830 74526 135210
rect 74146 119710 74526 120090
rect 74146 104590 74526 104970
rect 74146 89470 74526 89850
rect 74146 74350 74526 74730
rect 74146 70426 74526 70806
rect 74146 70034 74526 70414
rect 68430 69026 68810 69406
rect 68822 69026 69202 69406
rect 68430 68634 68810 69014
rect 68822 68634 69202 69014
rect 75386 154762 75766 155142
rect 75386 154370 75766 154750
rect 75386 151190 75766 151570
rect 75386 136070 75766 136450
rect 75386 120950 75766 121330
rect 75386 105830 75766 106210
rect 75386 90710 75766 91090
rect 75386 75590 75766 75970
rect 75386 69026 75766 69406
rect 75386 68634 75766 69014
rect 89266 153362 89646 153742
rect 89266 152970 89646 153350
rect 89266 149950 89646 150330
rect 89266 134830 89646 135210
rect 89266 119710 89646 120090
rect 89266 104590 89646 104970
rect 89266 89470 89646 89850
rect 89266 74350 89646 74730
rect 89266 70426 89646 70806
rect 89266 70034 89646 70414
rect 90506 154762 90886 155142
rect 90506 154370 90886 154750
rect 90506 151190 90886 151570
rect 90506 136070 90886 136450
rect 90506 120950 90886 121330
rect 90506 105830 90886 106210
rect 90506 90710 90886 91090
rect 90506 75590 90886 75970
rect 90506 69026 90886 69406
rect 90506 68634 90886 69014
rect 104386 153362 104766 153742
rect 104386 152970 104766 153350
rect 104386 149950 104766 150330
rect 104386 134830 104766 135210
rect 104386 119710 104766 120090
rect 104386 104590 104766 104970
rect 104386 89470 104766 89850
rect 104386 74350 104766 74730
rect 104386 70426 104766 70806
rect 104386 70034 104766 70414
rect 105626 154762 106006 155142
rect 105626 154370 106006 154750
rect 105626 151190 106006 151570
rect 105626 136070 106006 136450
rect 105626 120950 106006 121330
rect 105626 105830 106006 106210
rect 105626 90710 106006 91090
rect 105626 75590 106006 75970
rect 105626 69026 106006 69406
rect 105626 68634 106006 69014
rect 119506 153362 119886 153742
rect 119506 152970 119886 153350
rect 119506 149950 119886 150330
rect 119506 134830 119886 135210
rect 119506 119710 119886 120090
rect 119506 104590 119886 104970
rect 119506 89470 119886 89850
rect 119506 74350 119886 74730
rect 119506 70426 119886 70806
rect 119506 70034 119886 70414
rect 120746 154762 121126 155142
rect 120746 154370 121126 154750
rect 120746 151190 121126 151570
rect 120746 136070 121126 136450
rect 120746 120950 121126 121330
rect 120746 105830 121126 106210
rect 120746 90710 121126 91090
rect 120746 75590 121126 75970
rect 120746 69026 121126 69406
rect 120746 68634 121126 69014
rect 134626 153362 135006 153742
rect 134626 152970 135006 153350
rect 134626 149950 135006 150330
rect 134626 134830 135006 135210
rect 134626 119710 135006 120090
rect 134626 104590 135006 104970
rect 134626 89470 135006 89850
rect 134626 74350 135006 74730
rect 134626 70426 135006 70806
rect 134626 70034 135006 70414
rect 135866 154762 136246 155142
rect 135866 154370 136246 154750
rect 135866 151190 136246 151570
rect 135866 136070 136246 136450
rect 135866 120950 136246 121330
rect 135866 105830 136246 106210
rect 135866 90710 136246 91090
rect 135866 75590 136246 75970
rect 135866 69026 136246 69406
rect 135866 68634 136246 69014
rect 149746 153362 150126 153742
rect 149746 152970 150126 153350
rect 149746 149950 150126 150330
rect 149746 134830 150126 135210
rect 149746 119710 150126 120090
rect 149746 104590 150126 104970
rect 149746 89470 150126 89850
rect 149746 74350 150126 74730
rect 149746 70426 150126 70806
rect 149746 70034 150126 70414
rect 150986 154762 151366 155142
rect 150986 154370 151366 154750
rect 154766 154762 155146 155142
rect 155158 154762 155538 155142
rect 154766 154370 155146 154750
rect 155158 154370 155538 154750
rect 150986 151190 151366 151570
rect 150986 136070 151366 136450
rect 150986 120950 151366 121330
rect 150986 105830 151366 106210
rect 150986 90710 151366 91090
rect 150986 75590 151366 75970
rect 153366 153362 153746 153742
rect 153758 153362 154138 153742
rect 153366 152970 153746 153350
rect 153758 152970 154138 153350
rect 153366 148789 153746 149169
rect 153758 148789 154138 149169
rect 153366 148397 153746 148777
rect 153758 148397 154138 148777
rect 153366 148005 153746 148385
rect 153758 148005 154138 148385
rect 153366 147613 153746 147993
rect 153758 147613 154138 147993
rect 153366 147221 153746 147601
rect 153758 147221 154138 147601
rect 153366 146829 153746 147209
rect 153758 146829 154138 147209
rect 153366 134830 153746 135210
rect 153758 134830 154138 135210
rect 153366 132789 153746 133169
rect 153758 132789 154138 133169
rect 153366 132397 153746 132777
rect 153758 132397 154138 132777
rect 153366 132005 153746 132385
rect 153758 132005 154138 132385
rect 153366 131613 153746 131993
rect 153758 131613 154138 131993
rect 153366 131221 153746 131601
rect 153758 131221 154138 131601
rect 153366 130829 153746 131209
rect 153758 130829 154138 131209
rect 153366 119710 153746 120090
rect 153758 119710 154138 120090
rect 153366 116789 153746 117169
rect 153758 116789 154138 117169
rect 153366 116397 153746 116777
rect 153758 116397 154138 116777
rect 153366 116005 153746 116385
rect 153758 116005 154138 116385
rect 153366 115613 153746 115993
rect 153758 115613 154138 115993
rect 153366 115221 153746 115601
rect 153758 115221 154138 115601
rect 153366 114829 153746 115209
rect 153758 114829 154138 115209
rect 153366 104590 153746 104970
rect 153758 104590 154138 104970
rect 153366 100789 153746 101169
rect 153758 100789 154138 101169
rect 153366 100397 153746 100777
rect 153758 100397 154138 100777
rect 153366 100005 153746 100385
rect 153758 100005 154138 100385
rect 153366 99613 153746 99993
rect 153758 99613 154138 99993
rect 153366 99221 153746 99601
rect 153758 99221 154138 99601
rect 153366 98829 153746 99209
rect 153758 98829 154138 99209
rect 153366 89470 153746 89850
rect 153758 89470 154138 89850
rect 153366 84789 153746 85169
rect 153758 84789 154138 85169
rect 153366 84397 153746 84777
rect 153758 84397 154138 84777
rect 153366 84005 153746 84385
rect 153758 84005 154138 84385
rect 153366 83613 153746 83993
rect 153758 83613 154138 83993
rect 153366 83221 153746 83601
rect 153758 83221 154138 83601
rect 153366 82829 153746 83209
rect 153758 82829 154138 83209
rect 153366 74350 153746 74730
rect 153758 74350 154138 74730
rect 153366 70426 153746 70806
rect 153758 70426 154138 70806
rect 153366 70034 153746 70414
rect 153758 70034 154138 70414
rect 160442 154121 160822 154501
rect 160834 154121 161214 154501
rect 161226 154121 161606 154501
rect 161618 154121 161998 154501
rect 162010 154121 162390 154501
rect 162402 154121 162782 154501
rect 162794 154121 163174 154501
rect 163186 154121 163566 154501
rect 163578 154121 163958 154501
rect 160442 153729 160822 154109
rect 160834 153729 161214 154109
rect 161226 153729 161606 154109
rect 161618 153729 161998 154109
rect 162010 153729 162390 154109
rect 162402 153729 162782 154109
rect 162794 153729 163174 154109
rect 163186 153729 163566 154109
rect 163578 153729 163958 154109
rect 160442 153337 160822 153717
rect 160834 153337 161214 153717
rect 161226 153337 161606 153717
rect 161618 153337 161998 153717
rect 162010 153337 162390 153717
rect 162402 153337 162782 153717
rect 162794 153337 163174 153717
rect 163186 153337 163566 153717
rect 163578 153337 163958 153717
rect 160442 152945 160822 153325
rect 160834 152945 161214 153325
rect 161226 152945 161606 153325
rect 161618 152945 161998 153325
rect 162010 152945 162390 153325
rect 162402 152945 162782 153325
rect 162794 152945 163174 153325
rect 163186 152945 163566 153325
rect 163578 152945 163958 153325
rect 160442 152553 160822 152933
rect 160834 152553 161214 152933
rect 161226 152553 161606 152933
rect 161618 152553 161998 152933
rect 162010 152553 162390 152933
rect 162402 152553 162782 152933
rect 162794 152553 163174 152933
rect 163186 152553 163566 152933
rect 163578 152553 163958 152933
rect 160442 152161 160822 152541
rect 160834 152161 161214 152541
rect 161226 152161 161606 152541
rect 161618 152161 161998 152541
rect 162010 152161 162390 152541
rect 162402 152161 162782 152541
rect 162794 152161 163174 152541
rect 163186 152161 163566 152541
rect 163578 152161 163958 152541
rect 154766 151190 155146 151570
rect 155158 151190 155538 151570
rect 164442 148789 164822 149169
rect 164834 148789 165214 149169
rect 165226 148789 165606 149169
rect 165618 148789 165998 149169
rect 166010 148789 166390 149169
rect 166402 148789 166782 149169
rect 166794 148789 167174 149169
rect 167186 148789 167566 149169
rect 167578 148789 167958 149169
rect 164442 148397 164822 148777
rect 164834 148397 165214 148777
rect 165226 148397 165606 148777
rect 165618 148397 165998 148777
rect 166010 148397 166390 148777
rect 166402 148397 166782 148777
rect 166794 148397 167174 148777
rect 167186 148397 167566 148777
rect 167578 148397 167958 148777
rect 164442 148005 164822 148385
rect 164834 148005 165214 148385
rect 165226 148005 165606 148385
rect 165618 148005 165998 148385
rect 166010 148005 166390 148385
rect 166402 148005 166782 148385
rect 166794 148005 167174 148385
rect 167186 148005 167566 148385
rect 167578 148005 167958 148385
rect 164442 147613 164822 147993
rect 164834 147613 165214 147993
rect 165226 147613 165606 147993
rect 165618 147613 165998 147993
rect 166010 147613 166390 147993
rect 166402 147613 166782 147993
rect 166794 147613 167174 147993
rect 167186 147613 167566 147993
rect 167578 147613 167958 147993
rect 164442 147221 164822 147601
rect 164834 147221 165214 147601
rect 165226 147221 165606 147601
rect 165618 147221 165998 147601
rect 166010 147221 166390 147601
rect 166402 147221 166782 147601
rect 166794 147221 167174 147601
rect 167186 147221 167566 147601
rect 167578 147221 167958 147601
rect 164442 146829 164822 147209
rect 164834 146829 165214 147209
rect 165226 146829 165606 147209
rect 165618 146829 165998 147209
rect 166010 146829 166390 147209
rect 166402 146829 166782 147209
rect 166794 146829 167174 147209
rect 167186 146829 167566 147209
rect 167578 146829 167958 147209
rect 154766 138121 155146 138501
rect 155158 138121 155538 138501
rect 154766 137729 155146 138109
rect 155158 137729 155538 138109
rect 154766 137337 155146 137717
rect 155158 137337 155538 137717
rect 154766 136945 155146 137325
rect 155158 136945 155538 137325
rect 154766 136553 155146 136933
rect 155158 136553 155538 136933
rect 154766 136161 155146 136541
rect 155158 136161 155538 136541
rect 160442 138121 160822 138501
rect 160834 138121 161214 138501
rect 161226 138121 161606 138501
rect 161618 138121 161998 138501
rect 162010 138121 162390 138501
rect 162402 138121 162782 138501
rect 162794 138121 163174 138501
rect 163186 138121 163566 138501
rect 163578 138121 163958 138501
rect 160442 137729 160822 138109
rect 160834 137729 161214 138109
rect 161226 137729 161606 138109
rect 161618 137729 161998 138109
rect 162010 137729 162390 138109
rect 162402 137729 162782 138109
rect 162794 137729 163174 138109
rect 163186 137729 163566 138109
rect 163578 137729 163958 138109
rect 160442 137337 160822 137717
rect 160834 137337 161214 137717
rect 161226 137337 161606 137717
rect 161618 137337 161998 137717
rect 162010 137337 162390 137717
rect 162402 137337 162782 137717
rect 162794 137337 163174 137717
rect 163186 137337 163566 137717
rect 163578 137337 163958 137717
rect 160442 136945 160822 137325
rect 160834 136945 161214 137325
rect 161226 136945 161606 137325
rect 161618 136945 161998 137325
rect 162010 136945 162390 137325
rect 162402 136945 162782 137325
rect 162794 136945 163174 137325
rect 163186 136945 163566 137325
rect 163578 136945 163958 137325
rect 160442 136553 160822 136933
rect 160834 136553 161214 136933
rect 161226 136553 161606 136933
rect 161618 136553 161998 136933
rect 162010 136553 162390 136933
rect 162402 136553 162782 136933
rect 162794 136553 163174 136933
rect 163186 136553 163566 136933
rect 163578 136553 163958 136933
rect 160442 136161 160822 136541
rect 160834 136161 161214 136541
rect 161226 136161 161606 136541
rect 161618 136161 161998 136541
rect 162010 136161 162390 136541
rect 162402 136161 162782 136541
rect 162794 136161 163174 136541
rect 163186 136161 163566 136541
rect 163578 136161 163958 136541
rect 164442 132789 164822 133169
rect 164834 132789 165214 133169
rect 165226 132789 165606 133169
rect 165618 132789 165998 133169
rect 166010 132789 166390 133169
rect 166402 132789 166782 133169
rect 166794 132789 167174 133169
rect 167186 132789 167566 133169
rect 167578 132789 167958 133169
rect 164442 132397 164822 132777
rect 164834 132397 165214 132777
rect 165226 132397 165606 132777
rect 165618 132397 165998 132777
rect 166010 132397 166390 132777
rect 166402 132397 166782 132777
rect 166794 132397 167174 132777
rect 167186 132397 167566 132777
rect 167578 132397 167958 132777
rect 164442 132005 164822 132385
rect 164834 132005 165214 132385
rect 165226 132005 165606 132385
rect 165618 132005 165998 132385
rect 166010 132005 166390 132385
rect 166402 132005 166782 132385
rect 166794 132005 167174 132385
rect 167186 132005 167566 132385
rect 167578 132005 167958 132385
rect 164442 131613 164822 131993
rect 164834 131613 165214 131993
rect 165226 131613 165606 131993
rect 165618 131613 165998 131993
rect 166010 131613 166390 131993
rect 166402 131613 166782 131993
rect 166794 131613 167174 131993
rect 167186 131613 167566 131993
rect 167578 131613 167958 131993
rect 164442 131221 164822 131601
rect 164834 131221 165214 131601
rect 165226 131221 165606 131601
rect 165618 131221 165998 131601
rect 166010 131221 166390 131601
rect 166402 131221 166782 131601
rect 166794 131221 167174 131601
rect 167186 131221 167566 131601
rect 167578 131221 167958 131601
rect 164442 130829 164822 131209
rect 164834 130829 165214 131209
rect 165226 130829 165606 131209
rect 165618 130829 165998 131209
rect 166010 130829 166390 131209
rect 166402 130829 166782 131209
rect 166794 130829 167174 131209
rect 167186 130829 167566 131209
rect 167578 130829 167958 131209
rect 154766 122121 155146 122501
rect 155158 122121 155538 122501
rect 154766 121729 155146 122109
rect 155158 121729 155538 122109
rect 154766 121337 155146 121717
rect 155158 121337 155538 121717
rect 154766 120945 155146 121325
rect 155158 120945 155538 121325
rect 154766 120553 155146 120933
rect 155158 120553 155538 120933
rect 154766 120161 155146 120541
rect 155158 120161 155538 120541
rect 160442 122121 160822 122501
rect 160834 122121 161214 122501
rect 161226 122121 161606 122501
rect 161618 122121 161998 122501
rect 162010 122121 162390 122501
rect 162402 122121 162782 122501
rect 162794 122121 163174 122501
rect 163186 122121 163566 122501
rect 163578 122121 163958 122501
rect 160442 121729 160822 122109
rect 160834 121729 161214 122109
rect 161226 121729 161606 122109
rect 161618 121729 161998 122109
rect 162010 121729 162390 122109
rect 162402 121729 162782 122109
rect 162794 121729 163174 122109
rect 163186 121729 163566 122109
rect 163578 121729 163958 122109
rect 160442 121337 160822 121717
rect 160834 121337 161214 121717
rect 161226 121337 161606 121717
rect 161618 121337 161998 121717
rect 162010 121337 162390 121717
rect 162402 121337 162782 121717
rect 162794 121337 163174 121717
rect 163186 121337 163566 121717
rect 163578 121337 163958 121717
rect 160442 120945 160822 121325
rect 160834 120945 161214 121325
rect 161226 120945 161606 121325
rect 161618 120945 161998 121325
rect 162010 120945 162390 121325
rect 162402 120945 162782 121325
rect 162794 120945 163174 121325
rect 163186 120945 163566 121325
rect 163578 120945 163958 121325
rect 160442 120553 160822 120933
rect 160834 120553 161214 120933
rect 161226 120553 161606 120933
rect 161618 120553 161998 120933
rect 162010 120553 162390 120933
rect 162402 120553 162782 120933
rect 162794 120553 163174 120933
rect 163186 120553 163566 120933
rect 163578 120553 163958 120933
rect 160442 120161 160822 120541
rect 160834 120161 161214 120541
rect 161226 120161 161606 120541
rect 161618 120161 161998 120541
rect 162010 120161 162390 120541
rect 162402 120161 162782 120541
rect 162794 120161 163174 120541
rect 163186 120161 163566 120541
rect 163578 120161 163958 120541
rect 164442 116789 164822 117169
rect 164834 116789 165214 117169
rect 165226 116789 165606 117169
rect 165618 116789 165998 117169
rect 166010 116789 166390 117169
rect 166402 116789 166782 117169
rect 166794 116789 167174 117169
rect 167186 116789 167566 117169
rect 167578 116789 167958 117169
rect 164442 116397 164822 116777
rect 164834 116397 165214 116777
rect 165226 116397 165606 116777
rect 165618 116397 165998 116777
rect 166010 116397 166390 116777
rect 166402 116397 166782 116777
rect 166794 116397 167174 116777
rect 167186 116397 167566 116777
rect 167578 116397 167958 116777
rect 164442 116005 164822 116385
rect 164834 116005 165214 116385
rect 165226 116005 165606 116385
rect 165618 116005 165998 116385
rect 166010 116005 166390 116385
rect 166402 116005 166782 116385
rect 166794 116005 167174 116385
rect 167186 116005 167566 116385
rect 167578 116005 167958 116385
rect 164442 115613 164822 115993
rect 164834 115613 165214 115993
rect 165226 115613 165606 115993
rect 165618 115613 165998 115993
rect 166010 115613 166390 115993
rect 166402 115613 166782 115993
rect 166794 115613 167174 115993
rect 167186 115613 167566 115993
rect 167578 115613 167958 115993
rect 164442 115221 164822 115601
rect 164834 115221 165214 115601
rect 165226 115221 165606 115601
rect 165618 115221 165998 115601
rect 166010 115221 166390 115601
rect 166402 115221 166782 115601
rect 166794 115221 167174 115601
rect 167186 115221 167566 115601
rect 167578 115221 167958 115601
rect 164442 114829 164822 115209
rect 164834 114829 165214 115209
rect 165226 114829 165606 115209
rect 165618 114829 165998 115209
rect 166010 114829 166390 115209
rect 166402 114829 166782 115209
rect 166794 114829 167174 115209
rect 167186 114829 167566 115209
rect 167578 114829 167958 115209
rect 154766 106121 155146 106501
rect 155158 106121 155538 106501
rect 154766 105729 155146 106109
rect 155158 105729 155538 106109
rect 154766 105337 155146 105717
rect 155158 105337 155538 105717
rect 154766 104945 155146 105325
rect 155158 104945 155538 105325
rect 154766 104553 155146 104933
rect 155158 104553 155538 104933
rect 154766 104161 155146 104541
rect 155158 104161 155538 104541
rect 160442 106121 160822 106501
rect 160834 106121 161214 106501
rect 161226 106121 161606 106501
rect 161618 106121 161998 106501
rect 162010 106121 162390 106501
rect 162402 106121 162782 106501
rect 162794 106121 163174 106501
rect 163186 106121 163566 106501
rect 163578 106121 163958 106501
rect 160442 105729 160822 106109
rect 160834 105729 161214 106109
rect 161226 105729 161606 106109
rect 161618 105729 161998 106109
rect 162010 105729 162390 106109
rect 162402 105729 162782 106109
rect 162794 105729 163174 106109
rect 163186 105729 163566 106109
rect 163578 105729 163958 106109
rect 160442 105337 160822 105717
rect 160834 105337 161214 105717
rect 161226 105337 161606 105717
rect 161618 105337 161998 105717
rect 162010 105337 162390 105717
rect 162402 105337 162782 105717
rect 162794 105337 163174 105717
rect 163186 105337 163566 105717
rect 163578 105337 163958 105717
rect 160442 104945 160822 105325
rect 160834 104945 161214 105325
rect 161226 104945 161606 105325
rect 161618 104945 161998 105325
rect 162010 104945 162390 105325
rect 162402 104945 162782 105325
rect 162794 104945 163174 105325
rect 163186 104945 163566 105325
rect 163578 104945 163958 105325
rect 160442 104553 160822 104933
rect 160834 104553 161214 104933
rect 161226 104553 161606 104933
rect 161618 104553 161998 104933
rect 162010 104553 162390 104933
rect 162402 104553 162782 104933
rect 162794 104553 163174 104933
rect 163186 104553 163566 104933
rect 163578 104553 163958 104933
rect 160442 104161 160822 104541
rect 160834 104161 161214 104541
rect 161226 104161 161606 104541
rect 161618 104161 161998 104541
rect 162010 104161 162390 104541
rect 162402 104161 162782 104541
rect 162794 104161 163174 104541
rect 163186 104161 163566 104541
rect 163578 104161 163958 104541
rect 164442 100789 164822 101169
rect 164834 100789 165214 101169
rect 165226 100789 165606 101169
rect 165618 100789 165998 101169
rect 166010 100789 166390 101169
rect 166402 100789 166782 101169
rect 166794 100789 167174 101169
rect 167186 100789 167566 101169
rect 167578 100789 167958 101169
rect 164442 100397 164822 100777
rect 164834 100397 165214 100777
rect 165226 100397 165606 100777
rect 165618 100397 165998 100777
rect 166010 100397 166390 100777
rect 166402 100397 166782 100777
rect 166794 100397 167174 100777
rect 167186 100397 167566 100777
rect 167578 100397 167958 100777
rect 164442 100005 164822 100385
rect 164834 100005 165214 100385
rect 165226 100005 165606 100385
rect 165618 100005 165998 100385
rect 166010 100005 166390 100385
rect 166402 100005 166782 100385
rect 166794 100005 167174 100385
rect 167186 100005 167566 100385
rect 167578 100005 167958 100385
rect 164442 99613 164822 99993
rect 164834 99613 165214 99993
rect 165226 99613 165606 99993
rect 165618 99613 165998 99993
rect 166010 99613 166390 99993
rect 166402 99613 166782 99993
rect 166794 99613 167174 99993
rect 167186 99613 167566 99993
rect 167578 99613 167958 99993
rect 164442 99221 164822 99601
rect 164834 99221 165214 99601
rect 165226 99221 165606 99601
rect 165618 99221 165998 99601
rect 166010 99221 166390 99601
rect 166402 99221 166782 99601
rect 166794 99221 167174 99601
rect 167186 99221 167566 99601
rect 167578 99221 167958 99601
rect 164442 98829 164822 99209
rect 164834 98829 165214 99209
rect 165226 98829 165606 99209
rect 165618 98829 165998 99209
rect 166010 98829 166390 99209
rect 166402 98829 166782 99209
rect 166794 98829 167174 99209
rect 167186 98829 167566 99209
rect 167578 98829 167958 99209
rect 154766 90121 155146 90501
rect 155158 90121 155538 90501
rect 154766 89729 155146 90109
rect 155158 89729 155538 90109
rect 154766 89337 155146 89717
rect 155158 89337 155538 89717
rect 154766 88945 155146 89325
rect 155158 88945 155538 89325
rect 154766 88553 155146 88933
rect 155158 88553 155538 88933
rect 154766 88161 155146 88541
rect 155158 88161 155538 88541
rect 160442 90121 160822 90501
rect 160834 90121 161214 90501
rect 161226 90121 161606 90501
rect 161618 90121 161998 90501
rect 162010 90121 162390 90501
rect 162402 90121 162782 90501
rect 162794 90121 163174 90501
rect 163186 90121 163566 90501
rect 163578 90121 163958 90501
rect 160442 89729 160822 90109
rect 160834 89729 161214 90109
rect 161226 89729 161606 90109
rect 161618 89729 161998 90109
rect 162010 89729 162390 90109
rect 162402 89729 162782 90109
rect 162794 89729 163174 90109
rect 163186 89729 163566 90109
rect 163578 89729 163958 90109
rect 160442 89337 160822 89717
rect 160834 89337 161214 89717
rect 161226 89337 161606 89717
rect 161618 89337 161998 89717
rect 162010 89337 162390 89717
rect 162402 89337 162782 89717
rect 162794 89337 163174 89717
rect 163186 89337 163566 89717
rect 163578 89337 163958 89717
rect 160442 88945 160822 89325
rect 160834 88945 161214 89325
rect 161226 88945 161606 89325
rect 161618 88945 161998 89325
rect 162010 88945 162390 89325
rect 162402 88945 162782 89325
rect 162794 88945 163174 89325
rect 163186 88945 163566 89325
rect 163578 88945 163958 89325
rect 160442 88553 160822 88933
rect 160834 88553 161214 88933
rect 161226 88553 161606 88933
rect 161618 88553 161998 88933
rect 162010 88553 162390 88933
rect 162402 88553 162782 88933
rect 162794 88553 163174 88933
rect 163186 88553 163566 88933
rect 163578 88553 163958 88933
rect 160442 88161 160822 88541
rect 160834 88161 161214 88541
rect 161226 88161 161606 88541
rect 161618 88161 161998 88541
rect 162010 88161 162390 88541
rect 162402 88161 162782 88541
rect 162794 88161 163174 88541
rect 163186 88161 163566 88541
rect 163578 88161 163958 88541
rect 164442 84789 164822 85169
rect 164834 84789 165214 85169
rect 165226 84789 165606 85169
rect 165618 84789 165998 85169
rect 166010 84789 166390 85169
rect 166402 84789 166782 85169
rect 166794 84789 167174 85169
rect 167186 84789 167566 85169
rect 167578 84789 167958 85169
rect 164442 84397 164822 84777
rect 164834 84397 165214 84777
rect 165226 84397 165606 84777
rect 165618 84397 165998 84777
rect 166010 84397 166390 84777
rect 166402 84397 166782 84777
rect 166794 84397 167174 84777
rect 167186 84397 167566 84777
rect 167578 84397 167958 84777
rect 164442 84005 164822 84385
rect 164834 84005 165214 84385
rect 165226 84005 165606 84385
rect 165618 84005 165998 84385
rect 166010 84005 166390 84385
rect 166402 84005 166782 84385
rect 166794 84005 167174 84385
rect 167186 84005 167566 84385
rect 167578 84005 167958 84385
rect 164442 83613 164822 83993
rect 164834 83613 165214 83993
rect 165226 83613 165606 83993
rect 165618 83613 165998 83993
rect 166010 83613 166390 83993
rect 166402 83613 166782 83993
rect 166794 83613 167174 83993
rect 167186 83613 167566 83993
rect 167578 83613 167958 83993
rect 164442 83221 164822 83601
rect 164834 83221 165214 83601
rect 165226 83221 165606 83601
rect 165618 83221 165998 83601
rect 166010 83221 166390 83601
rect 166402 83221 166782 83601
rect 166794 83221 167174 83601
rect 167186 83221 167566 83601
rect 167578 83221 167958 83601
rect 164442 82829 164822 83209
rect 164834 82829 165214 83209
rect 165226 82829 165606 83209
rect 165618 82829 165998 83209
rect 166010 82829 166390 83209
rect 166402 82829 166782 83209
rect 166794 82829 167174 83209
rect 167186 82829 167566 83209
rect 167578 82829 167958 83209
rect 154766 75590 155146 75970
rect 155158 75590 155538 75970
rect 154766 74121 155146 74501
rect 155158 74121 155538 74501
rect 154766 73729 155146 74109
rect 155158 73729 155538 74109
rect 154766 73337 155146 73717
rect 155158 73337 155538 73717
rect 154766 72945 155146 73325
rect 155158 72945 155538 73325
rect 154766 72553 155146 72933
rect 155158 72553 155538 72933
rect 154766 72161 155146 72541
rect 155158 72161 155538 72541
rect 150986 69026 151366 69406
rect 150986 68634 151366 69014
rect 160442 74121 160822 74501
rect 160834 74121 161214 74501
rect 161226 74121 161606 74501
rect 161618 74121 161998 74501
rect 162010 74121 162390 74501
rect 162402 74121 162782 74501
rect 162794 74121 163174 74501
rect 163186 74121 163566 74501
rect 163578 74121 163958 74501
rect 160442 73729 160822 74109
rect 160834 73729 161214 74109
rect 161226 73729 161606 74109
rect 161618 73729 161998 74109
rect 162010 73729 162390 74109
rect 162402 73729 162782 74109
rect 162794 73729 163174 74109
rect 163186 73729 163566 74109
rect 163578 73729 163958 74109
rect 160442 73337 160822 73717
rect 160834 73337 161214 73717
rect 161226 73337 161606 73717
rect 161618 73337 161998 73717
rect 162010 73337 162390 73717
rect 162402 73337 162782 73717
rect 162794 73337 163174 73717
rect 163186 73337 163566 73717
rect 163578 73337 163958 73717
rect 160442 72945 160822 73325
rect 160834 72945 161214 73325
rect 161226 72945 161606 73325
rect 161618 72945 161998 73325
rect 162010 72945 162390 73325
rect 162402 72945 162782 73325
rect 162794 72945 163174 73325
rect 163186 72945 163566 73325
rect 163578 72945 163958 73325
rect 160442 72553 160822 72933
rect 160834 72553 161214 72933
rect 161226 72553 161606 72933
rect 161618 72553 161998 72933
rect 162010 72553 162390 72933
rect 162402 72553 162782 72933
rect 162794 72553 163174 72933
rect 163186 72553 163566 72933
rect 163578 72553 163958 72933
rect 160442 72161 160822 72541
rect 160834 72161 161214 72541
rect 161226 72161 161606 72541
rect 161618 72161 161998 72541
rect 162010 72161 162390 72541
rect 162402 72161 162782 72541
rect 162794 72161 163174 72541
rect 163186 72161 163566 72541
rect 163578 72161 163958 72541
rect 154766 69026 155146 69406
rect 155158 69026 155538 69406
rect 154766 68634 155146 69014
rect 155158 68634 155538 69014
rect 72161 63178 72541 63558
rect 72553 63178 72933 63558
rect 72945 63178 73325 63558
rect 73337 63178 73717 63558
rect 73729 63178 74109 63558
rect 74121 63178 74501 63558
rect 72161 62786 72541 63166
rect 72553 62786 72933 63166
rect 72945 62786 73325 63166
rect 73337 62786 73717 63166
rect 73729 62786 74109 63166
rect 74121 62786 74501 63166
rect 72161 62394 72541 62774
rect 72553 62394 72933 62774
rect 72945 62394 73325 62774
rect 73337 62394 73717 62774
rect 73729 62394 74109 62774
rect 74121 62394 74501 62774
rect 72161 62002 72541 62382
rect 72553 62002 72933 62382
rect 72945 62002 73325 62382
rect 73337 62002 73717 62382
rect 73729 62002 74109 62382
rect 74121 62002 74501 62382
rect 72161 61610 72541 61990
rect 72553 61610 72933 61990
rect 72945 61610 73325 61990
rect 73337 61610 73717 61990
rect 73729 61610 74109 61990
rect 74121 61610 74501 61990
rect 72161 61218 72541 61598
rect 72553 61218 72933 61598
rect 72945 61218 73325 61598
rect 73337 61218 73717 61598
rect 73729 61218 74109 61598
rect 74121 61218 74501 61598
rect 72161 60826 72541 61206
rect 72553 60826 72933 61206
rect 72945 60826 73325 61206
rect 73337 60826 73717 61206
rect 73729 60826 74109 61206
rect 74121 60826 74501 61206
rect 72161 60434 72541 60814
rect 72553 60434 72933 60814
rect 72945 60434 73325 60814
rect 73337 60434 73717 60814
rect 73729 60434 74109 60814
rect 74121 60434 74501 60814
rect 72161 60042 72541 60422
rect 72553 60042 72933 60422
rect 72945 60042 73325 60422
rect 73337 60042 73717 60422
rect 73729 60042 74109 60422
rect 74121 60042 74501 60422
rect 88161 63178 88541 63558
rect 88553 63178 88933 63558
rect 88945 63178 89325 63558
rect 89337 63178 89717 63558
rect 89729 63178 90109 63558
rect 90121 63178 90501 63558
rect 88161 62786 88541 63166
rect 88553 62786 88933 63166
rect 88945 62786 89325 63166
rect 89337 62786 89717 63166
rect 89729 62786 90109 63166
rect 90121 62786 90501 63166
rect 88161 62394 88541 62774
rect 88553 62394 88933 62774
rect 88945 62394 89325 62774
rect 89337 62394 89717 62774
rect 89729 62394 90109 62774
rect 90121 62394 90501 62774
rect 88161 62002 88541 62382
rect 88553 62002 88933 62382
rect 88945 62002 89325 62382
rect 89337 62002 89717 62382
rect 89729 62002 90109 62382
rect 90121 62002 90501 62382
rect 88161 61610 88541 61990
rect 88553 61610 88933 61990
rect 88945 61610 89325 61990
rect 89337 61610 89717 61990
rect 89729 61610 90109 61990
rect 90121 61610 90501 61990
rect 88161 61218 88541 61598
rect 88553 61218 88933 61598
rect 88945 61218 89325 61598
rect 89337 61218 89717 61598
rect 89729 61218 90109 61598
rect 90121 61218 90501 61598
rect 88161 60826 88541 61206
rect 88553 60826 88933 61206
rect 88945 60826 89325 61206
rect 89337 60826 89717 61206
rect 89729 60826 90109 61206
rect 90121 60826 90501 61206
rect 88161 60434 88541 60814
rect 88553 60434 88933 60814
rect 88945 60434 89325 60814
rect 89337 60434 89717 60814
rect 89729 60434 90109 60814
rect 90121 60434 90501 60814
rect 88161 60042 88541 60422
rect 88553 60042 88933 60422
rect 88945 60042 89325 60422
rect 89337 60042 89717 60422
rect 89729 60042 90109 60422
rect 90121 60042 90501 60422
rect 104161 63178 104541 63558
rect 104553 63178 104933 63558
rect 104945 63178 105325 63558
rect 105337 63178 105717 63558
rect 105729 63178 106109 63558
rect 106121 63178 106501 63558
rect 104161 62786 104541 63166
rect 104553 62786 104933 63166
rect 104945 62786 105325 63166
rect 105337 62786 105717 63166
rect 105729 62786 106109 63166
rect 106121 62786 106501 63166
rect 104161 62394 104541 62774
rect 104553 62394 104933 62774
rect 104945 62394 105325 62774
rect 105337 62394 105717 62774
rect 105729 62394 106109 62774
rect 106121 62394 106501 62774
rect 104161 62002 104541 62382
rect 104553 62002 104933 62382
rect 104945 62002 105325 62382
rect 105337 62002 105717 62382
rect 105729 62002 106109 62382
rect 106121 62002 106501 62382
rect 104161 61610 104541 61990
rect 104553 61610 104933 61990
rect 104945 61610 105325 61990
rect 105337 61610 105717 61990
rect 105729 61610 106109 61990
rect 106121 61610 106501 61990
rect 104161 61218 104541 61598
rect 104553 61218 104933 61598
rect 104945 61218 105325 61598
rect 105337 61218 105717 61598
rect 105729 61218 106109 61598
rect 106121 61218 106501 61598
rect 104161 60826 104541 61206
rect 104553 60826 104933 61206
rect 104945 60826 105325 61206
rect 105337 60826 105717 61206
rect 105729 60826 106109 61206
rect 106121 60826 106501 61206
rect 104161 60434 104541 60814
rect 104553 60434 104933 60814
rect 104945 60434 105325 60814
rect 105337 60434 105717 60814
rect 105729 60434 106109 60814
rect 106121 60434 106501 60814
rect 104161 60042 104541 60422
rect 104553 60042 104933 60422
rect 104945 60042 105325 60422
rect 105337 60042 105717 60422
rect 105729 60042 106109 60422
rect 106121 60042 106501 60422
rect 120161 63178 120541 63558
rect 120553 63178 120933 63558
rect 120945 63178 121325 63558
rect 121337 63178 121717 63558
rect 121729 63178 122109 63558
rect 122121 63178 122501 63558
rect 120161 62786 120541 63166
rect 120553 62786 120933 63166
rect 120945 62786 121325 63166
rect 121337 62786 121717 63166
rect 121729 62786 122109 63166
rect 122121 62786 122501 63166
rect 120161 62394 120541 62774
rect 120553 62394 120933 62774
rect 120945 62394 121325 62774
rect 121337 62394 121717 62774
rect 121729 62394 122109 62774
rect 122121 62394 122501 62774
rect 120161 62002 120541 62382
rect 120553 62002 120933 62382
rect 120945 62002 121325 62382
rect 121337 62002 121717 62382
rect 121729 62002 122109 62382
rect 122121 62002 122501 62382
rect 120161 61610 120541 61990
rect 120553 61610 120933 61990
rect 120945 61610 121325 61990
rect 121337 61610 121717 61990
rect 121729 61610 122109 61990
rect 122121 61610 122501 61990
rect 120161 61218 120541 61598
rect 120553 61218 120933 61598
rect 120945 61218 121325 61598
rect 121337 61218 121717 61598
rect 121729 61218 122109 61598
rect 122121 61218 122501 61598
rect 120161 60826 120541 61206
rect 120553 60826 120933 61206
rect 120945 60826 121325 61206
rect 121337 60826 121717 61206
rect 121729 60826 122109 61206
rect 122121 60826 122501 61206
rect 120161 60434 120541 60814
rect 120553 60434 120933 60814
rect 120945 60434 121325 60814
rect 121337 60434 121717 60814
rect 121729 60434 122109 60814
rect 122121 60434 122501 60814
rect 120161 60042 120541 60422
rect 120553 60042 120933 60422
rect 120945 60042 121325 60422
rect 121337 60042 121717 60422
rect 121729 60042 122109 60422
rect 122121 60042 122501 60422
rect 132046 63178 132426 63558
rect 132438 63178 132818 63558
rect 132830 63178 133210 63558
rect 133222 63178 133602 63558
rect 133614 63178 133994 63558
rect 134006 63178 134386 63558
rect 134398 63178 134778 63558
rect 134790 63178 135170 63558
rect 135182 63178 135562 63558
rect 135574 63178 135954 63558
rect 132046 62786 132426 63166
rect 132438 62786 132818 63166
rect 132830 62786 133210 63166
rect 133222 62786 133602 63166
rect 133614 62786 133994 63166
rect 134006 62786 134386 63166
rect 134398 62786 134778 63166
rect 134790 62786 135170 63166
rect 135182 62786 135562 63166
rect 135574 62786 135954 63166
rect 132046 62394 132426 62774
rect 132438 62394 132818 62774
rect 132830 62394 133210 62774
rect 133222 62394 133602 62774
rect 133614 62394 133994 62774
rect 134006 62394 134386 62774
rect 134398 62394 134778 62774
rect 134790 62394 135170 62774
rect 135182 62394 135562 62774
rect 135574 62394 135954 62774
rect 132046 62002 132426 62382
rect 132438 62002 132818 62382
rect 132830 62002 133210 62382
rect 133222 62002 133602 62382
rect 133614 62002 133994 62382
rect 134006 62002 134386 62382
rect 134398 62002 134778 62382
rect 134790 62002 135170 62382
rect 135182 62002 135562 62382
rect 135574 62002 135954 62382
rect 132046 61610 132426 61990
rect 132438 61610 132818 61990
rect 132830 61610 133210 61990
rect 133222 61610 133602 61990
rect 133614 61610 133994 61990
rect 134006 61610 134386 61990
rect 134398 61610 134778 61990
rect 134790 61610 135170 61990
rect 135182 61610 135562 61990
rect 135574 61610 135954 61990
rect 132046 61218 132426 61598
rect 132438 61218 132818 61598
rect 132830 61218 133210 61598
rect 133222 61218 133602 61598
rect 133614 61218 133994 61598
rect 134006 61218 134386 61598
rect 134398 61218 134778 61598
rect 134790 61218 135170 61598
rect 135182 61218 135562 61598
rect 135574 61218 135954 61598
rect 132046 60826 132426 61206
rect 132438 60826 132818 61206
rect 132830 60826 133210 61206
rect 133222 60826 133602 61206
rect 133614 60826 133994 61206
rect 134006 60826 134386 61206
rect 134398 60826 134778 61206
rect 134790 60826 135170 61206
rect 135182 60826 135562 61206
rect 135574 60826 135954 61206
rect 132046 60434 132426 60814
rect 132438 60434 132818 60814
rect 132830 60434 133210 60814
rect 133222 60434 133602 60814
rect 133614 60434 133994 60814
rect 134006 60434 134386 60814
rect 134398 60434 134778 60814
rect 134790 60434 135170 60814
rect 135182 60434 135562 60814
rect 135574 60434 135954 60814
rect 132046 60042 132426 60422
rect 132438 60042 132818 60422
rect 132830 60042 133210 60422
rect 133222 60042 133602 60422
rect 133614 60042 133994 60422
rect 134006 60042 134386 60422
rect 134398 60042 134778 60422
rect 134790 60042 135170 60422
rect 135182 60042 135562 60422
rect 135574 60042 135954 60422
rect 152161 63178 152541 63558
rect 152553 63178 152933 63558
rect 152945 63178 153325 63558
rect 153337 63178 153717 63558
rect 153729 63178 154109 63558
rect 154121 63178 154501 63558
rect 152161 62786 152541 63166
rect 152553 62786 152933 63166
rect 152945 62786 153325 63166
rect 153337 62786 153717 63166
rect 153729 62786 154109 63166
rect 154121 62786 154501 63166
rect 152161 62394 152541 62774
rect 152553 62394 152933 62774
rect 152945 62394 153325 62774
rect 153337 62394 153717 62774
rect 153729 62394 154109 62774
rect 154121 62394 154501 62774
rect 152161 62002 152541 62382
rect 152553 62002 152933 62382
rect 152945 62002 153325 62382
rect 153337 62002 153717 62382
rect 153729 62002 154109 62382
rect 154121 62002 154501 62382
rect 152161 61610 152541 61990
rect 152553 61610 152933 61990
rect 152945 61610 153325 61990
rect 153337 61610 153717 61990
rect 153729 61610 154109 61990
rect 154121 61610 154501 61990
rect 152161 61218 152541 61598
rect 152553 61218 152933 61598
rect 152945 61218 153325 61598
rect 153337 61218 153717 61598
rect 153729 61218 154109 61598
rect 154121 61218 154501 61598
rect 152161 60826 152541 61206
rect 152553 60826 152933 61206
rect 152945 60826 153325 61206
rect 153337 60826 153717 61206
rect 153729 60826 154109 61206
rect 154121 60826 154501 61206
rect 152161 60434 152541 60814
rect 152553 60434 152933 60814
rect 152945 60434 153325 60814
rect 153337 60434 153717 60814
rect 153729 60434 154109 60814
rect 154121 60434 154501 60814
rect 152161 60042 152541 60422
rect 152553 60042 152933 60422
rect 152945 60042 153325 60422
rect 153337 60042 153717 60422
rect 153729 60042 154109 60422
rect 154121 60042 154501 60422
rect 82829 59178 83209 59558
rect 83221 59178 83601 59558
rect 83613 59178 83993 59558
rect 84005 59178 84385 59558
rect 84397 59178 84777 59558
rect 84789 59178 85169 59558
rect 82829 58786 83209 59166
rect 83221 58786 83601 59166
rect 83613 58786 83993 59166
rect 84005 58786 84385 59166
rect 84397 58786 84777 59166
rect 84789 58786 85169 59166
rect 82829 58394 83209 58774
rect 83221 58394 83601 58774
rect 83613 58394 83993 58774
rect 84005 58394 84385 58774
rect 84397 58394 84777 58774
rect 84789 58394 85169 58774
rect 82829 58002 83209 58382
rect 83221 58002 83601 58382
rect 83613 58002 83993 58382
rect 84005 58002 84385 58382
rect 84397 58002 84777 58382
rect 84789 58002 85169 58382
rect 82829 57610 83209 57990
rect 83221 57610 83601 57990
rect 83613 57610 83993 57990
rect 84005 57610 84385 57990
rect 84397 57610 84777 57990
rect 84789 57610 85169 57990
rect 82829 57218 83209 57598
rect 83221 57218 83601 57598
rect 83613 57218 83993 57598
rect 84005 57218 84385 57598
rect 84397 57218 84777 57598
rect 84789 57218 85169 57598
rect 82829 56826 83209 57206
rect 83221 56826 83601 57206
rect 83613 56826 83993 57206
rect 84005 56826 84385 57206
rect 84397 56826 84777 57206
rect 84789 56826 85169 57206
rect 82829 56434 83209 56814
rect 83221 56434 83601 56814
rect 83613 56434 83993 56814
rect 84005 56434 84385 56814
rect 84397 56434 84777 56814
rect 84789 56434 85169 56814
rect 82829 56042 83209 56422
rect 83221 56042 83601 56422
rect 83613 56042 83993 56422
rect 84005 56042 84385 56422
rect 84397 56042 84777 56422
rect 84789 56042 85169 56422
rect 98829 59178 99209 59558
rect 99221 59178 99601 59558
rect 99613 59178 99993 59558
rect 100005 59178 100385 59558
rect 100397 59178 100777 59558
rect 100789 59178 101169 59558
rect 98829 58786 99209 59166
rect 99221 58786 99601 59166
rect 99613 58786 99993 59166
rect 100005 58786 100385 59166
rect 100397 58786 100777 59166
rect 100789 58786 101169 59166
rect 98829 58394 99209 58774
rect 99221 58394 99601 58774
rect 99613 58394 99993 58774
rect 100005 58394 100385 58774
rect 100397 58394 100777 58774
rect 100789 58394 101169 58774
rect 98829 58002 99209 58382
rect 99221 58002 99601 58382
rect 99613 58002 99993 58382
rect 100005 58002 100385 58382
rect 100397 58002 100777 58382
rect 100789 58002 101169 58382
rect 98829 57610 99209 57990
rect 99221 57610 99601 57990
rect 99613 57610 99993 57990
rect 100005 57610 100385 57990
rect 100397 57610 100777 57990
rect 100789 57610 101169 57990
rect 98829 57218 99209 57598
rect 99221 57218 99601 57598
rect 99613 57218 99993 57598
rect 100005 57218 100385 57598
rect 100397 57218 100777 57598
rect 100789 57218 101169 57598
rect 98829 56826 99209 57206
rect 99221 56826 99601 57206
rect 99613 56826 99993 57206
rect 100005 56826 100385 57206
rect 100397 56826 100777 57206
rect 100789 56826 101169 57206
rect 98829 56434 99209 56814
rect 99221 56434 99601 56814
rect 99613 56434 99993 56814
rect 100005 56434 100385 56814
rect 100397 56434 100777 56814
rect 100789 56434 101169 56814
rect 98829 56042 99209 56422
rect 99221 56042 99601 56422
rect 99613 56042 99993 56422
rect 100005 56042 100385 56422
rect 100397 56042 100777 56422
rect 100789 56042 101169 56422
rect 114829 59178 115209 59558
rect 115221 59178 115601 59558
rect 115613 59178 115993 59558
rect 116005 59178 116385 59558
rect 116397 59178 116777 59558
rect 116789 59178 117169 59558
rect 114829 58786 115209 59166
rect 115221 58786 115601 59166
rect 115613 58786 115993 59166
rect 116005 58786 116385 59166
rect 116397 58786 116777 59166
rect 116789 58786 117169 59166
rect 114829 58394 115209 58774
rect 115221 58394 115601 58774
rect 115613 58394 115993 58774
rect 116005 58394 116385 58774
rect 116397 58394 116777 58774
rect 116789 58394 117169 58774
rect 114829 58002 115209 58382
rect 115221 58002 115601 58382
rect 115613 58002 115993 58382
rect 116005 58002 116385 58382
rect 116397 58002 116777 58382
rect 116789 58002 117169 58382
rect 114829 57610 115209 57990
rect 115221 57610 115601 57990
rect 115613 57610 115993 57990
rect 116005 57610 116385 57990
rect 116397 57610 116777 57990
rect 116789 57610 117169 57990
rect 114829 57218 115209 57598
rect 115221 57218 115601 57598
rect 115613 57218 115993 57598
rect 116005 57218 116385 57598
rect 116397 57218 116777 57598
rect 116789 57218 117169 57598
rect 114829 56826 115209 57206
rect 115221 56826 115601 57206
rect 115613 56826 115993 57206
rect 116005 56826 116385 57206
rect 116397 56826 116777 57206
rect 116789 56826 117169 57206
rect 114829 56434 115209 56814
rect 115221 56434 115601 56814
rect 115613 56434 115993 56814
rect 116005 56434 116385 56814
rect 116397 56434 116777 56814
rect 116789 56434 117169 56814
rect 114829 56042 115209 56422
rect 115221 56042 115601 56422
rect 115613 56042 115993 56422
rect 116005 56042 116385 56422
rect 116397 56042 116777 56422
rect 116789 56042 117169 56422
rect 146829 59178 147209 59558
rect 147221 59178 147601 59558
rect 147613 59178 147993 59558
rect 148005 59178 148385 59558
rect 148397 59178 148777 59558
rect 148789 59178 149169 59558
rect 146829 58786 147209 59166
rect 147221 58786 147601 59166
rect 147613 58786 147993 59166
rect 148005 58786 148385 59166
rect 148397 58786 148777 59166
rect 148789 58786 149169 59166
rect 146829 58394 147209 58774
rect 147221 58394 147601 58774
rect 147613 58394 147993 58774
rect 148005 58394 148385 58774
rect 148397 58394 148777 58774
rect 148789 58394 149169 58774
rect 146829 58002 147209 58382
rect 147221 58002 147601 58382
rect 147613 58002 147993 58382
rect 148005 58002 148385 58382
rect 148397 58002 148777 58382
rect 148789 58002 149169 58382
rect 146829 57610 147209 57990
rect 147221 57610 147601 57990
rect 147613 57610 147993 57990
rect 148005 57610 148385 57990
rect 148397 57610 148777 57990
rect 148789 57610 149169 57990
rect 146829 57218 147209 57598
rect 147221 57218 147601 57598
rect 147613 57218 147993 57598
rect 148005 57218 148385 57598
rect 148397 57218 148777 57598
rect 148789 57218 149169 57598
rect 146829 56826 147209 57206
rect 147221 56826 147601 57206
rect 147613 56826 147993 57206
rect 148005 56826 148385 57206
rect 148397 56826 148777 57206
rect 148789 56826 149169 57206
rect 146829 56434 147209 56814
rect 147221 56434 147601 56814
rect 147613 56434 147993 56814
rect 148005 56434 148385 56814
rect 148397 56434 148777 56814
rect 148789 56434 149169 56814
rect 146829 56042 147209 56422
rect 147221 56042 147601 56422
rect 147613 56042 147993 56422
rect 148005 56042 148385 56422
rect 148397 56042 148777 56422
rect 148789 56042 149169 56422
<< metal7 >>
rect 65000 196000 79000 210000
rect 81000 196000 95000 210000
rect 97000 196000 111000 210000
rect 113000 196000 127000 210000
rect 129000 196000 143000 210000
rect 145000 196000 159000 210000
rect 82666 167958 85332 168000
rect 82666 167578 82829 167958
rect 83209 167578 83221 167958
rect 83601 167578 83613 167958
rect 83993 167578 84005 167958
rect 84385 167578 84397 167958
rect 84777 167578 84789 167958
rect 85169 167578 85332 167958
rect 82666 167566 85332 167578
rect 82666 167186 82829 167566
rect 83209 167186 83221 167566
rect 83601 167186 83613 167566
rect 83993 167186 84005 167566
rect 84385 167186 84397 167566
rect 84777 167186 84789 167566
rect 85169 167186 85332 167566
rect 82666 167174 85332 167186
rect 82666 166794 82829 167174
rect 83209 166794 83221 167174
rect 83601 166794 83613 167174
rect 83993 166794 84005 167174
rect 84385 166794 84397 167174
rect 84777 166794 84789 167174
rect 85169 166794 85332 167174
rect 82666 166782 85332 166794
rect 82666 166402 82829 166782
rect 83209 166402 83221 166782
rect 83601 166402 83613 166782
rect 83993 166402 84005 166782
rect 84385 166402 84397 166782
rect 84777 166402 84789 166782
rect 85169 166402 85332 166782
rect 82666 166390 85332 166402
rect 82666 166010 82829 166390
rect 83209 166010 83221 166390
rect 83601 166010 83613 166390
rect 83993 166010 84005 166390
rect 84385 166010 84397 166390
rect 84777 166010 84789 166390
rect 85169 166010 85332 166390
rect 82666 165998 85332 166010
rect 82666 165618 82829 165998
rect 83209 165618 83221 165998
rect 83601 165618 83613 165998
rect 83993 165618 84005 165998
rect 84385 165618 84397 165998
rect 84777 165618 84789 165998
rect 85169 165618 85332 165998
rect 82666 165606 85332 165618
rect 82666 165226 82829 165606
rect 83209 165226 83221 165606
rect 83601 165226 83613 165606
rect 83993 165226 84005 165606
rect 84385 165226 84397 165606
rect 84777 165226 84789 165606
rect 85169 165226 85332 165606
rect 82666 165214 85332 165226
rect 82666 164834 82829 165214
rect 83209 164834 83221 165214
rect 83601 164834 83613 165214
rect 83993 164834 84005 165214
rect 84385 164834 84397 165214
rect 84777 164834 84789 165214
rect 85169 164834 85332 165214
rect 82666 164822 85332 164834
rect 82666 164442 82829 164822
rect 83209 164442 83221 164822
rect 83601 164442 83613 164822
rect 83993 164442 84005 164822
rect 84385 164442 84397 164822
rect 84777 164442 84789 164822
rect 85169 164442 85332 164822
rect 71998 163958 74664 164000
rect 71998 163578 72161 163958
rect 72541 163578 72553 163958
rect 72933 163578 72945 163958
rect 73325 163578 73337 163958
rect 73717 163578 73729 163958
rect 74109 163578 74121 163958
rect 74501 163578 74664 163958
rect 71998 163566 74664 163578
rect 71998 163186 72161 163566
rect 72541 163186 72553 163566
rect 72933 163186 72945 163566
rect 73325 163186 73337 163566
rect 73717 163186 73729 163566
rect 74109 163186 74121 163566
rect 74501 163186 74664 163566
rect 71998 163174 74664 163186
rect 71998 162794 72161 163174
rect 72541 162794 72553 163174
rect 72933 162794 72945 163174
rect 73325 162794 73337 163174
rect 73717 162794 73729 163174
rect 74109 162794 74121 163174
rect 74501 162794 74664 163174
rect 71998 162782 74664 162794
rect 71998 162402 72161 162782
rect 72541 162402 72553 162782
rect 72933 162402 72945 162782
rect 73325 162402 73337 162782
rect 73717 162402 73729 162782
rect 74109 162402 74121 162782
rect 74501 162402 74664 162782
rect 71998 162390 74664 162402
rect 71998 162010 72161 162390
rect 72541 162010 72553 162390
rect 72933 162010 72945 162390
rect 73325 162010 73337 162390
rect 73717 162010 73729 162390
rect 74109 162010 74121 162390
rect 74501 162010 74664 162390
rect 71998 161998 74664 162010
rect 71998 161618 72161 161998
rect 72541 161618 72553 161998
rect 72933 161618 72945 161998
rect 73325 161618 73337 161998
rect 73717 161618 73729 161998
rect 74109 161618 74121 161998
rect 74501 161618 74664 161998
rect 71998 161606 74664 161618
rect 71998 161226 72161 161606
rect 72541 161226 72553 161606
rect 72933 161226 72945 161606
rect 73325 161226 73337 161606
rect 73717 161226 73729 161606
rect 74109 161226 74121 161606
rect 74501 161226 74664 161606
rect 71998 161214 74664 161226
rect 71998 160834 72161 161214
rect 72541 160834 72553 161214
rect 72933 160834 72945 161214
rect 73325 160834 73337 161214
rect 73717 160834 73729 161214
rect 74109 160834 74121 161214
rect 74501 160834 74664 161214
rect 71998 160822 74664 160834
rect 71998 160442 72161 160822
rect 72541 160442 72553 160822
rect 72933 160442 72945 160822
rect 73325 160442 73337 160822
rect 73717 160442 73729 160822
rect 74109 160442 74121 160822
rect 74501 160442 74664 160822
rect 14000 145000 28000 159000
rect 71998 155656 74664 160442
rect 82666 155656 85332 164442
rect 98666 167958 101332 168000
rect 98666 167578 98829 167958
rect 99209 167578 99221 167958
rect 99601 167578 99613 167958
rect 99993 167578 100005 167958
rect 100385 167578 100397 167958
rect 100777 167578 100789 167958
rect 101169 167578 101332 167958
rect 98666 167566 101332 167578
rect 98666 167186 98829 167566
rect 99209 167186 99221 167566
rect 99601 167186 99613 167566
rect 99993 167186 100005 167566
rect 100385 167186 100397 167566
rect 100777 167186 100789 167566
rect 101169 167186 101332 167566
rect 98666 167174 101332 167186
rect 98666 166794 98829 167174
rect 99209 166794 99221 167174
rect 99601 166794 99613 167174
rect 99993 166794 100005 167174
rect 100385 166794 100397 167174
rect 100777 166794 100789 167174
rect 101169 166794 101332 167174
rect 98666 166782 101332 166794
rect 98666 166402 98829 166782
rect 99209 166402 99221 166782
rect 99601 166402 99613 166782
rect 99993 166402 100005 166782
rect 100385 166402 100397 166782
rect 100777 166402 100789 166782
rect 101169 166402 101332 166782
rect 98666 166390 101332 166402
rect 98666 166010 98829 166390
rect 99209 166010 99221 166390
rect 99601 166010 99613 166390
rect 99993 166010 100005 166390
rect 100385 166010 100397 166390
rect 100777 166010 100789 166390
rect 101169 166010 101332 166390
rect 98666 165998 101332 166010
rect 98666 165618 98829 165998
rect 99209 165618 99221 165998
rect 99601 165618 99613 165998
rect 99993 165618 100005 165998
rect 100385 165618 100397 165998
rect 100777 165618 100789 165998
rect 101169 165618 101332 165998
rect 98666 165606 101332 165618
rect 98666 165226 98829 165606
rect 99209 165226 99221 165606
rect 99601 165226 99613 165606
rect 99993 165226 100005 165606
rect 100385 165226 100397 165606
rect 100777 165226 100789 165606
rect 101169 165226 101332 165606
rect 98666 165214 101332 165226
rect 98666 164834 98829 165214
rect 99209 164834 99221 165214
rect 99601 164834 99613 165214
rect 99993 164834 100005 165214
rect 100385 164834 100397 165214
rect 100777 164834 100789 165214
rect 101169 164834 101332 165214
rect 98666 164822 101332 164834
rect 98666 164442 98829 164822
rect 99209 164442 99221 164822
rect 99601 164442 99613 164822
rect 99993 164442 100005 164822
rect 100385 164442 100397 164822
rect 100777 164442 100789 164822
rect 101169 164442 101332 164822
rect 87998 163958 90664 164000
rect 87998 163578 88161 163958
rect 88541 163578 88553 163958
rect 88933 163578 88945 163958
rect 89325 163578 89337 163958
rect 89717 163578 89729 163958
rect 90109 163578 90121 163958
rect 90501 163578 90664 163958
rect 87998 163566 90664 163578
rect 87998 163186 88161 163566
rect 88541 163186 88553 163566
rect 88933 163186 88945 163566
rect 89325 163186 89337 163566
rect 89717 163186 89729 163566
rect 90109 163186 90121 163566
rect 90501 163186 90664 163566
rect 87998 163174 90664 163186
rect 87998 162794 88161 163174
rect 88541 162794 88553 163174
rect 88933 162794 88945 163174
rect 89325 162794 89337 163174
rect 89717 162794 89729 163174
rect 90109 162794 90121 163174
rect 90501 162794 90664 163174
rect 87998 162782 90664 162794
rect 87998 162402 88161 162782
rect 88541 162402 88553 162782
rect 88933 162402 88945 162782
rect 89325 162402 89337 162782
rect 89717 162402 89729 162782
rect 90109 162402 90121 162782
rect 90501 162402 90664 162782
rect 87998 162390 90664 162402
rect 87998 162010 88161 162390
rect 88541 162010 88553 162390
rect 88933 162010 88945 162390
rect 89325 162010 89337 162390
rect 89717 162010 89729 162390
rect 90109 162010 90121 162390
rect 90501 162010 90664 162390
rect 87998 161998 90664 162010
rect 87998 161618 88161 161998
rect 88541 161618 88553 161998
rect 88933 161618 88945 161998
rect 89325 161618 89337 161998
rect 89717 161618 89729 161998
rect 90109 161618 90121 161998
rect 90501 161618 90664 161998
rect 87998 161606 90664 161618
rect 87998 161226 88161 161606
rect 88541 161226 88553 161606
rect 88933 161226 88945 161606
rect 89325 161226 89337 161606
rect 89717 161226 89729 161606
rect 90109 161226 90121 161606
rect 90501 161226 90664 161606
rect 87998 161214 90664 161226
rect 87998 160834 88161 161214
rect 88541 160834 88553 161214
rect 88933 160834 88945 161214
rect 89325 160834 89337 161214
rect 89717 160834 89729 161214
rect 90109 160834 90121 161214
rect 90501 160834 90664 161214
rect 87998 160822 90664 160834
rect 87998 160442 88161 160822
rect 88541 160442 88553 160822
rect 88933 160442 88945 160822
rect 89325 160442 89337 160822
rect 89717 160442 89729 160822
rect 90109 160442 90121 160822
rect 90501 160442 90664 160822
rect 87998 155656 90664 160442
rect 98666 155656 101332 164442
rect 114666 167958 117332 168000
rect 114666 167578 114829 167958
rect 115209 167578 115221 167958
rect 115601 167578 115613 167958
rect 115993 167578 116005 167958
rect 116385 167578 116397 167958
rect 116777 167578 116789 167958
rect 117169 167578 117332 167958
rect 114666 167566 117332 167578
rect 114666 167186 114829 167566
rect 115209 167186 115221 167566
rect 115601 167186 115613 167566
rect 115993 167186 116005 167566
rect 116385 167186 116397 167566
rect 116777 167186 116789 167566
rect 117169 167186 117332 167566
rect 114666 167174 117332 167186
rect 114666 166794 114829 167174
rect 115209 166794 115221 167174
rect 115601 166794 115613 167174
rect 115993 166794 116005 167174
rect 116385 166794 116397 167174
rect 116777 166794 116789 167174
rect 117169 166794 117332 167174
rect 114666 166782 117332 166794
rect 114666 166402 114829 166782
rect 115209 166402 115221 166782
rect 115601 166402 115613 166782
rect 115993 166402 116005 166782
rect 116385 166402 116397 166782
rect 116777 166402 116789 166782
rect 117169 166402 117332 166782
rect 114666 166390 117332 166402
rect 114666 166010 114829 166390
rect 115209 166010 115221 166390
rect 115601 166010 115613 166390
rect 115993 166010 116005 166390
rect 116385 166010 116397 166390
rect 116777 166010 116789 166390
rect 117169 166010 117332 166390
rect 114666 165998 117332 166010
rect 114666 165618 114829 165998
rect 115209 165618 115221 165998
rect 115601 165618 115613 165998
rect 115993 165618 116005 165998
rect 116385 165618 116397 165998
rect 116777 165618 116789 165998
rect 117169 165618 117332 165998
rect 114666 165606 117332 165618
rect 114666 165226 114829 165606
rect 115209 165226 115221 165606
rect 115601 165226 115613 165606
rect 115993 165226 116005 165606
rect 116385 165226 116397 165606
rect 116777 165226 116789 165606
rect 117169 165226 117332 165606
rect 114666 165214 117332 165226
rect 114666 164834 114829 165214
rect 115209 164834 115221 165214
rect 115601 164834 115613 165214
rect 115993 164834 116005 165214
rect 116385 164834 116397 165214
rect 116777 164834 116789 165214
rect 117169 164834 117332 165214
rect 114666 164822 117332 164834
rect 114666 164442 114829 164822
rect 115209 164442 115221 164822
rect 115601 164442 115613 164822
rect 115993 164442 116005 164822
rect 116385 164442 116397 164822
rect 116777 164442 116789 164822
rect 117169 164442 117332 164822
rect 103998 163958 106664 164000
rect 103998 163578 104161 163958
rect 104541 163578 104553 163958
rect 104933 163578 104945 163958
rect 105325 163578 105337 163958
rect 105717 163578 105729 163958
rect 106109 163578 106121 163958
rect 106501 163578 106664 163958
rect 103998 163566 106664 163578
rect 103998 163186 104161 163566
rect 104541 163186 104553 163566
rect 104933 163186 104945 163566
rect 105325 163186 105337 163566
rect 105717 163186 105729 163566
rect 106109 163186 106121 163566
rect 106501 163186 106664 163566
rect 103998 163174 106664 163186
rect 103998 162794 104161 163174
rect 104541 162794 104553 163174
rect 104933 162794 104945 163174
rect 105325 162794 105337 163174
rect 105717 162794 105729 163174
rect 106109 162794 106121 163174
rect 106501 162794 106664 163174
rect 103998 162782 106664 162794
rect 103998 162402 104161 162782
rect 104541 162402 104553 162782
rect 104933 162402 104945 162782
rect 105325 162402 105337 162782
rect 105717 162402 105729 162782
rect 106109 162402 106121 162782
rect 106501 162402 106664 162782
rect 103998 162390 106664 162402
rect 103998 162010 104161 162390
rect 104541 162010 104553 162390
rect 104933 162010 104945 162390
rect 105325 162010 105337 162390
rect 105717 162010 105729 162390
rect 106109 162010 106121 162390
rect 106501 162010 106664 162390
rect 103998 161998 106664 162010
rect 103998 161618 104161 161998
rect 104541 161618 104553 161998
rect 104933 161618 104945 161998
rect 105325 161618 105337 161998
rect 105717 161618 105729 161998
rect 106109 161618 106121 161998
rect 106501 161618 106664 161998
rect 103998 161606 106664 161618
rect 103998 161226 104161 161606
rect 104541 161226 104553 161606
rect 104933 161226 104945 161606
rect 105325 161226 105337 161606
rect 105717 161226 105729 161606
rect 106109 161226 106121 161606
rect 106501 161226 106664 161606
rect 103998 161214 106664 161226
rect 103998 160834 104161 161214
rect 104541 160834 104553 161214
rect 104933 160834 104945 161214
rect 105325 160834 105337 161214
rect 105717 160834 105729 161214
rect 106109 160834 106121 161214
rect 106501 160834 106664 161214
rect 103998 160822 106664 160834
rect 103998 160442 104161 160822
rect 104541 160442 104553 160822
rect 104933 160442 104945 160822
rect 105325 160442 105337 160822
rect 105717 160442 105729 160822
rect 106109 160442 106121 160822
rect 106501 160442 106664 160822
rect 103998 155656 106664 160442
rect 114666 155656 117332 164442
rect 130666 167958 133332 168000
rect 130666 167578 130829 167958
rect 131209 167578 131221 167958
rect 131601 167578 131613 167958
rect 131993 167578 132005 167958
rect 132385 167578 132397 167958
rect 132777 167578 132789 167958
rect 133169 167578 133332 167958
rect 130666 167566 133332 167578
rect 130666 167186 130829 167566
rect 131209 167186 131221 167566
rect 131601 167186 131613 167566
rect 131993 167186 132005 167566
rect 132385 167186 132397 167566
rect 132777 167186 132789 167566
rect 133169 167186 133332 167566
rect 130666 167174 133332 167186
rect 130666 166794 130829 167174
rect 131209 166794 131221 167174
rect 131601 166794 131613 167174
rect 131993 166794 132005 167174
rect 132385 166794 132397 167174
rect 132777 166794 132789 167174
rect 133169 166794 133332 167174
rect 130666 166782 133332 166794
rect 130666 166402 130829 166782
rect 131209 166402 131221 166782
rect 131601 166402 131613 166782
rect 131993 166402 132005 166782
rect 132385 166402 132397 166782
rect 132777 166402 132789 166782
rect 133169 166402 133332 166782
rect 130666 166390 133332 166402
rect 130666 166010 130829 166390
rect 131209 166010 131221 166390
rect 131601 166010 131613 166390
rect 131993 166010 132005 166390
rect 132385 166010 132397 166390
rect 132777 166010 132789 166390
rect 133169 166010 133332 166390
rect 130666 165998 133332 166010
rect 130666 165618 130829 165998
rect 131209 165618 131221 165998
rect 131601 165618 131613 165998
rect 131993 165618 132005 165998
rect 132385 165618 132397 165998
rect 132777 165618 132789 165998
rect 133169 165618 133332 165998
rect 130666 165606 133332 165618
rect 130666 165226 130829 165606
rect 131209 165226 131221 165606
rect 131601 165226 131613 165606
rect 131993 165226 132005 165606
rect 132385 165226 132397 165606
rect 132777 165226 132789 165606
rect 133169 165226 133332 165606
rect 130666 165214 133332 165226
rect 130666 164834 130829 165214
rect 131209 164834 131221 165214
rect 131601 164834 131613 165214
rect 131993 164834 132005 165214
rect 132385 164834 132397 165214
rect 132777 164834 132789 165214
rect 133169 164834 133332 165214
rect 130666 164822 133332 164834
rect 130666 164442 130829 164822
rect 131209 164442 131221 164822
rect 131601 164442 131613 164822
rect 131993 164442 132005 164822
rect 132385 164442 132397 164822
rect 132777 164442 132789 164822
rect 133169 164442 133332 164822
rect 119998 163958 122664 164000
rect 119998 163578 120161 163958
rect 120541 163578 120553 163958
rect 120933 163578 120945 163958
rect 121325 163578 121337 163958
rect 121717 163578 121729 163958
rect 122109 163578 122121 163958
rect 122501 163578 122664 163958
rect 119998 163566 122664 163578
rect 119998 163186 120161 163566
rect 120541 163186 120553 163566
rect 120933 163186 120945 163566
rect 121325 163186 121337 163566
rect 121717 163186 121729 163566
rect 122109 163186 122121 163566
rect 122501 163186 122664 163566
rect 119998 163174 122664 163186
rect 119998 162794 120161 163174
rect 120541 162794 120553 163174
rect 120933 162794 120945 163174
rect 121325 162794 121337 163174
rect 121717 162794 121729 163174
rect 122109 162794 122121 163174
rect 122501 162794 122664 163174
rect 119998 162782 122664 162794
rect 119998 162402 120161 162782
rect 120541 162402 120553 162782
rect 120933 162402 120945 162782
rect 121325 162402 121337 162782
rect 121717 162402 121729 162782
rect 122109 162402 122121 162782
rect 122501 162402 122664 162782
rect 119998 162390 122664 162402
rect 119998 162010 120161 162390
rect 120541 162010 120553 162390
rect 120933 162010 120945 162390
rect 121325 162010 121337 162390
rect 121717 162010 121729 162390
rect 122109 162010 122121 162390
rect 122501 162010 122664 162390
rect 119998 161998 122664 162010
rect 119998 161618 120161 161998
rect 120541 161618 120553 161998
rect 120933 161618 120945 161998
rect 121325 161618 121337 161998
rect 121717 161618 121729 161998
rect 122109 161618 122121 161998
rect 122501 161618 122664 161998
rect 119998 161606 122664 161618
rect 119998 161226 120161 161606
rect 120541 161226 120553 161606
rect 120933 161226 120945 161606
rect 121325 161226 121337 161606
rect 121717 161226 121729 161606
rect 122109 161226 122121 161606
rect 122501 161226 122664 161606
rect 119998 161214 122664 161226
rect 119998 160834 120161 161214
rect 120541 160834 120553 161214
rect 120933 160834 120945 161214
rect 121325 160834 121337 161214
rect 121717 160834 121729 161214
rect 122109 160834 122121 161214
rect 122501 160834 122664 161214
rect 119998 160822 122664 160834
rect 119998 160442 120161 160822
rect 120541 160442 120553 160822
rect 120933 160442 120945 160822
rect 121325 160442 121337 160822
rect 121717 160442 121729 160822
rect 122109 160442 122121 160822
rect 122501 160442 122664 160822
rect 119998 155656 122664 160442
rect 130666 155656 133332 164442
rect 146666 167958 149332 168000
rect 146666 167578 146829 167958
rect 147209 167578 147221 167958
rect 147601 167578 147613 167958
rect 147993 167578 148005 167958
rect 148385 167578 148397 167958
rect 148777 167578 148789 167958
rect 149169 167578 149332 167958
rect 146666 167566 149332 167578
rect 146666 167186 146829 167566
rect 147209 167186 147221 167566
rect 147601 167186 147613 167566
rect 147993 167186 148005 167566
rect 148385 167186 148397 167566
rect 148777 167186 148789 167566
rect 149169 167186 149332 167566
rect 146666 167174 149332 167186
rect 146666 166794 146829 167174
rect 147209 166794 147221 167174
rect 147601 166794 147613 167174
rect 147993 166794 148005 167174
rect 148385 166794 148397 167174
rect 148777 166794 148789 167174
rect 149169 166794 149332 167174
rect 146666 166782 149332 166794
rect 146666 166402 146829 166782
rect 147209 166402 147221 166782
rect 147601 166402 147613 166782
rect 147993 166402 148005 166782
rect 148385 166402 148397 166782
rect 148777 166402 148789 166782
rect 149169 166402 149332 166782
rect 146666 166390 149332 166402
rect 146666 166010 146829 166390
rect 147209 166010 147221 166390
rect 147601 166010 147613 166390
rect 147993 166010 148005 166390
rect 148385 166010 148397 166390
rect 148777 166010 148789 166390
rect 149169 166010 149332 166390
rect 146666 165998 149332 166010
rect 146666 165618 146829 165998
rect 147209 165618 147221 165998
rect 147601 165618 147613 165998
rect 147993 165618 148005 165998
rect 148385 165618 148397 165998
rect 148777 165618 148789 165998
rect 149169 165618 149332 165998
rect 146666 165606 149332 165618
rect 146666 165226 146829 165606
rect 147209 165226 147221 165606
rect 147601 165226 147613 165606
rect 147993 165226 148005 165606
rect 148385 165226 148397 165606
rect 148777 165226 148789 165606
rect 149169 165226 149332 165606
rect 146666 165214 149332 165226
rect 146666 164834 146829 165214
rect 147209 164834 147221 165214
rect 147601 164834 147613 165214
rect 147993 164834 148005 165214
rect 148385 164834 148397 165214
rect 148777 164834 148789 165214
rect 149169 164834 149332 165214
rect 146666 164822 149332 164834
rect 146666 164442 146829 164822
rect 147209 164442 147221 164822
rect 147601 164442 147613 164822
rect 147993 164442 148005 164822
rect 148385 164442 148397 164822
rect 148777 164442 148789 164822
rect 149169 164442 149332 164822
rect 135998 163958 138664 164000
rect 135998 163578 136161 163958
rect 136541 163578 136553 163958
rect 136933 163578 136945 163958
rect 137325 163578 137337 163958
rect 137717 163578 137729 163958
rect 138109 163578 138121 163958
rect 138501 163578 138664 163958
rect 135998 163566 138664 163578
rect 135998 163186 136161 163566
rect 136541 163186 136553 163566
rect 136933 163186 136945 163566
rect 137325 163186 137337 163566
rect 137717 163186 137729 163566
rect 138109 163186 138121 163566
rect 138501 163186 138664 163566
rect 135998 163174 138664 163186
rect 135998 162794 136161 163174
rect 136541 162794 136553 163174
rect 136933 162794 136945 163174
rect 137325 162794 137337 163174
rect 137717 162794 137729 163174
rect 138109 162794 138121 163174
rect 138501 162794 138664 163174
rect 135998 162782 138664 162794
rect 135998 162402 136161 162782
rect 136541 162402 136553 162782
rect 136933 162402 136945 162782
rect 137325 162402 137337 162782
rect 137717 162402 137729 162782
rect 138109 162402 138121 162782
rect 138501 162402 138664 162782
rect 135998 162390 138664 162402
rect 135998 162010 136161 162390
rect 136541 162010 136553 162390
rect 136933 162010 136945 162390
rect 137325 162010 137337 162390
rect 137717 162010 137729 162390
rect 138109 162010 138121 162390
rect 138501 162010 138664 162390
rect 135998 161998 138664 162010
rect 135998 161618 136161 161998
rect 136541 161618 136553 161998
rect 136933 161618 136945 161998
rect 137325 161618 137337 161998
rect 137717 161618 137729 161998
rect 138109 161618 138121 161998
rect 138501 161618 138664 161998
rect 135998 161606 138664 161618
rect 135998 161226 136161 161606
rect 136541 161226 136553 161606
rect 136933 161226 136945 161606
rect 137325 161226 137337 161606
rect 137717 161226 137729 161606
rect 138109 161226 138121 161606
rect 138501 161226 138664 161606
rect 135998 161214 138664 161226
rect 135998 160834 136161 161214
rect 136541 160834 136553 161214
rect 136933 160834 136945 161214
rect 137325 160834 137337 161214
rect 137717 160834 137729 161214
rect 138109 160834 138121 161214
rect 138501 160834 138664 161214
rect 135998 160822 138664 160834
rect 135998 160442 136161 160822
rect 136541 160442 136553 160822
rect 136933 160442 136945 160822
rect 137325 160442 137337 160822
rect 137717 160442 137729 160822
rect 138109 160442 138121 160822
rect 138501 160442 138664 160822
rect 135998 155656 138664 160442
rect 146666 155656 149332 164442
rect 151998 163958 154664 164000
rect 151998 163578 152161 163958
rect 152541 163578 152553 163958
rect 152933 163578 152945 163958
rect 153325 163578 153337 163958
rect 153717 163578 153729 163958
rect 154109 163578 154121 163958
rect 154501 163578 154664 163958
rect 151998 163566 154664 163578
rect 151998 163186 152161 163566
rect 152541 163186 152553 163566
rect 152933 163186 152945 163566
rect 153325 163186 153337 163566
rect 153717 163186 153729 163566
rect 154109 163186 154121 163566
rect 154501 163186 154664 163566
rect 151998 163174 154664 163186
rect 151998 162794 152161 163174
rect 152541 162794 152553 163174
rect 152933 162794 152945 163174
rect 153325 162794 153337 163174
rect 153717 162794 153729 163174
rect 154109 162794 154121 163174
rect 154501 162794 154664 163174
rect 151998 162782 154664 162794
rect 151998 162402 152161 162782
rect 152541 162402 152553 162782
rect 152933 162402 152945 162782
rect 153325 162402 153337 162782
rect 153717 162402 153729 162782
rect 154109 162402 154121 162782
rect 154501 162402 154664 162782
rect 151998 162390 154664 162402
rect 151998 162010 152161 162390
rect 152541 162010 152553 162390
rect 152933 162010 152945 162390
rect 153325 162010 153337 162390
rect 153717 162010 153729 162390
rect 154109 162010 154121 162390
rect 154501 162010 154664 162390
rect 151998 161998 154664 162010
rect 151998 161618 152161 161998
rect 152541 161618 152553 161998
rect 152933 161618 152945 161998
rect 153325 161618 153337 161998
rect 153717 161618 153729 161998
rect 154109 161618 154121 161998
rect 154501 161618 154664 161998
rect 151998 161606 154664 161618
rect 151998 161226 152161 161606
rect 152541 161226 152553 161606
rect 152933 161226 152945 161606
rect 153325 161226 153337 161606
rect 153717 161226 153729 161606
rect 154109 161226 154121 161606
rect 154501 161226 154664 161606
rect 151998 161214 154664 161226
rect 151998 160834 152161 161214
rect 152541 160834 152553 161214
rect 152933 160834 152945 161214
rect 153325 160834 153337 161214
rect 153717 160834 153729 161214
rect 154109 160834 154121 161214
rect 154501 160834 154664 161214
rect 151998 160822 154664 160834
rect 151998 160442 152161 160822
rect 152541 160442 152553 160822
rect 152933 160442 152945 160822
rect 153325 160442 153337 160822
rect 153717 160442 153729 160822
rect 154109 160442 154121 160822
rect 154501 160442 154664 160822
rect 151998 155656 154664 160442
rect 68316 155142 155652 155256
rect 68316 154762 68430 155142
rect 68810 154762 68822 155142
rect 69202 154762 75386 155142
rect 75766 154762 90506 155142
rect 90886 154762 105626 155142
rect 106006 154762 120746 155142
rect 121126 154762 135866 155142
rect 136246 154762 150986 155142
rect 151366 154762 154766 155142
rect 155146 154762 155158 155142
rect 155538 154762 155652 155142
rect 68316 154750 155652 154762
rect 60000 154501 67916 154664
rect 60000 154121 60042 154501
rect 60422 154121 60434 154501
rect 60814 154121 60826 154501
rect 61206 154121 61218 154501
rect 61598 154121 61610 154501
rect 61990 154121 62002 154501
rect 62382 154121 62394 154501
rect 62774 154121 62786 154501
rect 63166 154121 63178 154501
rect 63558 154121 67916 154501
rect 68316 154370 68430 154750
rect 68810 154370 68822 154750
rect 69202 154370 75386 154750
rect 75766 154370 90506 154750
rect 90886 154370 105626 154750
rect 106006 154370 120746 154750
rect 121126 154370 135866 154750
rect 136246 154370 150986 154750
rect 151366 154370 154766 154750
rect 155146 154370 155158 154750
rect 155538 154370 155652 154750
rect 68316 154256 155652 154370
rect 156052 154501 164000 154664
rect 60000 154109 67916 154121
rect 60000 153729 60042 154109
rect 60422 153729 60434 154109
rect 60814 153729 60826 154109
rect 61206 153729 61218 154109
rect 61598 153729 61610 154109
rect 61990 153729 62002 154109
rect 62382 153729 62394 154109
rect 62774 153729 62786 154109
rect 63166 153729 63178 154109
rect 63558 153729 67916 154109
rect 156052 154121 160442 154501
rect 160822 154121 160834 154501
rect 161214 154121 161226 154501
rect 161606 154121 161618 154501
rect 161998 154121 162010 154501
rect 162390 154121 162402 154501
rect 162782 154121 162794 154501
rect 163174 154121 163186 154501
rect 163566 154121 163578 154501
rect 163958 154121 164000 154501
rect 156052 154109 164000 154121
rect 60000 153717 67916 153729
rect 60000 153337 60042 153717
rect 60422 153337 60434 153717
rect 60814 153337 60826 153717
rect 61206 153337 61218 153717
rect 61598 153337 61610 153717
rect 61990 153337 62002 153717
rect 62382 153337 62394 153717
rect 62774 153337 62786 153717
rect 63166 153337 63178 153717
rect 63558 153337 67916 153717
rect 60000 153325 67916 153337
rect 60000 152945 60042 153325
rect 60422 152945 60434 153325
rect 60814 152945 60826 153325
rect 61206 152945 61218 153325
rect 61598 152945 61610 153325
rect 61990 152945 62002 153325
rect 62382 152945 62394 153325
rect 62774 152945 62786 153325
rect 63166 152945 63178 153325
rect 63558 152945 67916 153325
rect 60000 152933 67916 152945
rect 60000 152553 60042 152933
rect 60422 152553 60434 152933
rect 60814 152553 60826 152933
rect 61206 152553 61218 152933
rect 61598 152553 61610 152933
rect 61990 152553 62002 152933
rect 62382 152553 62394 152933
rect 62774 152553 62786 152933
rect 63166 152553 63178 152933
rect 63558 152553 67916 152933
rect 69716 153742 154252 153856
rect 69716 153362 69830 153742
rect 70210 153362 70222 153742
rect 70602 153362 74146 153742
rect 74526 153362 89266 153742
rect 89646 153362 104386 153742
rect 104766 153362 119506 153742
rect 119886 153362 134626 153742
rect 135006 153362 149746 153742
rect 150126 153362 153366 153742
rect 153746 153362 153758 153742
rect 154138 153362 154252 153742
rect 69716 153350 154252 153362
rect 69716 152970 69830 153350
rect 70210 152970 70222 153350
rect 70602 152970 74146 153350
rect 74526 152970 89266 153350
rect 89646 152970 104386 153350
rect 104766 152970 119506 153350
rect 119886 152970 134626 153350
rect 135006 152970 149746 153350
rect 150126 152970 153366 153350
rect 153746 152970 153758 153350
rect 154138 152970 154252 153350
rect 69716 152856 154252 152970
rect 156052 153729 160442 154109
rect 160822 153729 160834 154109
rect 161214 153729 161226 154109
rect 161606 153729 161618 154109
rect 161998 153729 162010 154109
rect 162390 153729 162402 154109
rect 162782 153729 162794 154109
rect 163174 153729 163186 154109
rect 163566 153729 163578 154109
rect 163958 153729 164000 154109
rect 156052 153717 164000 153729
rect 156052 153337 160442 153717
rect 160822 153337 160834 153717
rect 161214 153337 161226 153717
rect 161606 153337 161618 153717
rect 161998 153337 162010 153717
rect 162390 153337 162402 153717
rect 162782 153337 162794 153717
rect 163174 153337 163186 153717
rect 163566 153337 163578 153717
rect 163958 153337 164000 153717
rect 156052 153325 164000 153337
rect 156052 152945 160442 153325
rect 160822 152945 160834 153325
rect 161214 152945 161226 153325
rect 161606 152945 161618 153325
rect 161998 152945 162010 153325
rect 162390 152945 162402 153325
rect 162782 152945 162794 153325
rect 163174 152945 163186 153325
rect 163566 152945 163578 153325
rect 163958 152945 164000 153325
rect 156052 152933 164000 152945
rect 60000 152541 67916 152553
rect 60000 152161 60042 152541
rect 60422 152161 60434 152541
rect 60814 152161 60826 152541
rect 61206 152161 61218 152541
rect 61598 152161 61610 152541
rect 61990 152161 62002 152541
rect 62382 152161 62394 152541
rect 62774 152161 62786 152541
rect 63166 152161 63178 152541
rect 63558 152161 67916 152541
rect 60000 151998 67916 152161
rect 156052 152553 160442 152933
rect 160822 152553 160834 152933
rect 161214 152553 161226 152933
rect 161606 152553 161618 152933
rect 161998 152553 162010 152933
rect 162390 152553 162402 152933
rect 162782 152553 162794 152933
rect 163174 152553 163186 152933
rect 163566 152553 163578 152933
rect 163958 152553 164000 152933
rect 156052 152541 164000 152553
rect 156052 152161 160442 152541
rect 160822 152161 160834 152541
rect 161214 152161 161226 152541
rect 161606 152161 161618 152541
rect 161998 152161 162010 152541
rect 162390 152161 162402 152541
rect 162782 152161 162794 152541
rect 163174 152161 163186 152541
rect 163566 152161 163578 152541
rect 163958 152161 164000 152541
rect 156052 151998 164000 152161
rect 68316 151570 155652 151600
rect 68316 151190 68430 151570
rect 68810 151190 68822 151570
rect 69202 151190 75386 151570
rect 75766 151190 90506 151570
rect 90886 151190 105626 151570
rect 106006 151190 120746 151570
rect 121126 151190 135866 151570
rect 136246 151190 150986 151570
rect 151366 151190 154766 151570
rect 155146 151190 155158 151570
rect 155538 151190 155652 151570
rect 68316 151160 155652 151190
rect 71116 150330 152852 150360
rect 71116 149950 74146 150330
rect 74526 149950 89266 150330
rect 89646 149950 104386 150330
rect 104766 149950 119506 150330
rect 119886 149950 134626 150330
rect 135006 149950 149746 150330
rect 150126 149950 152852 150330
rect 71116 149920 152852 149950
rect 56000 149169 70716 149332
rect 56000 148789 56042 149169
rect 56422 148789 56434 149169
rect 56814 148789 56826 149169
rect 57206 148789 57218 149169
rect 57598 148789 57610 149169
rect 57990 148789 58002 149169
rect 58382 148789 58394 149169
rect 58774 148789 58786 149169
rect 59166 148789 59178 149169
rect 59558 148789 69830 149169
rect 70210 148789 70222 149169
rect 70602 148789 70716 149169
rect 56000 148777 70716 148789
rect 56000 148397 56042 148777
rect 56422 148397 56434 148777
rect 56814 148397 56826 148777
rect 57206 148397 57218 148777
rect 57598 148397 57610 148777
rect 57990 148397 58002 148777
rect 58382 148397 58394 148777
rect 58774 148397 58786 148777
rect 59166 148397 59178 148777
rect 59558 148397 69830 148777
rect 70210 148397 70222 148777
rect 70602 148397 70716 148777
rect 56000 148385 70716 148397
rect 56000 148005 56042 148385
rect 56422 148005 56434 148385
rect 56814 148005 56826 148385
rect 57206 148005 57218 148385
rect 57598 148005 57610 148385
rect 57990 148005 58002 148385
rect 58382 148005 58394 148385
rect 58774 148005 58786 148385
rect 59166 148005 59178 148385
rect 59558 148005 69830 148385
rect 70210 148005 70222 148385
rect 70602 148005 70716 148385
rect 56000 147993 70716 148005
rect 56000 147613 56042 147993
rect 56422 147613 56434 147993
rect 56814 147613 56826 147993
rect 57206 147613 57218 147993
rect 57598 147613 57610 147993
rect 57990 147613 58002 147993
rect 58382 147613 58394 147993
rect 58774 147613 58786 147993
rect 59166 147613 59178 147993
rect 59558 147613 69830 147993
rect 70210 147613 70222 147993
rect 70602 147613 70716 147993
rect 56000 147601 70716 147613
rect 56000 147221 56042 147601
rect 56422 147221 56434 147601
rect 56814 147221 56826 147601
rect 57206 147221 57218 147601
rect 57598 147221 57610 147601
rect 57990 147221 58002 147601
rect 58382 147221 58394 147601
rect 58774 147221 58786 147601
rect 59166 147221 59178 147601
rect 59558 147221 69830 147601
rect 70210 147221 70222 147601
rect 70602 147221 70716 147601
rect 56000 147209 70716 147221
rect 56000 146829 56042 147209
rect 56422 146829 56434 147209
rect 56814 146829 56826 147209
rect 57206 146829 57218 147209
rect 57598 146829 57610 147209
rect 57990 146829 58002 147209
rect 58382 146829 58394 147209
rect 58774 146829 58786 147209
rect 59166 146829 59178 147209
rect 59558 146829 69830 147209
rect 70210 146829 70222 147209
rect 70602 146829 70716 147209
rect 56000 146666 70716 146829
rect 153252 149169 168000 149332
rect 153252 148789 153366 149169
rect 153746 148789 153758 149169
rect 154138 148789 164442 149169
rect 164822 148789 164834 149169
rect 165214 148789 165226 149169
rect 165606 148789 165618 149169
rect 165998 148789 166010 149169
rect 166390 148789 166402 149169
rect 166782 148789 166794 149169
rect 167174 148789 167186 149169
rect 167566 148789 167578 149169
rect 167958 148789 168000 149169
rect 153252 148777 168000 148789
rect 153252 148397 153366 148777
rect 153746 148397 153758 148777
rect 154138 148397 164442 148777
rect 164822 148397 164834 148777
rect 165214 148397 165226 148777
rect 165606 148397 165618 148777
rect 165998 148397 166010 148777
rect 166390 148397 166402 148777
rect 166782 148397 166794 148777
rect 167174 148397 167186 148777
rect 167566 148397 167578 148777
rect 167958 148397 168000 148777
rect 153252 148385 168000 148397
rect 153252 148005 153366 148385
rect 153746 148005 153758 148385
rect 154138 148005 164442 148385
rect 164822 148005 164834 148385
rect 165214 148005 165226 148385
rect 165606 148005 165618 148385
rect 165998 148005 166010 148385
rect 166390 148005 166402 148385
rect 166782 148005 166794 148385
rect 167174 148005 167186 148385
rect 167566 148005 167578 148385
rect 167958 148005 168000 148385
rect 153252 147993 168000 148005
rect 153252 147613 153366 147993
rect 153746 147613 153758 147993
rect 154138 147613 164442 147993
rect 164822 147613 164834 147993
rect 165214 147613 165226 147993
rect 165606 147613 165618 147993
rect 165998 147613 166010 147993
rect 166390 147613 166402 147993
rect 166782 147613 166794 147993
rect 167174 147613 167186 147993
rect 167566 147613 167578 147993
rect 167958 147613 168000 147993
rect 153252 147601 168000 147613
rect 153252 147221 153366 147601
rect 153746 147221 153758 147601
rect 154138 147221 164442 147601
rect 164822 147221 164834 147601
rect 165214 147221 165226 147601
rect 165606 147221 165618 147601
rect 165998 147221 166010 147601
rect 166390 147221 166402 147601
rect 166782 147221 166794 147601
rect 167174 147221 167186 147601
rect 167566 147221 167578 147601
rect 167958 147221 168000 147601
rect 153252 147209 168000 147221
rect 153252 146829 153366 147209
rect 153746 146829 153758 147209
rect 154138 146829 164442 147209
rect 164822 146829 164834 147209
rect 165214 146829 165226 147209
rect 165606 146829 165618 147209
rect 165998 146829 166010 147209
rect 166390 146829 166402 147209
rect 166782 146829 166794 147209
rect 167174 146829 167186 147209
rect 167566 146829 167578 147209
rect 167958 146829 168000 147209
rect 153252 146666 168000 146829
rect 196000 145000 210000 159000
rect 14000 129000 28000 143000
rect 60000 138501 69316 138664
rect 60000 138121 60042 138501
rect 60422 138121 60434 138501
rect 60814 138121 60826 138501
rect 61206 138121 61218 138501
rect 61598 138121 61610 138501
rect 61990 138121 62002 138501
rect 62382 138121 62394 138501
rect 62774 138121 62786 138501
rect 63166 138121 63178 138501
rect 63558 138121 68430 138501
rect 68810 138121 68822 138501
rect 69202 138121 69316 138501
rect 60000 138109 69316 138121
rect 60000 137729 60042 138109
rect 60422 137729 60434 138109
rect 60814 137729 60826 138109
rect 61206 137729 61218 138109
rect 61598 137729 61610 138109
rect 61990 137729 62002 138109
rect 62382 137729 62394 138109
rect 62774 137729 62786 138109
rect 63166 137729 63178 138109
rect 63558 137729 68430 138109
rect 68810 137729 68822 138109
rect 69202 137729 69316 138109
rect 60000 137717 69316 137729
rect 60000 137337 60042 137717
rect 60422 137337 60434 137717
rect 60814 137337 60826 137717
rect 61206 137337 61218 137717
rect 61598 137337 61610 137717
rect 61990 137337 62002 137717
rect 62382 137337 62394 137717
rect 62774 137337 62786 137717
rect 63166 137337 63178 137717
rect 63558 137337 68430 137717
rect 68810 137337 68822 137717
rect 69202 137337 69316 137717
rect 60000 137325 69316 137337
rect 60000 136945 60042 137325
rect 60422 136945 60434 137325
rect 60814 136945 60826 137325
rect 61206 136945 61218 137325
rect 61598 136945 61610 137325
rect 61990 136945 62002 137325
rect 62382 136945 62394 137325
rect 62774 136945 62786 137325
rect 63166 136945 63178 137325
rect 63558 136945 68430 137325
rect 68810 136945 68822 137325
rect 69202 136945 69316 137325
rect 60000 136933 69316 136945
rect 60000 136553 60042 136933
rect 60422 136553 60434 136933
rect 60814 136553 60826 136933
rect 61206 136553 61218 136933
rect 61598 136553 61610 136933
rect 61990 136553 62002 136933
rect 62382 136553 62394 136933
rect 62774 136553 62786 136933
rect 63166 136553 63178 136933
rect 63558 136553 68430 136933
rect 68810 136553 68822 136933
rect 69202 136553 69316 136933
rect 60000 136541 69316 136553
rect 60000 136161 60042 136541
rect 60422 136161 60434 136541
rect 60814 136161 60826 136541
rect 61206 136161 61218 136541
rect 61598 136161 61610 136541
rect 61990 136161 62002 136541
rect 62382 136161 62394 136541
rect 62774 136161 62786 136541
rect 63166 136161 63178 136541
rect 63558 136161 68430 136541
rect 68810 136161 68822 136541
rect 69202 136161 69316 136541
rect 154652 138501 164000 138664
rect 154652 138121 154766 138501
rect 155146 138121 155158 138501
rect 155538 138121 160442 138501
rect 160822 138121 160834 138501
rect 161214 138121 161226 138501
rect 161606 138121 161618 138501
rect 161998 138121 162010 138501
rect 162390 138121 162402 138501
rect 162782 138121 162794 138501
rect 163174 138121 163186 138501
rect 163566 138121 163578 138501
rect 163958 138121 164000 138501
rect 154652 138109 164000 138121
rect 154652 137729 154766 138109
rect 155146 137729 155158 138109
rect 155538 137729 160442 138109
rect 160822 137729 160834 138109
rect 161214 137729 161226 138109
rect 161606 137729 161618 138109
rect 161998 137729 162010 138109
rect 162390 137729 162402 138109
rect 162782 137729 162794 138109
rect 163174 137729 163186 138109
rect 163566 137729 163578 138109
rect 163958 137729 164000 138109
rect 154652 137717 164000 137729
rect 154652 137337 154766 137717
rect 155146 137337 155158 137717
rect 155538 137337 160442 137717
rect 160822 137337 160834 137717
rect 161214 137337 161226 137717
rect 161606 137337 161618 137717
rect 161998 137337 162010 137717
rect 162390 137337 162402 137717
rect 162782 137337 162794 137717
rect 163174 137337 163186 137717
rect 163566 137337 163578 137717
rect 163958 137337 164000 137717
rect 154652 137325 164000 137337
rect 154652 136945 154766 137325
rect 155146 136945 155158 137325
rect 155538 136945 160442 137325
rect 160822 136945 160834 137325
rect 161214 136945 161226 137325
rect 161606 136945 161618 137325
rect 161998 136945 162010 137325
rect 162390 136945 162402 137325
rect 162782 136945 162794 137325
rect 163174 136945 163186 137325
rect 163566 136945 163578 137325
rect 163958 136945 164000 137325
rect 154652 136933 164000 136945
rect 154652 136553 154766 136933
rect 155146 136553 155158 136933
rect 155538 136553 160442 136933
rect 160822 136553 160834 136933
rect 161214 136553 161226 136933
rect 161606 136553 161618 136933
rect 161998 136553 162010 136933
rect 162390 136553 162402 136933
rect 162782 136553 162794 136933
rect 163174 136553 163186 136933
rect 163566 136553 163578 136933
rect 163958 136553 164000 136933
rect 154652 136541 164000 136553
rect 60000 135998 69316 136161
rect 69716 136450 154252 136480
rect 69716 136070 75386 136450
rect 75766 136070 90506 136450
rect 90886 136070 105626 136450
rect 106006 136070 120746 136450
rect 121126 136070 135866 136450
rect 136246 136070 150986 136450
rect 151366 136070 154252 136450
rect 69716 136040 154252 136070
rect 154652 136161 154766 136541
rect 155146 136161 155158 136541
rect 155538 136161 160442 136541
rect 160822 136161 160834 136541
rect 161214 136161 161226 136541
rect 161606 136161 161618 136541
rect 161998 136161 162010 136541
rect 162390 136161 162402 136541
rect 162782 136161 162794 136541
rect 163174 136161 163186 136541
rect 163566 136161 163578 136541
rect 163958 136161 164000 136541
rect 154652 135998 164000 136161
rect 69716 135210 154252 135240
rect 69716 134830 69830 135210
rect 70210 134830 70222 135210
rect 70602 134830 74146 135210
rect 74526 134830 89266 135210
rect 89646 134830 104386 135210
rect 104766 134830 119506 135210
rect 119886 134830 134626 135210
rect 135006 134830 149746 135210
rect 150126 134830 153366 135210
rect 153746 134830 153758 135210
rect 154138 134830 154252 135210
rect 69716 134800 154252 134830
rect 56000 133169 70716 133332
rect 56000 132789 56042 133169
rect 56422 132789 56434 133169
rect 56814 132789 56826 133169
rect 57206 132789 57218 133169
rect 57598 132789 57610 133169
rect 57990 132789 58002 133169
rect 58382 132789 58394 133169
rect 58774 132789 58786 133169
rect 59166 132789 59178 133169
rect 59558 132789 69830 133169
rect 70210 132789 70222 133169
rect 70602 132789 70716 133169
rect 56000 132777 70716 132789
rect 56000 132397 56042 132777
rect 56422 132397 56434 132777
rect 56814 132397 56826 132777
rect 57206 132397 57218 132777
rect 57598 132397 57610 132777
rect 57990 132397 58002 132777
rect 58382 132397 58394 132777
rect 58774 132397 58786 132777
rect 59166 132397 59178 132777
rect 59558 132397 69830 132777
rect 70210 132397 70222 132777
rect 70602 132397 70716 132777
rect 56000 132385 70716 132397
rect 56000 132005 56042 132385
rect 56422 132005 56434 132385
rect 56814 132005 56826 132385
rect 57206 132005 57218 132385
rect 57598 132005 57610 132385
rect 57990 132005 58002 132385
rect 58382 132005 58394 132385
rect 58774 132005 58786 132385
rect 59166 132005 59178 132385
rect 59558 132005 69830 132385
rect 70210 132005 70222 132385
rect 70602 132005 70716 132385
rect 56000 131993 70716 132005
rect 56000 131613 56042 131993
rect 56422 131613 56434 131993
rect 56814 131613 56826 131993
rect 57206 131613 57218 131993
rect 57598 131613 57610 131993
rect 57990 131613 58002 131993
rect 58382 131613 58394 131993
rect 58774 131613 58786 131993
rect 59166 131613 59178 131993
rect 59558 131613 69830 131993
rect 70210 131613 70222 131993
rect 70602 131613 70716 131993
rect 56000 131601 70716 131613
rect 56000 131221 56042 131601
rect 56422 131221 56434 131601
rect 56814 131221 56826 131601
rect 57206 131221 57218 131601
rect 57598 131221 57610 131601
rect 57990 131221 58002 131601
rect 58382 131221 58394 131601
rect 58774 131221 58786 131601
rect 59166 131221 59178 131601
rect 59558 131221 69830 131601
rect 70210 131221 70222 131601
rect 70602 131221 70716 131601
rect 56000 131209 70716 131221
rect 56000 130829 56042 131209
rect 56422 130829 56434 131209
rect 56814 130829 56826 131209
rect 57206 130829 57218 131209
rect 57598 130829 57610 131209
rect 57990 130829 58002 131209
rect 58382 130829 58394 131209
rect 58774 130829 58786 131209
rect 59166 130829 59178 131209
rect 59558 130829 69830 131209
rect 70210 130829 70222 131209
rect 70602 130829 70716 131209
rect 56000 130666 70716 130829
rect 153252 133169 168000 133332
rect 153252 132789 153366 133169
rect 153746 132789 153758 133169
rect 154138 132789 164442 133169
rect 164822 132789 164834 133169
rect 165214 132789 165226 133169
rect 165606 132789 165618 133169
rect 165998 132789 166010 133169
rect 166390 132789 166402 133169
rect 166782 132789 166794 133169
rect 167174 132789 167186 133169
rect 167566 132789 167578 133169
rect 167958 132789 168000 133169
rect 153252 132777 168000 132789
rect 153252 132397 153366 132777
rect 153746 132397 153758 132777
rect 154138 132397 164442 132777
rect 164822 132397 164834 132777
rect 165214 132397 165226 132777
rect 165606 132397 165618 132777
rect 165998 132397 166010 132777
rect 166390 132397 166402 132777
rect 166782 132397 166794 132777
rect 167174 132397 167186 132777
rect 167566 132397 167578 132777
rect 167958 132397 168000 132777
rect 153252 132385 168000 132397
rect 153252 132005 153366 132385
rect 153746 132005 153758 132385
rect 154138 132005 164442 132385
rect 164822 132005 164834 132385
rect 165214 132005 165226 132385
rect 165606 132005 165618 132385
rect 165998 132005 166010 132385
rect 166390 132005 166402 132385
rect 166782 132005 166794 132385
rect 167174 132005 167186 132385
rect 167566 132005 167578 132385
rect 167958 132005 168000 132385
rect 153252 131993 168000 132005
rect 153252 131613 153366 131993
rect 153746 131613 153758 131993
rect 154138 131613 164442 131993
rect 164822 131613 164834 131993
rect 165214 131613 165226 131993
rect 165606 131613 165618 131993
rect 165998 131613 166010 131993
rect 166390 131613 166402 131993
rect 166782 131613 166794 131993
rect 167174 131613 167186 131993
rect 167566 131613 167578 131993
rect 167958 131613 168000 131993
rect 153252 131601 168000 131613
rect 153252 131221 153366 131601
rect 153746 131221 153758 131601
rect 154138 131221 164442 131601
rect 164822 131221 164834 131601
rect 165214 131221 165226 131601
rect 165606 131221 165618 131601
rect 165998 131221 166010 131601
rect 166390 131221 166402 131601
rect 166782 131221 166794 131601
rect 167174 131221 167186 131601
rect 167566 131221 167578 131601
rect 167958 131221 168000 131601
rect 153252 131209 168000 131221
rect 153252 130829 153366 131209
rect 153746 130829 153758 131209
rect 154138 130829 164442 131209
rect 164822 130829 164834 131209
rect 165214 130829 165226 131209
rect 165606 130829 165618 131209
rect 165998 130829 166010 131209
rect 166390 130829 166402 131209
rect 166782 130829 166794 131209
rect 167174 130829 167186 131209
rect 167566 130829 167578 131209
rect 167958 130829 168000 131209
rect 153252 130666 168000 130829
rect 196000 129000 210000 143000
rect 14000 113000 28000 127000
rect 60000 122501 69316 122664
rect 60000 122121 60042 122501
rect 60422 122121 60434 122501
rect 60814 122121 60826 122501
rect 61206 122121 61218 122501
rect 61598 122121 61610 122501
rect 61990 122121 62002 122501
rect 62382 122121 62394 122501
rect 62774 122121 62786 122501
rect 63166 122121 63178 122501
rect 63558 122121 68430 122501
rect 68810 122121 68822 122501
rect 69202 122121 69316 122501
rect 60000 122109 69316 122121
rect 60000 121729 60042 122109
rect 60422 121729 60434 122109
rect 60814 121729 60826 122109
rect 61206 121729 61218 122109
rect 61598 121729 61610 122109
rect 61990 121729 62002 122109
rect 62382 121729 62394 122109
rect 62774 121729 62786 122109
rect 63166 121729 63178 122109
rect 63558 121729 68430 122109
rect 68810 121729 68822 122109
rect 69202 121729 69316 122109
rect 60000 121717 69316 121729
rect 60000 121337 60042 121717
rect 60422 121337 60434 121717
rect 60814 121337 60826 121717
rect 61206 121337 61218 121717
rect 61598 121337 61610 121717
rect 61990 121337 62002 121717
rect 62382 121337 62394 121717
rect 62774 121337 62786 121717
rect 63166 121337 63178 121717
rect 63558 121337 68430 121717
rect 68810 121337 68822 121717
rect 69202 121337 69316 121717
rect 154652 122501 164000 122664
rect 154652 122121 154766 122501
rect 155146 122121 155158 122501
rect 155538 122121 160442 122501
rect 160822 122121 160834 122501
rect 161214 122121 161226 122501
rect 161606 122121 161618 122501
rect 161998 122121 162010 122501
rect 162390 122121 162402 122501
rect 162782 122121 162794 122501
rect 163174 122121 163186 122501
rect 163566 122121 163578 122501
rect 163958 122121 164000 122501
rect 154652 122109 164000 122121
rect 154652 121729 154766 122109
rect 155146 121729 155158 122109
rect 155538 121729 160442 122109
rect 160822 121729 160834 122109
rect 161214 121729 161226 122109
rect 161606 121729 161618 122109
rect 161998 121729 162010 122109
rect 162390 121729 162402 122109
rect 162782 121729 162794 122109
rect 163174 121729 163186 122109
rect 163566 121729 163578 122109
rect 163958 121729 164000 122109
rect 154652 121717 164000 121729
rect 60000 121325 69316 121337
rect 60000 120945 60042 121325
rect 60422 120945 60434 121325
rect 60814 120945 60826 121325
rect 61206 120945 61218 121325
rect 61598 120945 61610 121325
rect 61990 120945 62002 121325
rect 62382 120945 62394 121325
rect 62774 120945 62786 121325
rect 63166 120945 63178 121325
rect 63558 120945 68430 121325
rect 68810 120945 68822 121325
rect 69202 120945 69316 121325
rect 60000 120933 69316 120945
rect 60000 120553 60042 120933
rect 60422 120553 60434 120933
rect 60814 120553 60826 120933
rect 61206 120553 61218 120933
rect 61598 120553 61610 120933
rect 61990 120553 62002 120933
rect 62382 120553 62394 120933
rect 62774 120553 62786 120933
rect 63166 120553 63178 120933
rect 63558 120553 68430 120933
rect 68810 120553 68822 120933
rect 69202 120553 69316 120933
rect 69716 121330 154252 121360
rect 69716 120950 75386 121330
rect 75766 120950 90506 121330
rect 90886 120950 105626 121330
rect 106006 120950 120746 121330
rect 121126 120950 135866 121330
rect 136246 120950 150986 121330
rect 151366 120950 154252 121330
rect 69716 120920 154252 120950
rect 154652 121337 154766 121717
rect 155146 121337 155158 121717
rect 155538 121337 160442 121717
rect 160822 121337 160834 121717
rect 161214 121337 161226 121717
rect 161606 121337 161618 121717
rect 161998 121337 162010 121717
rect 162390 121337 162402 121717
rect 162782 121337 162794 121717
rect 163174 121337 163186 121717
rect 163566 121337 163578 121717
rect 163958 121337 164000 121717
rect 154652 121325 164000 121337
rect 154652 120945 154766 121325
rect 155146 120945 155158 121325
rect 155538 120945 160442 121325
rect 160822 120945 160834 121325
rect 161214 120945 161226 121325
rect 161606 120945 161618 121325
rect 161998 120945 162010 121325
rect 162390 120945 162402 121325
rect 162782 120945 162794 121325
rect 163174 120945 163186 121325
rect 163566 120945 163578 121325
rect 163958 120945 164000 121325
rect 154652 120933 164000 120945
rect 60000 120541 69316 120553
rect 60000 120161 60042 120541
rect 60422 120161 60434 120541
rect 60814 120161 60826 120541
rect 61206 120161 61218 120541
rect 61598 120161 61610 120541
rect 61990 120161 62002 120541
rect 62382 120161 62394 120541
rect 62774 120161 62786 120541
rect 63166 120161 63178 120541
rect 63558 120161 68430 120541
rect 68810 120161 68822 120541
rect 69202 120161 69316 120541
rect 60000 119998 69316 120161
rect 154652 120553 154766 120933
rect 155146 120553 155158 120933
rect 155538 120553 160442 120933
rect 160822 120553 160834 120933
rect 161214 120553 161226 120933
rect 161606 120553 161618 120933
rect 161998 120553 162010 120933
rect 162390 120553 162402 120933
rect 162782 120553 162794 120933
rect 163174 120553 163186 120933
rect 163566 120553 163578 120933
rect 163958 120553 164000 120933
rect 154652 120541 164000 120553
rect 154652 120161 154766 120541
rect 155146 120161 155158 120541
rect 155538 120161 160442 120541
rect 160822 120161 160834 120541
rect 161214 120161 161226 120541
rect 161606 120161 161618 120541
rect 161998 120161 162010 120541
rect 162390 120161 162402 120541
rect 162782 120161 162794 120541
rect 163174 120161 163186 120541
rect 163566 120161 163578 120541
rect 163958 120161 164000 120541
rect 69716 120090 154252 120120
rect 69716 119710 69830 120090
rect 70210 119710 70222 120090
rect 70602 119710 74146 120090
rect 74526 119710 89266 120090
rect 89646 119710 104386 120090
rect 104766 119710 119506 120090
rect 119886 119710 134626 120090
rect 135006 119710 149746 120090
rect 150126 119710 153366 120090
rect 153746 119710 153758 120090
rect 154138 119710 154252 120090
rect 154652 119998 164000 120161
rect 69716 119680 154252 119710
rect 56000 117169 70716 117332
rect 56000 116789 56042 117169
rect 56422 116789 56434 117169
rect 56814 116789 56826 117169
rect 57206 116789 57218 117169
rect 57598 116789 57610 117169
rect 57990 116789 58002 117169
rect 58382 116789 58394 117169
rect 58774 116789 58786 117169
rect 59166 116789 59178 117169
rect 59558 116789 69830 117169
rect 70210 116789 70222 117169
rect 70602 116789 70716 117169
rect 56000 116777 70716 116789
rect 56000 116397 56042 116777
rect 56422 116397 56434 116777
rect 56814 116397 56826 116777
rect 57206 116397 57218 116777
rect 57598 116397 57610 116777
rect 57990 116397 58002 116777
rect 58382 116397 58394 116777
rect 58774 116397 58786 116777
rect 59166 116397 59178 116777
rect 59558 116397 69830 116777
rect 70210 116397 70222 116777
rect 70602 116397 70716 116777
rect 56000 116385 70716 116397
rect 56000 116005 56042 116385
rect 56422 116005 56434 116385
rect 56814 116005 56826 116385
rect 57206 116005 57218 116385
rect 57598 116005 57610 116385
rect 57990 116005 58002 116385
rect 58382 116005 58394 116385
rect 58774 116005 58786 116385
rect 59166 116005 59178 116385
rect 59558 116005 69830 116385
rect 70210 116005 70222 116385
rect 70602 116005 70716 116385
rect 56000 115993 70716 116005
rect 56000 115613 56042 115993
rect 56422 115613 56434 115993
rect 56814 115613 56826 115993
rect 57206 115613 57218 115993
rect 57598 115613 57610 115993
rect 57990 115613 58002 115993
rect 58382 115613 58394 115993
rect 58774 115613 58786 115993
rect 59166 115613 59178 115993
rect 59558 115613 69830 115993
rect 70210 115613 70222 115993
rect 70602 115613 70716 115993
rect 56000 115601 70716 115613
rect 56000 115221 56042 115601
rect 56422 115221 56434 115601
rect 56814 115221 56826 115601
rect 57206 115221 57218 115601
rect 57598 115221 57610 115601
rect 57990 115221 58002 115601
rect 58382 115221 58394 115601
rect 58774 115221 58786 115601
rect 59166 115221 59178 115601
rect 59558 115221 69830 115601
rect 70210 115221 70222 115601
rect 70602 115221 70716 115601
rect 56000 115209 70716 115221
rect 56000 114829 56042 115209
rect 56422 114829 56434 115209
rect 56814 114829 56826 115209
rect 57206 114829 57218 115209
rect 57598 114829 57610 115209
rect 57990 114829 58002 115209
rect 58382 114829 58394 115209
rect 58774 114829 58786 115209
rect 59166 114829 59178 115209
rect 59558 114829 69830 115209
rect 70210 114829 70222 115209
rect 70602 114829 70716 115209
rect 56000 114666 70716 114829
rect 153252 117169 168000 117332
rect 153252 116789 153366 117169
rect 153746 116789 153758 117169
rect 154138 116789 164442 117169
rect 164822 116789 164834 117169
rect 165214 116789 165226 117169
rect 165606 116789 165618 117169
rect 165998 116789 166010 117169
rect 166390 116789 166402 117169
rect 166782 116789 166794 117169
rect 167174 116789 167186 117169
rect 167566 116789 167578 117169
rect 167958 116789 168000 117169
rect 153252 116777 168000 116789
rect 153252 116397 153366 116777
rect 153746 116397 153758 116777
rect 154138 116397 164442 116777
rect 164822 116397 164834 116777
rect 165214 116397 165226 116777
rect 165606 116397 165618 116777
rect 165998 116397 166010 116777
rect 166390 116397 166402 116777
rect 166782 116397 166794 116777
rect 167174 116397 167186 116777
rect 167566 116397 167578 116777
rect 167958 116397 168000 116777
rect 153252 116385 168000 116397
rect 153252 116005 153366 116385
rect 153746 116005 153758 116385
rect 154138 116005 164442 116385
rect 164822 116005 164834 116385
rect 165214 116005 165226 116385
rect 165606 116005 165618 116385
rect 165998 116005 166010 116385
rect 166390 116005 166402 116385
rect 166782 116005 166794 116385
rect 167174 116005 167186 116385
rect 167566 116005 167578 116385
rect 167958 116005 168000 116385
rect 153252 115993 168000 116005
rect 153252 115613 153366 115993
rect 153746 115613 153758 115993
rect 154138 115613 164442 115993
rect 164822 115613 164834 115993
rect 165214 115613 165226 115993
rect 165606 115613 165618 115993
rect 165998 115613 166010 115993
rect 166390 115613 166402 115993
rect 166782 115613 166794 115993
rect 167174 115613 167186 115993
rect 167566 115613 167578 115993
rect 167958 115613 168000 115993
rect 153252 115601 168000 115613
rect 153252 115221 153366 115601
rect 153746 115221 153758 115601
rect 154138 115221 164442 115601
rect 164822 115221 164834 115601
rect 165214 115221 165226 115601
rect 165606 115221 165618 115601
rect 165998 115221 166010 115601
rect 166390 115221 166402 115601
rect 166782 115221 166794 115601
rect 167174 115221 167186 115601
rect 167566 115221 167578 115601
rect 167958 115221 168000 115601
rect 153252 115209 168000 115221
rect 153252 114829 153366 115209
rect 153746 114829 153758 115209
rect 154138 114829 164442 115209
rect 164822 114829 164834 115209
rect 165214 114829 165226 115209
rect 165606 114829 165618 115209
rect 165998 114829 166010 115209
rect 166390 114829 166402 115209
rect 166782 114829 166794 115209
rect 167174 114829 167186 115209
rect 167566 114829 167578 115209
rect 167958 114829 168000 115209
rect 153252 114666 168000 114829
rect 196000 113000 210000 127000
rect 14000 97000 28000 111000
rect 60000 106501 69316 106664
rect 60000 106121 60042 106501
rect 60422 106121 60434 106501
rect 60814 106121 60826 106501
rect 61206 106121 61218 106501
rect 61598 106121 61610 106501
rect 61990 106121 62002 106501
rect 62382 106121 62394 106501
rect 62774 106121 62786 106501
rect 63166 106121 63178 106501
rect 63558 106121 68430 106501
rect 68810 106121 68822 106501
rect 69202 106121 69316 106501
rect 154652 106501 164000 106664
rect 60000 106109 69316 106121
rect 60000 105729 60042 106109
rect 60422 105729 60434 106109
rect 60814 105729 60826 106109
rect 61206 105729 61218 106109
rect 61598 105729 61610 106109
rect 61990 105729 62002 106109
rect 62382 105729 62394 106109
rect 62774 105729 62786 106109
rect 63166 105729 63178 106109
rect 63558 105729 68430 106109
rect 68810 105729 68822 106109
rect 69202 105729 69316 106109
rect 69716 106210 154252 106240
rect 69716 105830 75386 106210
rect 75766 105830 90506 106210
rect 90886 105830 105626 106210
rect 106006 105830 120746 106210
rect 121126 105830 135866 106210
rect 136246 105830 150986 106210
rect 151366 105830 154252 106210
rect 69716 105800 154252 105830
rect 154652 106121 154766 106501
rect 155146 106121 155158 106501
rect 155538 106121 160442 106501
rect 160822 106121 160834 106501
rect 161214 106121 161226 106501
rect 161606 106121 161618 106501
rect 161998 106121 162010 106501
rect 162390 106121 162402 106501
rect 162782 106121 162794 106501
rect 163174 106121 163186 106501
rect 163566 106121 163578 106501
rect 163958 106121 164000 106501
rect 154652 106109 164000 106121
rect 60000 105717 69316 105729
rect 60000 105337 60042 105717
rect 60422 105337 60434 105717
rect 60814 105337 60826 105717
rect 61206 105337 61218 105717
rect 61598 105337 61610 105717
rect 61990 105337 62002 105717
rect 62382 105337 62394 105717
rect 62774 105337 62786 105717
rect 63166 105337 63178 105717
rect 63558 105337 68430 105717
rect 68810 105337 68822 105717
rect 69202 105337 69316 105717
rect 60000 105325 69316 105337
rect 60000 104945 60042 105325
rect 60422 104945 60434 105325
rect 60814 104945 60826 105325
rect 61206 104945 61218 105325
rect 61598 104945 61610 105325
rect 61990 104945 62002 105325
rect 62382 104945 62394 105325
rect 62774 104945 62786 105325
rect 63166 104945 63178 105325
rect 63558 104945 68430 105325
rect 68810 104945 68822 105325
rect 69202 104945 69316 105325
rect 154652 105729 154766 106109
rect 155146 105729 155158 106109
rect 155538 105729 160442 106109
rect 160822 105729 160834 106109
rect 161214 105729 161226 106109
rect 161606 105729 161618 106109
rect 161998 105729 162010 106109
rect 162390 105729 162402 106109
rect 162782 105729 162794 106109
rect 163174 105729 163186 106109
rect 163566 105729 163578 106109
rect 163958 105729 164000 106109
rect 154652 105717 164000 105729
rect 154652 105337 154766 105717
rect 155146 105337 155158 105717
rect 155538 105337 160442 105717
rect 160822 105337 160834 105717
rect 161214 105337 161226 105717
rect 161606 105337 161618 105717
rect 161998 105337 162010 105717
rect 162390 105337 162402 105717
rect 162782 105337 162794 105717
rect 163174 105337 163186 105717
rect 163566 105337 163578 105717
rect 163958 105337 164000 105717
rect 154652 105325 164000 105337
rect 60000 104933 69316 104945
rect 60000 104553 60042 104933
rect 60422 104553 60434 104933
rect 60814 104553 60826 104933
rect 61206 104553 61218 104933
rect 61598 104553 61610 104933
rect 61990 104553 62002 104933
rect 62382 104553 62394 104933
rect 62774 104553 62786 104933
rect 63166 104553 63178 104933
rect 63558 104553 68430 104933
rect 68810 104553 68822 104933
rect 69202 104553 69316 104933
rect 69716 104970 154252 105000
rect 69716 104590 69830 104970
rect 70210 104590 70222 104970
rect 70602 104590 74146 104970
rect 74526 104590 89266 104970
rect 89646 104590 104386 104970
rect 104766 104590 119506 104970
rect 119886 104590 134626 104970
rect 135006 104590 149746 104970
rect 150126 104590 153366 104970
rect 153746 104590 153758 104970
rect 154138 104590 154252 104970
rect 69716 104560 154252 104590
rect 154652 104945 154766 105325
rect 155146 104945 155158 105325
rect 155538 104945 160442 105325
rect 160822 104945 160834 105325
rect 161214 104945 161226 105325
rect 161606 104945 161618 105325
rect 161998 104945 162010 105325
rect 162390 104945 162402 105325
rect 162782 104945 162794 105325
rect 163174 104945 163186 105325
rect 163566 104945 163578 105325
rect 163958 104945 164000 105325
rect 154652 104933 164000 104945
rect 60000 104541 69316 104553
rect 60000 104161 60042 104541
rect 60422 104161 60434 104541
rect 60814 104161 60826 104541
rect 61206 104161 61218 104541
rect 61598 104161 61610 104541
rect 61990 104161 62002 104541
rect 62382 104161 62394 104541
rect 62774 104161 62786 104541
rect 63166 104161 63178 104541
rect 63558 104161 68430 104541
rect 68810 104161 68822 104541
rect 69202 104161 69316 104541
rect 60000 103998 69316 104161
rect 154652 104553 154766 104933
rect 155146 104553 155158 104933
rect 155538 104553 160442 104933
rect 160822 104553 160834 104933
rect 161214 104553 161226 104933
rect 161606 104553 161618 104933
rect 161998 104553 162010 104933
rect 162390 104553 162402 104933
rect 162782 104553 162794 104933
rect 163174 104553 163186 104933
rect 163566 104553 163578 104933
rect 163958 104553 164000 104933
rect 154652 104541 164000 104553
rect 154652 104161 154766 104541
rect 155146 104161 155158 104541
rect 155538 104161 160442 104541
rect 160822 104161 160834 104541
rect 161214 104161 161226 104541
rect 161606 104161 161618 104541
rect 161998 104161 162010 104541
rect 162390 104161 162402 104541
rect 162782 104161 162794 104541
rect 163174 104161 163186 104541
rect 163566 104161 163578 104541
rect 163958 104161 164000 104541
rect 154652 103998 164000 104161
rect 56000 101169 70716 101332
rect 56000 100789 56042 101169
rect 56422 100789 56434 101169
rect 56814 100789 56826 101169
rect 57206 100789 57218 101169
rect 57598 100789 57610 101169
rect 57990 100789 58002 101169
rect 58382 100789 58394 101169
rect 58774 100789 58786 101169
rect 59166 100789 59178 101169
rect 59558 100789 69830 101169
rect 70210 100789 70222 101169
rect 70602 100789 70716 101169
rect 56000 100777 70716 100789
rect 56000 100397 56042 100777
rect 56422 100397 56434 100777
rect 56814 100397 56826 100777
rect 57206 100397 57218 100777
rect 57598 100397 57610 100777
rect 57990 100397 58002 100777
rect 58382 100397 58394 100777
rect 58774 100397 58786 100777
rect 59166 100397 59178 100777
rect 59558 100397 69830 100777
rect 70210 100397 70222 100777
rect 70602 100397 70716 100777
rect 56000 100385 70716 100397
rect 56000 100005 56042 100385
rect 56422 100005 56434 100385
rect 56814 100005 56826 100385
rect 57206 100005 57218 100385
rect 57598 100005 57610 100385
rect 57990 100005 58002 100385
rect 58382 100005 58394 100385
rect 58774 100005 58786 100385
rect 59166 100005 59178 100385
rect 59558 100005 69830 100385
rect 70210 100005 70222 100385
rect 70602 100005 70716 100385
rect 56000 99993 70716 100005
rect 56000 99613 56042 99993
rect 56422 99613 56434 99993
rect 56814 99613 56826 99993
rect 57206 99613 57218 99993
rect 57598 99613 57610 99993
rect 57990 99613 58002 99993
rect 58382 99613 58394 99993
rect 58774 99613 58786 99993
rect 59166 99613 59178 99993
rect 59558 99613 69830 99993
rect 70210 99613 70222 99993
rect 70602 99613 70716 99993
rect 56000 99601 70716 99613
rect 56000 99221 56042 99601
rect 56422 99221 56434 99601
rect 56814 99221 56826 99601
rect 57206 99221 57218 99601
rect 57598 99221 57610 99601
rect 57990 99221 58002 99601
rect 58382 99221 58394 99601
rect 58774 99221 58786 99601
rect 59166 99221 59178 99601
rect 59558 99221 69830 99601
rect 70210 99221 70222 99601
rect 70602 99221 70716 99601
rect 56000 99209 70716 99221
rect 56000 98829 56042 99209
rect 56422 98829 56434 99209
rect 56814 98829 56826 99209
rect 57206 98829 57218 99209
rect 57598 98829 57610 99209
rect 57990 98829 58002 99209
rect 58382 98829 58394 99209
rect 58774 98829 58786 99209
rect 59166 98829 59178 99209
rect 59558 98829 69830 99209
rect 70210 98829 70222 99209
rect 70602 98829 70716 99209
rect 56000 98666 70716 98829
rect 153252 101169 168000 101332
rect 153252 100789 153366 101169
rect 153746 100789 153758 101169
rect 154138 100789 164442 101169
rect 164822 100789 164834 101169
rect 165214 100789 165226 101169
rect 165606 100789 165618 101169
rect 165998 100789 166010 101169
rect 166390 100789 166402 101169
rect 166782 100789 166794 101169
rect 167174 100789 167186 101169
rect 167566 100789 167578 101169
rect 167958 100789 168000 101169
rect 153252 100777 168000 100789
rect 153252 100397 153366 100777
rect 153746 100397 153758 100777
rect 154138 100397 164442 100777
rect 164822 100397 164834 100777
rect 165214 100397 165226 100777
rect 165606 100397 165618 100777
rect 165998 100397 166010 100777
rect 166390 100397 166402 100777
rect 166782 100397 166794 100777
rect 167174 100397 167186 100777
rect 167566 100397 167578 100777
rect 167958 100397 168000 100777
rect 153252 100385 168000 100397
rect 153252 100005 153366 100385
rect 153746 100005 153758 100385
rect 154138 100005 164442 100385
rect 164822 100005 164834 100385
rect 165214 100005 165226 100385
rect 165606 100005 165618 100385
rect 165998 100005 166010 100385
rect 166390 100005 166402 100385
rect 166782 100005 166794 100385
rect 167174 100005 167186 100385
rect 167566 100005 167578 100385
rect 167958 100005 168000 100385
rect 153252 99993 168000 100005
rect 153252 99613 153366 99993
rect 153746 99613 153758 99993
rect 154138 99613 164442 99993
rect 164822 99613 164834 99993
rect 165214 99613 165226 99993
rect 165606 99613 165618 99993
rect 165998 99613 166010 99993
rect 166390 99613 166402 99993
rect 166782 99613 166794 99993
rect 167174 99613 167186 99993
rect 167566 99613 167578 99993
rect 167958 99613 168000 99993
rect 153252 99601 168000 99613
rect 153252 99221 153366 99601
rect 153746 99221 153758 99601
rect 154138 99221 164442 99601
rect 164822 99221 164834 99601
rect 165214 99221 165226 99601
rect 165606 99221 165618 99601
rect 165998 99221 166010 99601
rect 166390 99221 166402 99601
rect 166782 99221 166794 99601
rect 167174 99221 167186 99601
rect 167566 99221 167578 99601
rect 167958 99221 168000 99601
rect 153252 99209 168000 99221
rect 153252 98829 153366 99209
rect 153746 98829 153758 99209
rect 154138 98829 164442 99209
rect 164822 98829 164834 99209
rect 165214 98829 165226 99209
rect 165606 98829 165618 99209
rect 165998 98829 166010 99209
rect 166390 98829 166402 99209
rect 166782 98829 166794 99209
rect 167174 98829 167186 99209
rect 167566 98829 167578 99209
rect 167958 98829 168000 99209
rect 153252 98666 168000 98829
rect 196000 97000 210000 111000
rect 14000 81000 28000 95000
rect 69716 91090 154252 91120
rect 69716 90710 75386 91090
rect 75766 90710 90506 91090
rect 90886 90710 105626 91090
rect 106006 90710 120746 91090
rect 121126 90710 135866 91090
rect 136246 90710 150986 91090
rect 151366 90710 154252 91090
rect 69716 90680 154252 90710
rect 60000 90501 69316 90664
rect 60000 90121 60042 90501
rect 60422 90121 60434 90501
rect 60814 90121 60826 90501
rect 61206 90121 61218 90501
rect 61598 90121 61610 90501
rect 61990 90121 62002 90501
rect 62382 90121 62394 90501
rect 62774 90121 62786 90501
rect 63166 90121 63178 90501
rect 63558 90121 68430 90501
rect 68810 90121 68822 90501
rect 69202 90121 69316 90501
rect 60000 90109 69316 90121
rect 60000 89729 60042 90109
rect 60422 89729 60434 90109
rect 60814 89729 60826 90109
rect 61206 89729 61218 90109
rect 61598 89729 61610 90109
rect 61990 89729 62002 90109
rect 62382 89729 62394 90109
rect 62774 89729 62786 90109
rect 63166 89729 63178 90109
rect 63558 89729 68430 90109
rect 68810 89729 68822 90109
rect 69202 89729 69316 90109
rect 154652 90501 164000 90664
rect 154652 90121 154766 90501
rect 155146 90121 155158 90501
rect 155538 90121 160442 90501
rect 160822 90121 160834 90501
rect 161214 90121 161226 90501
rect 161606 90121 161618 90501
rect 161998 90121 162010 90501
rect 162390 90121 162402 90501
rect 162782 90121 162794 90501
rect 163174 90121 163186 90501
rect 163566 90121 163578 90501
rect 163958 90121 164000 90501
rect 154652 90109 164000 90121
rect 60000 89717 69316 89729
rect 60000 89337 60042 89717
rect 60422 89337 60434 89717
rect 60814 89337 60826 89717
rect 61206 89337 61218 89717
rect 61598 89337 61610 89717
rect 61990 89337 62002 89717
rect 62382 89337 62394 89717
rect 62774 89337 62786 89717
rect 63166 89337 63178 89717
rect 63558 89337 68430 89717
rect 68810 89337 68822 89717
rect 69202 89337 69316 89717
rect 69716 89850 154252 89880
rect 69716 89470 69830 89850
rect 70210 89470 70222 89850
rect 70602 89470 74146 89850
rect 74526 89470 89266 89850
rect 89646 89470 104386 89850
rect 104766 89470 119506 89850
rect 119886 89470 134626 89850
rect 135006 89470 149746 89850
rect 150126 89470 153366 89850
rect 153746 89470 153758 89850
rect 154138 89470 154252 89850
rect 69716 89440 154252 89470
rect 154652 89729 154766 90109
rect 155146 89729 155158 90109
rect 155538 89729 160442 90109
rect 160822 89729 160834 90109
rect 161214 89729 161226 90109
rect 161606 89729 161618 90109
rect 161998 89729 162010 90109
rect 162390 89729 162402 90109
rect 162782 89729 162794 90109
rect 163174 89729 163186 90109
rect 163566 89729 163578 90109
rect 163958 89729 164000 90109
rect 154652 89717 164000 89729
rect 60000 89325 69316 89337
rect 60000 88945 60042 89325
rect 60422 88945 60434 89325
rect 60814 88945 60826 89325
rect 61206 88945 61218 89325
rect 61598 88945 61610 89325
rect 61990 88945 62002 89325
rect 62382 88945 62394 89325
rect 62774 88945 62786 89325
rect 63166 88945 63178 89325
rect 63558 88945 68430 89325
rect 68810 88945 68822 89325
rect 69202 88945 69316 89325
rect 60000 88933 69316 88945
rect 60000 88553 60042 88933
rect 60422 88553 60434 88933
rect 60814 88553 60826 88933
rect 61206 88553 61218 88933
rect 61598 88553 61610 88933
rect 61990 88553 62002 88933
rect 62382 88553 62394 88933
rect 62774 88553 62786 88933
rect 63166 88553 63178 88933
rect 63558 88553 68430 88933
rect 68810 88553 68822 88933
rect 69202 88553 69316 88933
rect 60000 88541 69316 88553
rect 60000 88161 60042 88541
rect 60422 88161 60434 88541
rect 60814 88161 60826 88541
rect 61206 88161 61218 88541
rect 61598 88161 61610 88541
rect 61990 88161 62002 88541
rect 62382 88161 62394 88541
rect 62774 88161 62786 88541
rect 63166 88161 63178 88541
rect 63558 88161 68430 88541
rect 68810 88161 68822 88541
rect 69202 88161 69316 88541
rect 60000 87998 69316 88161
rect 154652 89337 154766 89717
rect 155146 89337 155158 89717
rect 155538 89337 160442 89717
rect 160822 89337 160834 89717
rect 161214 89337 161226 89717
rect 161606 89337 161618 89717
rect 161998 89337 162010 89717
rect 162390 89337 162402 89717
rect 162782 89337 162794 89717
rect 163174 89337 163186 89717
rect 163566 89337 163578 89717
rect 163958 89337 164000 89717
rect 154652 89325 164000 89337
rect 154652 88945 154766 89325
rect 155146 88945 155158 89325
rect 155538 88945 160442 89325
rect 160822 88945 160834 89325
rect 161214 88945 161226 89325
rect 161606 88945 161618 89325
rect 161998 88945 162010 89325
rect 162390 88945 162402 89325
rect 162782 88945 162794 89325
rect 163174 88945 163186 89325
rect 163566 88945 163578 89325
rect 163958 88945 164000 89325
rect 154652 88933 164000 88945
rect 154652 88553 154766 88933
rect 155146 88553 155158 88933
rect 155538 88553 160442 88933
rect 160822 88553 160834 88933
rect 161214 88553 161226 88933
rect 161606 88553 161618 88933
rect 161998 88553 162010 88933
rect 162390 88553 162402 88933
rect 162782 88553 162794 88933
rect 163174 88553 163186 88933
rect 163566 88553 163578 88933
rect 163958 88553 164000 88933
rect 154652 88541 164000 88553
rect 154652 88161 154766 88541
rect 155146 88161 155158 88541
rect 155538 88161 160442 88541
rect 160822 88161 160834 88541
rect 161214 88161 161226 88541
rect 161606 88161 161618 88541
rect 161998 88161 162010 88541
rect 162390 88161 162402 88541
rect 162782 88161 162794 88541
rect 163174 88161 163186 88541
rect 163566 88161 163578 88541
rect 163958 88161 164000 88541
rect 154652 87998 164000 88161
rect 56000 85169 70716 85332
rect 56000 84789 56042 85169
rect 56422 84789 56434 85169
rect 56814 84789 56826 85169
rect 57206 84789 57218 85169
rect 57598 84789 57610 85169
rect 57990 84789 58002 85169
rect 58382 84789 58394 85169
rect 58774 84789 58786 85169
rect 59166 84789 59178 85169
rect 59558 84789 69830 85169
rect 70210 84789 70222 85169
rect 70602 84789 70716 85169
rect 56000 84777 70716 84789
rect 56000 84397 56042 84777
rect 56422 84397 56434 84777
rect 56814 84397 56826 84777
rect 57206 84397 57218 84777
rect 57598 84397 57610 84777
rect 57990 84397 58002 84777
rect 58382 84397 58394 84777
rect 58774 84397 58786 84777
rect 59166 84397 59178 84777
rect 59558 84397 69830 84777
rect 70210 84397 70222 84777
rect 70602 84397 70716 84777
rect 56000 84385 70716 84397
rect 56000 84005 56042 84385
rect 56422 84005 56434 84385
rect 56814 84005 56826 84385
rect 57206 84005 57218 84385
rect 57598 84005 57610 84385
rect 57990 84005 58002 84385
rect 58382 84005 58394 84385
rect 58774 84005 58786 84385
rect 59166 84005 59178 84385
rect 59558 84005 69830 84385
rect 70210 84005 70222 84385
rect 70602 84005 70716 84385
rect 56000 83993 70716 84005
rect 56000 83613 56042 83993
rect 56422 83613 56434 83993
rect 56814 83613 56826 83993
rect 57206 83613 57218 83993
rect 57598 83613 57610 83993
rect 57990 83613 58002 83993
rect 58382 83613 58394 83993
rect 58774 83613 58786 83993
rect 59166 83613 59178 83993
rect 59558 83613 69830 83993
rect 70210 83613 70222 83993
rect 70602 83613 70716 83993
rect 56000 83601 70716 83613
rect 56000 83221 56042 83601
rect 56422 83221 56434 83601
rect 56814 83221 56826 83601
rect 57206 83221 57218 83601
rect 57598 83221 57610 83601
rect 57990 83221 58002 83601
rect 58382 83221 58394 83601
rect 58774 83221 58786 83601
rect 59166 83221 59178 83601
rect 59558 83221 69830 83601
rect 70210 83221 70222 83601
rect 70602 83221 70716 83601
rect 56000 83209 70716 83221
rect 56000 82829 56042 83209
rect 56422 82829 56434 83209
rect 56814 82829 56826 83209
rect 57206 82829 57218 83209
rect 57598 82829 57610 83209
rect 57990 82829 58002 83209
rect 58382 82829 58394 83209
rect 58774 82829 58786 83209
rect 59166 82829 59178 83209
rect 59558 82829 69830 83209
rect 70210 82829 70222 83209
rect 70602 82829 70716 83209
rect 56000 82666 70716 82829
rect 153252 85169 168000 85332
rect 153252 84789 153366 85169
rect 153746 84789 153758 85169
rect 154138 84789 164442 85169
rect 164822 84789 164834 85169
rect 165214 84789 165226 85169
rect 165606 84789 165618 85169
rect 165998 84789 166010 85169
rect 166390 84789 166402 85169
rect 166782 84789 166794 85169
rect 167174 84789 167186 85169
rect 167566 84789 167578 85169
rect 167958 84789 168000 85169
rect 153252 84777 168000 84789
rect 153252 84397 153366 84777
rect 153746 84397 153758 84777
rect 154138 84397 164442 84777
rect 164822 84397 164834 84777
rect 165214 84397 165226 84777
rect 165606 84397 165618 84777
rect 165998 84397 166010 84777
rect 166390 84397 166402 84777
rect 166782 84397 166794 84777
rect 167174 84397 167186 84777
rect 167566 84397 167578 84777
rect 167958 84397 168000 84777
rect 153252 84385 168000 84397
rect 153252 84005 153366 84385
rect 153746 84005 153758 84385
rect 154138 84005 164442 84385
rect 164822 84005 164834 84385
rect 165214 84005 165226 84385
rect 165606 84005 165618 84385
rect 165998 84005 166010 84385
rect 166390 84005 166402 84385
rect 166782 84005 166794 84385
rect 167174 84005 167186 84385
rect 167566 84005 167578 84385
rect 167958 84005 168000 84385
rect 153252 83993 168000 84005
rect 153252 83613 153366 83993
rect 153746 83613 153758 83993
rect 154138 83613 164442 83993
rect 164822 83613 164834 83993
rect 165214 83613 165226 83993
rect 165606 83613 165618 83993
rect 165998 83613 166010 83993
rect 166390 83613 166402 83993
rect 166782 83613 166794 83993
rect 167174 83613 167186 83993
rect 167566 83613 167578 83993
rect 167958 83613 168000 83993
rect 153252 83601 168000 83613
rect 153252 83221 153366 83601
rect 153746 83221 153758 83601
rect 154138 83221 164442 83601
rect 164822 83221 164834 83601
rect 165214 83221 165226 83601
rect 165606 83221 165618 83601
rect 165998 83221 166010 83601
rect 166390 83221 166402 83601
rect 166782 83221 166794 83601
rect 167174 83221 167186 83601
rect 167566 83221 167578 83601
rect 167958 83221 168000 83601
rect 153252 83209 168000 83221
rect 153252 82829 153366 83209
rect 153746 82829 153758 83209
rect 154138 82829 164442 83209
rect 164822 82829 164834 83209
rect 165214 82829 165226 83209
rect 165606 82829 165618 83209
rect 165998 82829 166010 83209
rect 166390 82829 166402 83209
rect 166782 82829 166794 83209
rect 167174 82829 167186 83209
rect 167566 82829 167578 83209
rect 167958 82829 168000 83209
rect 153252 82666 168000 82829
rect 196000 81000 210000 95000
rect 14000 65000 28000 79000
rect 68316 75970 155652 76000
rect 68316 75590 68430 75970
rect 68810 75590 68822 75970
rect 69202 75590 75386 75970
rect 75766 75590 90506 75970
rect 90886 75590 105626 75970
rect 106006 75590 120746 75970
rect 121126 75590 135866 75970
rect 136246 75590 150986 75970
rect 151366 75590 154766 75970
rect 155146 75590 155158 75970
rect 155538 75590 155652 75970
rect 68316 75560 155652 75590
rect 69716 74730 154252 74760
rect 60000 74501 69316 74664
rect 60000 74121 60042 74501
rect 60422 74121 60434 74501
rect 60814 74121 60826 74501
rect 61206 74121 61218 74501
rect 61598 74121 61610 74501
rect 61990 74121 62002 74501
rect 62382 74121 62394 74501
rect 62774 74121 62786 74501
rect 63166 74121 63178 74501
rect 63558 74121 68430 74501
rect 68810 74121 68822 74501
rect 69202 74121 69316 74501
rect 69716 74350 69830 74730
rect 70210 74350 70222 74730
rect 70602 74350 74146 74730
rect 74526 74350 89266 74730
rect 89646 74350 104386 74730
rect 104766 74350 119506 74730
rect 119886 74350 134626 74730
rect 135006 74350 149746 74730
rect 150126 74350 153366 74730
rect 153746 74350 153758 74730
rect 154138 74350 154252 74730
rect 69716 74320 154252 74350
rect 154652 74501 164000 74664
rect 60000 74109 69316 74121
rect 60000 73729 60042 74109
rect 60422 73729 60434 74109
rect 60814 73729 60826 74109
rect 61206 73729 61218 74109
rect 61598 73729 61610 74109
rect 61990 73729 62002 74109
rect 62382 73729 62394 74109
rect 62774 73729 62786 74109
rect 63166 73729 63178 74109
rect 63558 73729 68430 74109
rect 68810 73729 68822 74109
rect 69202 73729 69316 74109
rect 60000 73717 69316 73729
rect 60000 73337 60042 73717
rect 60422 73337 60434 73717
rect 60814 73337 60826 73717
rect 61206 73337 61218 73717
rect 61598 73337 61610 73717
rect 61990 73337 62002 73717
rect 62382 73337 62394 73717
rect 62774 73337 62786 73717
rect 63166 73337 63178 73717
rect 63558 73337 68430 73717
rect 68810 73337 68822 73717
rect 69202 73337 69316 73717
rect 60000 73325 69316 73337
rect 60000 72945 60042 73325
rect 60422 72945 60434 73325
rect 60814 72945 60826 73325
rect 61206 72945 61218 73325
rect 61598 72945 61610 73325
rect 61990 72945 62002 73325
rect 62382 72945 62394 73325
rect 62774 72945 62786 73325
rect 63166 72945 63178 73325
rect 63558 72945 68430 73325
rect 68810 72945 68822 73325
rect 69202 72945 69316 73325
rect 60000 72933 69316 72945
rect 60000 72553 60042 72933
rect 60422 72553 60434 72933
rect 60814 72553 60826 72933
rect 61206 72553 61218 72933
rect 61598 72553 61610 72933
rect 61990 72553 62002 72933
rect 62382 72553 62394 72933
rect 62774 72553 62786 72933
rect 63166 72553 63178 72933
rect 63558 72553 68430 72933
rect 68810 72553 68822 72933
rect 69202 72553 69316 72933
rect 60000 72541 69316 72553
rect 60000 72161 60042 72541
rect 60422 72161 60434 72541
rect 60814 72161 60826 72541
rect 61206 72161 61218 72541
rect 61598 72161 61610 72541
rect 61990 72161 62002 72541
rect 62382 72161 62394 72541
rect 62774 72161 62786 72541
rect 63166 72161 63178 72541
rect 63558 72161 68430 72541
rect 68810 72161 68822 72541
rect 69202 72161 69316 72541
rect 60000 71998 69316 72161
rect 154652 74121 154766 74501
rect 155146 74121 155158 74501
rect 155538 74121 160442 74501
rect 160822 74121 160834 74501
rect 161214 74121 161226 74501
rect 161606 74121 161618 74501
rect 161998 74121 162010 74501
rect 162390 74121 162402 74501
rect 162782 74121 162794 74501
rect 163174 74121 163186 74501
rect 163566 74121 163578 74501
rect 163958 74121 164000 74501
rect 154652 74109 164000 74121
rect 154652 73729 154766 74109
rect 155146 73729 155158 74109
rect 155538 73729 160442 74109
rect 160822 73729 160834 74109
rect 161214 73729 161226 74109
rect 161606 73729 161618 74109
rect 161998 73729 162010 74109
rect 162390 73729 162402 74109
rect 162782 73729 162794 74109
rect 163174 73729 163186 74109
rect 163566 73729 163578 74109
rect 163958 73729 164000 74109
rect 154652 73717 164000 73729
rect 154652 73337 154766 73717
rect 155146 73337 155158 73717
rect 155538 73337 160442 73717
rect 160822 73337 160834 73717
rect 161214 73337 161226 73717
rect 161606 73337 161618 73717
rect 161998 73337 162010 73717
rect 162390 73337 162402 73717
rect 162782 73337 162794 73717
rect 163174 73337 163186 73717
rect 163566 73337 163578 73717
rect 163958 73337 164000 73717
rect 154652 73325 164000 73337
rect 154652 72945 154766 73325
rect 155146 72945 155158 73325
rect 155538 72945 160442 73325
rect 160822 72945 160834 73325
rect 161214 72945 161226 73325
rect 161606 72945 161618 73325
rect 161998 72945 162010 73325
rect 162390 72945 162402 73325
rect 162782 72945 162794 73325
rect 163174 72945 163186 73325
rect 163566 72945 163578 73325
rect 163958 72945 164000 73325
rect 154652 72933 164000 72945
rect 154652 72553 154766 72933
rect 155146 72553 155158 72933
rect 155538 72553 160442 72933
rect 160822 72553 160834 72933
rect 161214 72553 161226 72933
rect 161606 72553 161618 72933
rect 161998 72553 162010 72933
rect 162390 72553 162402 72933
rect 162782 72553 162794 72933
rect 163174 72553 163186 72933
rect 163566 72553 163578 72933
rect 163958 72553 164000 72933
rect 154652 72541 164000 72553
rect 154652 72161 154766 72541
rect 155146 72161 155158 72541
rect 155538 72161 160442 72541
rect 160822 72161 160834 72541
rect 161214 72161 161226 72541
rect 161606 72161 161618 72541
rect 161998 72161 162010 72541
rect 162390 72161 162402 72541
rect 162782 72161 162794 72541
rect 163174 72161 163186 72541
rect 163566 72161 163578 72541
rect 163958 72161 164000 72541
rect 154652 71998 164000 72161
rect 69716 70806 154252 70920
rect 69716 70426 69830 70806
rect 70210 70426 70222 70806
rect 70602 70426 74146 70806
rect 74526 70426 89266 70806
rect 89646 70426 104386 70806
rect 104766 70426 119506 70806
rect 119886 70426 134626 70806
rect 135006 70426 149746 70806
rect 150126 70426 153366 70806
rect 153746 70426 153758 70806
rect 154138 70426 154252 70806
rect 69716 70414 154252 70426
rect 69716 70034 69830 70414
rect 70210 70034 70222 70414
rect 70602 70034 74146 70414
rect 74526 70034 89266 70414
rect 89646 70034 104386 70414
rect 104766 70034 119506 70414
rect 119886 70034 134626 70414
rect 135006 70034 149746 70414
rect 150126 70034 153366 70414
rect 153746 70034 153758 70414
rect 154138 70034 154252 70414
rect 69716 69920 154252 70034
rect 68316 69406 155652 69520
rect 68316 69026 68430 69406
rect 68810 69026 68822 69406
rect 69202 69026 75386 69406
rect 75766 69026 90506 69406
rect 90886 69026 105626 69406
rect 106006 69026 120746 69406
rect 121126 69026 135866 69406
rect 136246 69026 150986 69406
rect 151366 69026 154766 69406
rect 155146 69026 155158 69406
rect 155538 69026 155652 69406
rect 68316 69014 155652 69026
rect 68316 68634 68430 69014
rect 68810 68634 68822 69014
rect 69202 68634 75386 69014
rect 75766 68634 90506 69014
rect 90886 68634 105626 69014
rect 106006 68634 120746 69014
rect 121126 68634 135866 69014
rect 136246 68634 150986 69014
rect 151366 68634 154766 69014
rect 155146 68634 155158 69014
rect 155538 68634 155652 69014
rect 68316 68520 155652 68634
rect 71998 63558 74664 68120
rect 71998 63178 72161 63558
rect 72541 63178 72553 63558
rect 72933 63178 72945 63558
rect 73325 63178 73337 63558
rect 73717 63178 73729 63558
rect 74109 63178 74121 63558
rect 74501 63178 74664 63558
rect 71998 63166 74664 63178
rect 71998 62786 72161 63166
rect 72541 62786 72553 63166
rect 72933 62786 72945 63166
rect 73325 62786 73337 63166
rect 73717 62786 73729 63166
rect 74109 62786 74121 63166
rect 74501 62786 74664 63166
rect 71998 62774 74664 62786
rect 71998 62394 72161 62774
rect 72541 62394 72553 62774
rect 72933 62394 72945 62774
rect 73325 62394 73337 62774
rect 73717 62394 73729 62774
rect 74109 62394 74121 62774
rect 74501 62394 74664 62774
rect 71998 62382 74664 62394
rect 71998 62002 72161 62382
rect 72541 62002 72553 62382
rect 72933 62002 72945 62382
rect 73325 62002 73337 62382
rect 73717 62002 73729 62382
rect 74109 62002 74121 62382
rect 74501 62002 74664 62382
rect 71998 61990 74664 62002
rect 71998 61610 72161 61990
rect 72541 61610 72553 61990
rect 72933 61610 72945 61990
rect 73325 61610 73337 61990
rect 73717 61610 73729 61990
rect 74109 61610 74121 61990
rect 74501 61610 74664 61990
rect 71998 61598 74664 61610
rect 71998 61218 72161 61598
rect 72541 61218 72553 61598
rect 72933 61218 72945 61598
rect 73325 61218 73337 61598
rect 73717 61218 73729 61598
rect 74109 61218 74121 61598
rect 74501 61218 74664 61598
rect 71998 61206 74664 61218
rect 71998 60826 72161 61206
rect 72541 60826 72553 61206
rect 72933 60826 72945 61206
rect 73325 60826 73337 61206
rect 73717 60826 73729 61206
rect 74109 60826 74121 61206
rect 74501 60826 74664 61206
rect 71998 60814 74664 60826
rect 71998 60434 72161 60814
rect 72541 60434 72553 60814
rect 72933 60434 72945 60814
rect 73325 60434 73337 60814
rect 73717 60434 73729 60814
rect 74109 60434 74121 60814
rect 74501 60434 74664 60814
rect 71998 60422 74664 60434
rect 71998 60042 72161 60422
rect 72541 60042 72553 60422
rect 72933 60042 72945 60422
rect 73325 60042 73337 60422
rect 73717 60042 73729 60422
rect 74109 60042 74121 60422
rect 74501 60042 74664 60422
rect 71998 60000 74664 60042
rect 82666 59558 85332 68120
rect 87998 63558 90664 68120
rect 87998 63178 88161 63558
rect 88541 63178 88553 63558
rect 88933 63178 88945 63558
rect 89325 63178 89337 63558
rect 89717 63178 89729 63558
rect 90109 63178 90121 63558
rect 90501 63178 90664 63558
rect 87998 63166 90664 63178
rect 87998 62786 88161 63166
rect 88541 62786 88553 63166
rect 88933 62786 88945 63166
rect 89325 62786 89337 63166
rect 89717 62786 89729 63166
rect 90109 62786 90121 63166
rect 90501 62786 90664 63166
rect 87998 62774 90664 62786
rect 87998 62394 88161 62774
rect 88541 62394 88553 62774
rect 88933 62394 88945 62774
rect 89325 62394 89337 62774
rect 89717 62394 89729 62774
rect 90109 62394 90121 62774
rect 90501 62394 90664 62774
rect 87998 62382 90664 62394
rect 87998 62002 88161 62382
rect 88541 62002 88553 62382
rect 88933 62002 88945 62382
rect 89325 62002 89337 62382
rect 89717 62002 89729 62382
rect 90109 62002 90121 62382
rect 90501 62002 90664 62382
rect 87998 61990 90664 62002
rect 87998 61610 88161 61990
rect 88541 61610 88553 61990
rect 88933 61610 88945 61990
rect 89325 61610 89337 61990
rect 89717 61610 89729 61990
rect 90109 61610 90121 61990
rect 90501 61610 90664 61990
rect 87998 61598 90664 61610
rect 87998 61218 88161 61598
rect 88541 61218 88553 61598
rect 88933 61218 88945 61598
rect 89325 61218 89337 61598
rect 89717 61218 89729 61598
rect 90109 61218 90121 61598
rect 90501 61218 90664 61598
rect 87998 61206 90664 61218
rect 87998 60826 88161 61206
rect 88541 60826 88553 61206
rect 88933 60826 88945 61206
rect 89325 60826 89337 61206
rect 89717 60826 89729 61206
rect 90109 60826 90121 61206
rect 90501 60826 90664 61206
rect 87998 60814 90664 60826
rect 87998 60434 88161 60814
rect 88541 60434 88553 60814
rect 88933 60434 88945 60814
rect 89325 60434 89337 60814
rect 89717 60434 89729 60814
rect 90109 60434 90121 60814
rect 90501 60434 90664 60814
rect 87998 60422 90664 60434
rect 87998 60042 88161 60422
rect 88541 60042 88553 60422
rect 88933 60042 88945 60422
rect 89325 60042 89337 60422
rect 89717 60042 89729 60422
rect 90109 60042 90121 60422
rect 90501 60042 90664 60422
rect 87998 60000 90664 60042
rect 82666 59178 82829 59558
rect 83209 59178 83221 59558
rect 83601 59178 83613 59558
rect 83993 59178 84005 59558
rect 84385 59178 84397 59558
rect 84777 59178 84789 59558
rect 85169 59178 85332 59558
rect 82666 59166 85332 59178
rect 82666 58786 82829 59166
rect 83209 58786 83221 59166
rect 83601 58786 83613 59166
rect 83993 58786 84005 59166
rect 84385 58786 84397 59166
rect 84777 58786 84789 59166
rect 85169 58786 85332 59166
rect 82666 58774 85332 58786
rect 82666 58394 82829 58774
rect 83209 58394 83221 58774
rect 83601 58394 83613 58774
rect 83993 58394 84005 58774
rect 84385 58394 84397 58774
rect 84777 58394 84789 58774
rect 85169 58394 85332 58774
rect 82666 58382 85332 58394
rect 82666 58002 82829 58382
rect 83209 58002 83221 58382
rect 83601 58002 83613 58382
rect 83993 58002 84005 58382
rect 84385 58002 84397 58382
rect 84777 58002 84789 58382
rect 85169 58002 85332 58382
rect 82666 57990 85332 58002
rect 82666 57610 82829 57990
rect 83209 57610 83221 57990
rect 83601 57610 83613 57990
rect 83993 57610 84005 57990
rect 84385 57610 84397 57990
rect 84777 57610 84789 57990
rect 85169 57610 85332 57990
rect 82666 57598 85332 57610
rect 82666 57218 82829 57598
rect 83209 57218 83221 57598
rect 83601 57218 83613 57598
rect 83993 57218 84005 57598
rect 84385 57218 84397 57598
rect 84777 57218 84789 57598
rect 85169 57218 85332 57598
rect 82666 57206 85332 57218
rect 82666 56826 82829 57206
rect 83209 56826 83221 57206
rect 83601 56826 83613 57206
rect 83993 56826 84005 57206
rect 84385 56826 84397 57206
rect 84777 56826 84789 57206
rect 85169 56826 85332 57206
rect 82666 56814 85332 56826
rect 82666 56434 82829 56814
rect 83209 56434 83221 56814
rect 83601 56434 83613 56814
rect 83993 56434 84005 56814
rect 84385 56434 84397 56814
rect 84777 56434 84789 56814
rect 85169 56434 85332 56814
rect 82666 56422 85332 56434
rect 82666 56042 82829 56422
rect 83209 56042 83221 56422
rect 83601 56042 83613 56422
rect 83993 56042 84005 56422
rect 84385 56042 84397 56422
rect 84777 56042 84789 56422
rect 85169 56042 85332 56422
rect 82666 56000 85332 56042
rect 98666 59558 101332 68120
rect 103998 63558 106664 68120
rect 103998 63178 104161 63558
rect 104541 63178 104553 63558
rect 104933 63178 104945 63558
rect 105325 63178 105337 63558
rect 105717 63178 105729 63558
rect 106109 63178 106121 63558
rect 106501 63178 106664 63558
rect 103998 63166 106664 63178
rect 103998 62786 104161 63166
rect 104541 62786 104553 63166
rect 104933 62786 104945 63166
rect 105325 62786 105337 63166
rect 105717 62786 105729 63166
rect 106109 62786 106121 63166
rect 106501 62786 106664 63166
rect 103998 62774 106664 62786
rect 103998 62394 104161 62774
rect 104541 62394 104553 62774
rect 104933 62394 104945 62774
rect 105325 62394 105337 62774
rect 105717 62394 105729 62774
rect 106109 62394 106121 62774
rect 106501 62394 106664 62774
rect 103998 62382 106664 62394
rect 103998 62002 104161 62382
rect 104541 62002 104553 62382
rect 104933 62002 104945 62382
rect 105325 62002 105337 62382
rect 105717 62002 105729 62382
rect 106109 62002 106121 62382
rect 106501 62002 106664 62382
rect 103998 61990 106664 62002
rect 103998 61610 104161 61990
rect 104541 61610 104553 61990
rect 104933 61610 104945 61990
rect 105325 61610 105337 61990
rect 105717 61610 105729 61990
rect 106109 61610 106121 61990
rect 106501 61610 106664 61990
rect 103998 61598 106664 61610
rect 103998 61218 104161 61598
rect 104541 61218 104553 61598
rect 104933 61218 104945 61598
rect 105325 61218 105337 61598
rect 105717 61218 105729 61598
rect 106109 61218 106121 61598
rect 106501 61218 106664 61598
rect 103998 61206 106664 61218
rect 103998 60826 104161 61206
rect 104541 60826 104553 61206
rect 104933 60826 104945 61206
rect 105325 60826 105337 61206
rect 105717 60826 105729 61206
rect 106109 60826 106121 61206
rect 106501 60826 106664 61206
rect 103998 60814 106664 60826
rect 103998 60434 104161 60814
rect 104541 60434 104553 60814
rect 104933 60434 104945 60814
rect 105325 60434 105337 60814
rect 105717 60434 105729 60814
rect 106109 60434 106121 60814
rect 106501 60434 106664 60814
rect 103998 60422 106664 60434
rect 103998 60042 104161 60422
rect 104541 60042 104553 60422
rect 104933 60042 104945 60422
rect 105325 60042 105337 60422
rect 105717 60042 105729 60422
rect 106109 60042 106121 60422
rect 106501 60042 106664 60422
rect 103998 60000 106664 60042
rect 98666 59178 98829 59558
rect 99209 59178 99221 59558
rect 99601 59178 99613 59558
rect 99993 59178 100005 59558
rect 100385 59178 100397 59558
rect 100777 59178 100789 59558
rect 101169 59178 101332 59558
rect 98666 59166 101332 59178
rect 98666 58786 98829 59166
rect 99209 58786 99221 59166
rect 99601 58786 99613 59166
rect 99993 58786 100005 59166
rect 100385 58786 100397 59166
rect 100777 58786 100789 59166
rect 101169 58786 101332 59166
rect 98666 58774 101332 58786
rect 98666 58394 98829 58774
rect 99209 58394 99221 58774
rect 99601 58394 99613 58774
rect 99993 58394 100005 58774
rect 100385 58394 100397 58774
rect 100777 58394 100789 58774
rect 101169 58394 101332 58774
rect 98666 58382 101332 58394
rect 98666 58002 98829 58382
rect 99209 58002 99221 58382
rect 99601 58002 99613 58382
rect 99993 58002 100005 58382
rect 100385 58002 100397 58382
rect 100777 58002 100789 58382
rect 101169 58002 101332 58382
rect 98666 57990 101332 58002
rect 98666 57610 98829 57990
rect 99209 57610 99221 57990
rect 99601 57610 99613 57990
rect 99993 57610 100005 57990
rect 100385 57610 100397 57990
rect 100777 57610 100789 57990
rect 101169 57610 101332 57990
rect 98666 57598 101332 57610
rect 98666 57218 98829 57598
rect 99209 57218 99221 57598
rect 99601 57218 99613 57598
rect 99993 57218 100005 57598
rect 100385 57218 100397 57598
rect 100777 57218 100789 57598
rect 101169 57218 101332 57598
rect 98666 57206 101332 57218
rect 98666 56826 98829 57206
rect 99209 56826 99221 57206
rect 99601 56826 99613 57206
rect 99993 56826 100005 57206
rect 100385 56826 100397 57206
rect 100777 56826 100789 57206
rect 101169 56826 101332 57206
rect 98666 56814 101332 56826
rect 98666 56434 98829 56814
rect 99209 56434 99221 56814
rect 99601 56434 99613 56814
rect 99993 56434 100005 56814
rect 100385 56434 100397 56814
rect 100777 56434 100789 56814
rect 101169 56434 101332 56814
rect 98666 56422 101332 56434
rect 98666 56042 98829 56422
rect 99209 56042 99221 56422
rect 99601 56042 99613 56422
rect 99993 56042 100005 56422
rect 100385 56042 100397 56422
rect 100777 56042 100789 56422
rect 101169 56042 101332 56422
rect 98666 56000 101332 56042
rect 114666 59558 117332 68120
rect 119998 63558 122664 68120
rect 119998 63178 120161 63558
rect 120541 63178 120553 63558
rect 120933 63178 120945 63558
rect 121325 63178 121337 63558
rect 121717 63178 121729 63558
rect 122109 63178 122121 63558
rect 122501 63178 122664 63558
rect 119998 63166 122664 63178
rect 119998 62786 120161 63166
rect 120541 62786 120553 63166
rect 120933 62786 120945 63166
rect 121325 62786 121337 63166
rect 121717 62786 121729 63166
rect 122109 62786 122121 63166
rect 122501 62786 122664 63166
rect 119998 62774 122664 62786
rect 119998 62394 120161 62774
rect 120541 62394 120553 62774
rect 120933 62394 120945 62774
rect 121325 62394 121337 62774
rect 121717 62394 121729 62774
rect 122109 62394 122121 62774
rect 122501 62394 122664 62774
rect 119998 62382 122664 62394
rect 119998 62002 120161 62382
rect 120541 62002 120553 62382
rect 120933 62002 120945 62382
rect 121325 62002 121337 62382
rect 121717 62002 121729 62382
rect 122109 62002 122121 62382
rect 122501 62002 122664 62382
rect 119998 61990 122664 62002
rect 119998 61610 120161 61990
rect 120541 61610 120553 61990
rect 120933 61610 120945 61990
rect 121325 61610 121337 61990
rect 121717 61610 121729 61990
rect 122109 61610 122121 61990
rect 122501 61610 122664 61990
rect 119998 61598 122664 61610
rect 119998 61218 120161 61598
rect 120541 61218 120553 61598
rect 120933 61218 120945 61598
rect 121325 61218 121337 61598
rect 121717 61218 121729 61598
rect 122109 61218 122121 61598
rect 122501 61218 122664 61598
rect 119998 61206 122664 61218
rect 119998 60826 120161 61206
rect 120541 60826 120553 61206
rect 120933 60826 120945 61206
rect 121325 60826 121337 61206
rect 121717 60826 121729 61206
rect 122109 60826 122121 61206
rect 122501 60826 122664 61206
rect 119998 60814 122664 60826
rect 119998 60434 120161 60814
rect 120541 60434 120553 60814
rect 120933 60434 120945 60814
rect 121325 60434 121337 60814
rect 121717 60434 121729 60814
rect 122109 60434 122121 60814
rect 122501 60434 122664 60814
rect 119998 60422 122664 60434
rect 119998 60042 120161 60422
rect 120541 60042 120553 60422
rect 120933 60042 120945 60422
rect 121325 60042 121337 60422
rect 121717 60042 121729 60422
rect 122109 60042 122121 60422
rect 122501 60042 122664 60422
rect 119998 60000 122664 60042
rect 132000 63558 136000 68120
rect 132000 63178 132046 63558
rect 132426 63178 132438 63558
rect 132818 63178 132830 63558
rect 133210 63178 133222 63558
rect 133602 63178 133614 63558
rect 133994 63178 134006 63558
rect 134386 63178 134398 63558
rect 134778 63178 134790 63558
rect 135170 63178 135182 63558
rect 135562 63178 135574 63558
rect 135954 63178 136000 63558
rect 132000 63166 136000 63178
rect 132000 62786 132046 63166
rect 132426 62786 132438 63166
rect 132818 62786 132830 63166
rect 133210 62786 133222 63166
rect 133602 62786 133614 63166
rect 133994 62786 134006 63166
rect 134386 62786 134398 63166
rect 134778 62786 134790 63166
rect 135170 62786 135182 63166
rect 135562 62786 135574 63166
rect 135954 62786 136000 63166
rect 132000 62774 136000 62786
rect 132000 62394 132046 62774
rect 132426 62394 132438 62774
rect 132818 62394 132830 62774
rect 133210 62394 133222 62774
rect 133602 62394 133614 62774
rect 133994 62394 134006 62774
rect 134386 62394 134398 62774
rect 134778 62394 134790 62774
rect 135170 62394 135182 62774
rect 135562 62394 135574 62774
rect 135954 62394 136000 62774
rect 132000 62382 136000 62394
rect 132000 62002 132046 62382
rect 132426 62002 132438 62382
rect 132818 62002 132830 62382
rect 133210 62002 133222 62382
rect 133602 62002 133614 62382
rect 133994 62002 134006 62382
rect 134386 62002 134398 62382
rect 134778 62002 134790 62382
rect 135170 62002 135182 62382
rect 135562 62002 135574 62382
rect 135954 62002 136000 62382
rect 132000 61990 136000 62002
rect 132000 61610 132046 61990
rect 132426 61610 132438 61990
rect 132818 61610 132830 61990
rect 133210 61610 133222 61990
rect 133602 61610 133614 61990
rect 133994 61610 134006 61990
rect 134386 61610 134398 61990
rect 134778 61610 134790 61990
rect 135170 61610 135182 61990
rect 135562 61610 135574 61990
rect 135954 61610 136000 61990
rect 132000 61598 136000 61610
rect 132000 61218 132046 61598
rect 132426 61218 132438 61598
rect 132818 61218 132830 61598
rect 133210 61218 133222 61598
rect 133602 61218 133614 61598
rect 133994 61218 134006 61598
rect 134386 61218 134398 61598
rect 134778 61218 134790 61598
rect 135170 61218 135182 61598
rect 135562 61218 135574 61598
rect 135954 61218 136000 61598
rect 132000 61206 136000 61218
rect 132000 60826 132046 61206
rect 132426 60826 132438 61206
rect 132818 60826 132830 61206
rect 133210 60826 133222 61206
rect 133602 60826 133614 61206
rect 133994 60826 134006 61206
rect 134386 60826 134398 61206
rect 134778 60826 134790 61206
rect 135170 60826 135182 61206
rect 135562 60826 135574 61206
rect 135954 60826 136000 61206
rect 132000 60814 136000 60826
rect 132000 60434 132046 60814
rect 132426 60434 132438 60814
rect 132818 60434 132830 60814
rect 133210 60434 133222 60814
rect 133602 60434 133614 60814
rect 133994 60434 134006 60814
rect 134386 60434 134398 60814
rect 134778 60434 134790 60814
rect 135170 60434 135182 60814
rect 135562 60434 135574 60814
rect 135954 60434 136000 60814
rect 132000 60422 136000 60434
rect 132000 60042 132046 60422
rect 132426 60042 132438 60422
rect 132818 60042 132830 60422
rect 133210 60042 133222 60422
rect 133602 60042 133614 60422
rect 133994 60042 134006 60422
rect 134386 60042 134398 60422
rect 134778 60042 134790 60422
rect 135170 60042 135182 60422
rect 135562 60042 135574 60422
rect 135954 60042 136000 60422
rect 132000 60000 136000 60042
rect 114666 59178 114829 59558
rect 115209 59178 115221 59558
rect 115601 59178 115613 59558
rect 115993 59178 116005 59558
rect 116385 59178 116397 59558
rect 116777 59178 116789 59558
rect 117169 59178 117332 59558
rect 114666 59166 117332 59178
rect 114666 58786 114829 59166
rect 115209 58786 115221 59166
rect 115601 58786 115613 59166
rect 115993 58786 116005 59166
rect 116385 58786 116397 59166
rect 116777 58786 116789 59166
rect 117169 58786 117332 59166
rect 114666 58774 117332 58786
rect 114666 58394 114829 58774
rect 115209 58394 115221 58774
rect 115601 58394 115613 58774
rect 115993 58394 116005 58774
rect 116385 58394 116397 58774
rect 116777 58394 116789 58774
rect 117169 58394 117332 58774
rect 114666 58382 117332 58394
rect 114666 58002 114829 58382
rect 115209 58002 115221 58382
rect 115601 58002 115613 58382
rect 115993 58002 116005 58382
rect 116385 58002 116397 58382
rect 116777 58002 116789 58382
rect 117169 58002 117332 58382
rect 114666 57990 117332 58002
rect 114666 57610 114829 57990
rect 115209 57610 115221 57990
rect 115601 57610 115613 57990
rect 115993 57610 116005 57990
rect 116385 57610 116397 57990
rect 116777 57610 116789 57990
rect 117169 57610 117332 57990
rect 114666 57598 117332 57610
rect 114666 57218 114829 57598
rect 115209 57218 115221 57598
rect 115601 57218 115613 57598
rect 115993 57218 116005 57598
rect 116385 57218 116397 57598
rect 116777 57218 116789 57598
rect 117169 57218 117332 57598
rect 114666 57206 117332 57218
rect 114666 56826 114829 57206
rect 115209 56826 115221 57206
rect 115601 56826 115613 57206
rect 115993 56826 116005 57206
rect 116385 56826 116397 57206
rect 116777 56826 116789 57206
rect 117169 56826 117332 57206
rect 114666 56814 117332 56826
rect 114666 56434 114829 56814
rect 115209 56434 115221 56814
rect 115601 56434 115613 56814
rect 115993 56434 116005 56814
rect 116385 56434 116397 56814
rect 116777 56434 116789 56814
rect 117169 56434 117332 56814
rect 114666 56422 117332 56434
rect 114666 56042 114829 56422
rect 115209 56042 115221 56422
rect 115601 56042 115613 56422
rect 115993 56042 116005 56422
rect 116385 56042 116397 56422
rect 116777 56042 116789 56422
rect 117169 56042 117332 56422
rect 114666 56000 117332 56042
rect 146666 59558 149332 68120
rect 151998 63558 154664 68120
rect 196000 65000 210000 79000
rect 151998 63178 152161 63558
rect 152541 63178 152553 63558
rect 152933 63178 152945 63558
rect 153325 63178 153337 63558
rect 153717 63178 153729 63558
rect 154109 63178 154121 63558
rect 154501 63178 154664 63558
rect 151998 63166 154664 63178
rect 151998 62786 152161 63166
rect 152541 62786 152553 63166
rect 152933 62786 152945 63166
rect 153325 62786 153337 63166
rect 153717 62786 153729 63166
rect 154109 62786 154121 63166
rect 154501 62786 154664 63166
rect 151998 62774 154664 62786
rect 151998 62394 152161 62774
rect 152541 62394 152553 62774
rect 152933 62394 152945 62774
rect 153325 62394 153337 62774
rect 153717 62394 153729 62774
rect 154109 62394 154121 62774
rect 154501 62394 154664 62774
rect 151998 62382 154664 62394
rect 151998 62002 152161 62382
rect 152541 62002 152553 62382
rect 152933 62002 152945 62382
rect 153325 62002 153337 62382
rect 153717 62002 153729 62382
rect 154109 62002 154121 62382
rect 154501 62002 154664 62382
rect 151998 61990 154664 62002
rect 151998 61610 152161 61990
rect 152541 61610 152553 61990
rect 152933 61610 152945 61990
rect 153325 61610 153337 61990
rect 153717 61610 153729 61990
rect 154109 61610 154121 61990
rect 154501 61610 154664 61990
rect 151998 61598 154664 61610
rect 151998 61218 152161 61598
rect 152541 61218 152553 61598
rect 152933 61218 152945 61598
rect 153325 61218 153337 61598
rect 153717 61218 153729 61598
rect 154109 61218 154121 61598
rect 154501 61218 154664 61598
rect 151998 61206 154664 61218
rect 151998 60826 152161 61206
rect 152541 60826 152553 61206
rect 152933 60826 152945 61206
rect 153325 60826 153337 61206
rect 153717 60826 153729 61206
rect 154109 60826 154121 61206
rect 154501 60826 154664 61206
rect 151998 60814 154664 60826
rect 151998 60434 152161 60814
rect 152541 60434 152553 60814
rect 152933 60434 152945 60814
rect 153325 60434 153337 60814
rect 153717 60434 153729 60814
rect 154109 60434 154121 60814
rect 154501 60434 154664 60814
rect 151998 60422 154664 60434
rect 151998 60042 152161 60422
rect 152541 60042 152553 60422
rect 152933 60042 152945 60422
rect 153325 60042 153337 60422
rect 153717 60042 153729 60422
rect 154109 60042 154121 60422
rect 154501 60042 154664 60422
rect 151998 60000 154664 60042
rect 146666 59178 146829 59558
rect 147209 59178 147221 59558
rect 147601 59178 147613 59558
rect 147993 59178 148005 59558
rect 148385 59178 148397 59558
rect 148777 59178 148789 59558
rect 149169 59178 149332 59558
rect 146666 59166 149332 59178
rect 146666 58786 146829 59166
rect 147209 58786 147221 59166
rect 147601 58786 147613 59166
rect 147993 58786 148005 59166
rect 148385 58786 148397 59166
rect 148777 58786 148789 59166
rect 149169 58786 149332 59166
rect 146666 58774 149332 58786
rect 146666 58394 146829 58774
rect 147209 58394 147221 58774
rect 147601 58394 147613 58774
rect 147993 58394 148005 58774
rect 148385 58394 148397 58774
rect 148777 58394 148789 58774
rect 149169 58394 149332 58774
rect 146666 58382 149332 58394
rect 146666 58002 146829 58382
rect 147209 58002 147221 58382
rect 147601 58002 147613 58382
rect 147993 58002 148005 58382
rect 148385 58002 148397 58382
rect 148777 58002 148789 58382
rect 149169 58002 149332 58382
rect 146666 57990 149332 58002
rect 146666 57610 146829 57990
rect 147209 57610 147221 57990
rect 147601 57610 147613 57990
rect 147993 57610 148005 57990
rect 148385 57610 148397 57990
rect 148777 57610 148789 57990
rect 149169 57610 149332 57990
rect 146666 57598 149332 57610
rect 146666 57218 146829 57598
rect 147209 57218 147221 57598
rect 147601 57218 147613 57598
rect 147993 57218 148005 57598
rect 148385 57218 148397 57598
rect 148777 57218 148789 57598
rect 149169 57218 149332 57598
rect 146666 57206 149332 57218
rect 146666 56826 146829 57206
rect 147209 56826 147221 57206
rect 147601 56826 147613 57206
rect 147993 56826 148005 57206
rect 148385 56826 148397 57206
rect 148777 56826 148789 57206
rect 149169 56826 149332 57206
rect 146666 56814 149332 56826
rect 146666 56434 146829 56814
rect 147209 56434 147221 56814
rect 147601 56434 147613 56814
rect 147993 56434 148005 56814
rect 148385 56434 148397 56814
rect 148777 56434 148789 56814
rect 149169 56434 149332 56814
rect 146666 56422 149332 56434
rect 146666 56042 146829 56422
rect 147209 56042 147221 56422
rect 147601 56042 147613 56422
rect 147993 56042 148005 56422
rect 148385 56042 148397 56422
rect 148777 56042 148789 56422
rect 149169 56042 149332 56422
rect 146666 56000 149332 56042
rect 65000 14000 79000 28000
rect 81000 14000 95000 28000
rect 97000 14000 111000 28000
rect 113000 14000 127000 28000
rect 129000 14000 143000 28000
rect 145000 14000 159000 28000
use sg13g2_decap_8  FILLER_0_0
timestamp 1679581782
transform 1 0 71616 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679581782
transform 1 0 72288 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679581782
transform 1 0 72960 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679581782
transform 1 0 73632 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679581782
transform 1 0 74304 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679581782
transform 1 0 74976 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679581782
transform 1 0 75648 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679581782
transform 1 0 76320 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679581782
transform 1 0 76992 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679581782
transform 1 0 77664 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679581782
transform 1 0 78336 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679581782
transform 1 0 79008 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679581782
transform 1 0 79680 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679581782
transform 1 0 80352 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679581782
transform 1 0 81024 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679581782
transform 1 0 81696 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679581782
transform 1 0 82368 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679581782
transform 1 0 83040 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679581782
transform 1 0 83712 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679581782
transform 1 0 84384 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679581782
transform 1 0 85056 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679581782
transform 1 0 85728 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679581782
transform 1 0 86400 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679581782
transform 1 0 87072 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679581782
transform 1 0 87744 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679581782
transform 1 0 88416 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679581782
transform 1 0 89088 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679581782
transform 1 0 89760 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679581782
transform 1 0 90432 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679581782
transform 1 0 91104 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679581782
transform 1 0 91776 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679581782
transform 1 0 92448 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679581782
transform 1 0 93120 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679581782
transform 1 0 93792 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679581782
transform 1 0 94464 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679581782
transform 1 0 95136 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679581782
transform 1 0 95808 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679581782
transform 1 0 96480 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679581782
transform 1 0 97152 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679581782
transform 1 0 97824 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679581782
transform 1 0 98496 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679581782
transform 1 0 99168 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679581782
transform 1 0 99840 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679581782
transform 1 0 100512 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679581782
transform 1 0 101184 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679581782
transform 1 0 101856 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679581782
transform 1 0 102528 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679581782
transform 1 0 103200 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679581782
transform 1 0 103872 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679581782
transform 1 0 104544 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679581782
transform 1 0 105216 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679581782
transform 1 0 105888 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679581782
transform 1 0 106560 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679581782
transform 1 0 107232 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679581782
transform 1 0 107904 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679581782
transform 1 0 108576 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679581782
transform 1 0 109248 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679581782
transform 1 0 109920 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679581782
transform 1 0 110592 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679581782
transform 1 0 111264 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679581782
transform 1 0 111936 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679581782
transform 1 0 112608 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679581782
transform 1 0 113280 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679581782
transform 1 0 113952 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679581782
transform 1 0 114624 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679581782
transform 1 0 115296 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679581782
transform 1 0 115968 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679581782
transform 1 0 116640 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679581782
transform 1 0 117312 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679581782
transform 1 0 117984 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679581782
transform 1 0 118656 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679581782
transform 1 0 119328 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679581782
transform 1 0 120000 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679581782
transform 1 0 120672 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679581782
transform 1 0 121344 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679581782
transform 1 0 122016 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679581782
transform 1 0 122688 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679581782
transform 1 0 123360 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679581782
transform 1 0 124032 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679581782
transform 1 0 124704 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679581782
transform 1 0 125376 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679581782
transform 1 0 126048 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679581782
transform 1 0 126720 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679581782
transform 1 0 127392 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679581782
transform 1 0 128064 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679581782
transform 1 0 128736 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679581782
transform 1 0 129408 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679581782
transform 1 0 130080 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679581782
transform 1 0 130752 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679581782
transform 1 0 131424 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679581782
transform 1 0 132096 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679581782
transform 1 0 132768 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679581782
transform 1 0 133440 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679581782
transform 1 0 134112 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679581782
transform 1 0 134784 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679581782
transform 1 0 135456 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679581782
transform 1 0 136128 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679581782
transform 1 0 136800 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679581782
transform 1 0 137472 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679581782
transform 1 0 138144 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679581782
transform 1 0 138816 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679581782
transform 1 0 139488 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679581782
transform 1 0 140160 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679581782
transform 1 0 140832 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679581782
transform 1 0 141504 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679581782
transform 1 0 142176 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679581782
transform 1 0 142848 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_749
timestamp 1679581782
transform 1 0 143520 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_756
timestamp 1679581782
transform 1 0 144192 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_763
timestamp 1679581782
transform 1 0 144864 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_770
timestamp 1679581782
transform 1 0 145536 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_777
timestamp 1679581782
transform 1 0 146208 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_784
timestamp 1679581782
transform 1 0 146880 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_791
timestamp 1679581782
transform 1 0 147552 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_798
timestamp 1679581782
transform 1 0 148224 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_805
timestamp 1679581782
transform 1 0 148896 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_812
timestamp 1679581782
transform 1 0 149568 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_819
timestamp 1679581782
transform 1 0 150240 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_826
timestamp 1679581782
transform 1 0 150912 0 1 71820
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_833
timestamp 1679581782
transform 1 0 151584 0 1 71820
box -48 -56 720 834
use sg13g2_fill_1  FILLER_0_840
timestamp 1677579658
transform 1 0 152256 0 1 71820
box -48 -56 144 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679581782
transform 1 0 71616 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679581782
transform 1 0 72288 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679581782
transform 1 0 72960 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679581782
transform 1 0 73632 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679581782
transform 1 0 74304 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679581782
transform 1 0 74976 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679581782
transform 1 0 75648 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679581782
transform 1 0 76320 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679581782
transform 1 0 76992 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679581782
transform 1 0 77664 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679581782
transform 1 0 78336 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679581782
transform 1 0 79008 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679581782
transform 1 0 79680 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679581782
transform 1 0 80352 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679581782
transform 1 0 81024 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679581782
transform 1 0 81696 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679581782
transform 1 0 82368 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679581782
transform 1 0 83040 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679581782
transform 1 0 83712 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679581782
transform 1 0 84384 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679581782
transform 1 0 85056 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679581782
transform 1 0 85728 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679581782
transform 1 0 86400 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679581782
transform 1 0 87072 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679581782
transform 1 0 87744 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679581782
transform 1 0 88416 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679581782
transform 1 0 89088 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679581782
transform 1 0 89760 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 90432 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679581782
transform 1 0 91104 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679581782
transform 1 0 91776 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679581782
transform 1 0 92448 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679581782
transform 1 0 93120 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679581782
transform 1 0 93792 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679581782
transform 1 0 94464 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679581782
transform 1 0 95136 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679581782
transform 1 0 95808 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679581782
transform 1 0 96480 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679581782
transform 1 0 97152 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679581782
transform 1 0 97824 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679581782
transform 1 0 98496 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679581782
transform 1 0 99168 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679581782
transform 1 0 99840 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679581782
transform 1 0 100512 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679581782
transform 1 0 101184 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679581782
transform 1 0 101856 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679581782
transform 1 0 102528 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679581782
transform 1 0 103200 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679581782
transform 1 0 103872 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679581782
transform 1 0 104544 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679581782
transform 1 0 105216 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679581782
transform 1 0 105888 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679581782
transform 1 0 106560 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679581782
transform 1 0 107232 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679581782
transform 1 0 107904 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679581782
transform 1 0 108576 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679581782
transform 1 0 109248 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679581782
transform 1 0 109920 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679581782
transform 1 0 110592 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679581782
transform 1 0 111264 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679581782
transform 1 0 111936 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679581782
transform 1 0 112608 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679581782
transform 1 0 113280 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679581782
transform 1 0 113952 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679581782
transform 1 0 114624 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679581782
transform 1 0 115296 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679581782
transform 1 0 115968 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679581782
transform 1 0 116640 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679581782
transform 1 0 117312 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679581782
transform 1 0 117984 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679581782
transform 1 0 118656 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679581782
transform 1 0 119328 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679581782
transform 1 0 120000 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679581782
transform 1 0 120672 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679581782
transform 1 0 121344 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679581782
transform 1 0 122016 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679581782
transform 1 0 122688 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679581782
transform 1 0 123360 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679581782
transform 1 0 124032 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679581782
transform 1 0 124704 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679581782
transform 1 0 125376 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679581782
transform 1 0 126048 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679581782
transform 1 0 126720 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679581782
transform 1 0 127392 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679581782
transform 1 0 128064 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_595
timestamp 1679581782
transform 1 0 128736 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_602
timestamp 1679581782
transform 1 0 129408 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679581782
transform 1 0 130080 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_616
timestamp 1679581782
transform 1 0 130752 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_623
timestamp 1679581782
transform 1 0 131424 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_630
timestamp 1679581782
transform 1 0 132096 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_637
timestamp 1679581782
transform 1 0 132768 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_644
timestamp 1679581782
transform 1 0 133440 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_651
timestamp 1679581782
transform 1 0 134112 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_658
timestamp 1679581782
transform 1 0 134784 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_665
timestamp 1679581782
transform 1 0 135456 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_672
timestamp 1679581782
transform 1 0 136128 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_679
timestamp 1679581782
transform 1 0 136800 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_686
timestamp 1679581782
transform 1 0 137472 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_693
timestamp 1679581782
transform 1 0 138144 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_700
timestamp 1679581782
transform 1 0 138816 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_707
timestamp 1679581782
transform 1 0 139488 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_714
timestamp 1679581782
transform 1 0 140160 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_721
timestamp 1679581782
transform 1 0 140832 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_728
timestamp 1679581782
transform 1 0 141504 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_735
timestamp 1679581782
transform 1 0 142176 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_742
timestamp 1679581782
transform 1 0 142848 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_749
timestamp 1679581782
transform 1 0 143520 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_756
timestamp 1679581782
transform 1 0 144192 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_763
timestamp 1679581782
transform 1 0 144864 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_770
timestamp 1679581782
transform 1 0 145536 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_777
timestamp 1679581782
transform 1 0 146208 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_784
timestamp 1679581782
transform 1 0 146880 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_791
timestamp 1679581782
transform 1 0 147552 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_798
timestamp 1679581782
transform 1 0 148224 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_805
timestamp 1679581782
transform 1 0 148896 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_812
timestamp 1679581782
transform 1 0 149568 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_819
timestamp 1679581782
transform 1 0 150240 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_826
timestamp 1679581782
transform 1 0 150912 0 -1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_833
timestamp 1679581782
transform 1 0 151584 0 -1 73332
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_840
timestamp 1677579658
transform 1 0 152256 0 -1 73332
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679581782
transform 1 0 71616 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679581782
transform 1 0 72288 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679581782
transform 1 0 72960 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679581782
transform 1 0 73632 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679581782
transform 1 0 74304 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679581782
transform 1 0 74976 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679581782
transform 1 0 75648 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679581782
transform 1 0 76320 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679581782
transform 1 0 76992 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679581782
transform 1 0 77664 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679581782
transform 1 0 78336 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679581782
transform 1 0 79008 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679581782
transform 1 0 79680 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679581782
transform 1 0 80352 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679581782
transform 1 0 81024 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679581782
transform 1 0 81696 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679581782
transform 1 0 82368 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679581782
transform 1 0 83040 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679581782
transform 1 0 83712 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1679581782
transform 1 0 84384 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_140
timestamp 1679581782
transform 1 0 85056 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1679581782
transform 1 0 85728 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1679581782
transform 1 0 86400 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1679581782
transform 1 0 87072 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679581782
transform 1 0 87744 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1679581782
transform 1 0 88416 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1679581782
transform 1 0 89088 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_189
timestamp 1679581782
transform 1 0 89760 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_196
timestamp 1679581782
transform 1 0 90432 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_203
timestamp 1679581782
transform 1 0 91104 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_210
timestamp 1679581782
transform 1 0 91776 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_217
timestamp 1679581782
transform 1 0 92448 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_224
timestamp 1679581782
transform 1 0 93120 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_231
timestamp 1679581782
transform 1 0 93792 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_238
timestamp 1679581782
transform 1 0 94464 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_245
timestamp 1679581782
transform 1 0 95136 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_252
timestamp 1679581782
transform 1 0 95808 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_259
timestamp 1679581782
transform 1 0 96480 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_266
timestamp 1679581782
transform 1 0 97152 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_273
timestamp 1679581782
transform 1 0 97824 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_280
timestamp 1679581782
transform 1 0 98496 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_287
timestamp 1679581782
transform 1 0 99168 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_294
timestamp 1679581782
transform 1 0 99840 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_301
timestamp 1679581782
transform 1 0 100512 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_308
timestamp 1679581782
transform 1 0 101184 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_315
timestamp 1679581782
transform 1 0 101856 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_322
timestamp 1679581782
transform 1 0 102528 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_329
timestamp 1679581782
transform 1 0 103200 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_336
timestamp 1679581782
transform 1 0 103872 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_343
timestamp 1679581782
transform 1 0 104544 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_350
timestamp 1679581782
transform 1 0 105216 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_357
timestamp 1679581782
transform 1 0 105888 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_364
timestamp 1679581782
transform 1 0 106560 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_371
timestamp 1679581782
transform 1 0 107232 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_378
timestamp 1679581782
transform 1 0 107904 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_385
timestamp 1679581782
transform 1 0 108576 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_392
timestamp 1679581782
transform 1 0 109248 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_399
timestamp 1679581782
transform 1 0 109920 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_406
timestamp 1679581782
transform 1 0 110592 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_413
timestamp 1679581782
transform 1 0 111264 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_420
timestamp 1679581782
transform 1 0 111936 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_427
timestamp 1679581782
transform 1 0 112608 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_434
timestamp 1679581782
transform 1 0 113280 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_441
timestamp 1679581782
transform 1 0 113952 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_448
timestamp 1679581782
transform 1 0 114624 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_455
timestamp 1679581782
transform 1 0 115296 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_462
timestamp 1679581782
transform 1 0 115968 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_469
timestamp 1679581782
transform 1 0 116640 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_476
timestamp 1679581782
transform 1 0 117312 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_483
timestamp 1679581782
transform 1 0 117984 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_490
timestamp 1679581782
transform 1 0 118656 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_497
timestamp 1679581782
transform 1 0 119328 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_504
timestamp 1679581782
transform 1 0 120000 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_511
timestamp 1679581782
transform 1 0 120672 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_518
timestamp 1679581782
transform 1 0 121344 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_525
timestamp 1679581782
transform 1 0 122016 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_532
timestamp 1679581782
transform 1 0 122688 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_539
timestamp 1679581782
transform 1 0 123360 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_546
timestamp 1679581782
transform 1 0 124032 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_553
timestamp 1679581782
transform 1 0 124704 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_560
timestamp 1679581782
transform 1 0 125376 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_567
timestamp 1679581782
transform 1 0 126048 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_574
timestamp 1679581782
transform 1 0 126720 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_581
timestamp 1679581782
transform 1 0 127392 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_588
timestamp 1679581782
transform 1 0 128064 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_595
timestamp 1679581782
transform 1 0 128736 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_602
timestamp 1679581782
transform 1 0 129408 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_609
timestamp 1679581782
transform 1 0 130080 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_616
timestamp 1679581782
transform 1 0 130752 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_623
timestamp 1679581782
transform 1 0 131424 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_630
timestamp 1679581782
transform 1 0 132096 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_637
timestamp 1679581782
transform 1 0 132768 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_644
timestamp 1679581782
transform 1 0 133440 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_651
timestamp 1679581782
transform 1 0 134112 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_658
timestamp 1679581782
transform 1 0 134784 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_665
timestamp 1679581782
transform 1 0 135456 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_672
timestamp 1679581782
transform 1 0 136128 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_679
timestamp 1679581782
transform 1 0 136800 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_686
timestamp 1679581782
transform 1 0 137472 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_693
timestamp 1679581782
transform 1 0 138144 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_700
timestamp 1679581782
transform 1 0 138816 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_707
timestamp 1679581782
transform 1 0 139488 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_714
timestamp 1679581782
transform 1 0 140160 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_721
timestamp 1679581782
transform 1 0 140832 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_728
timestamp 1679581782
transform 1 0 141504 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_735
timestamp 1679581782
transform 1 0 142176 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_742
timestamp 1679581782
transform 1 0 142848 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_749
timestamp 1679581782
transform 1 0 143520 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_756
timestamp 1679581782
transform 1 0 144192 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_763
timestamp 1679581782
transform 1 0 144864 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_770
timestamp 1679581782
transform 1 0 145536 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_777
timestamp 1679581782
transform 1 0 146208 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_784
timestamp 1679581782
transform 1 0 146880 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_791
timestamp 1679581782
transform 1 0 147552 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_798
timestamp 1679581782
transform 1 0 148224 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_805
timestamp 1679581782
transform 1 0 148896 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_812
timestamp 1679581782
transform 1 0 149568 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_819
timestamp 1679581782
transform 1 0 150240 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_826
timestamp 1679581782
transform 1 0 150912 0 1 73332
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_833
timestamp 1679581782
transform 1 0 151584 0 1 73332
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_840
timestamp 1677579658
transform 1 0 152256 0 1 73332
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679581782
transform 1 0 71616 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679581782
transform 1 0 72288 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679581782
transform 1 0 72960 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679581782
transform 1 0 73632 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679581782
transform 1 0 74304 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679581782
transform 1 0 74976 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679581782
transform 1 0 75648 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679581782
transform 1 0 76320 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679581782
transform 1 0 76992 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679581782
transform 1 0 77664 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679581782
transform 1 0 78336 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679581782
transform 1 0 79008 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679581782
transform 1 0 79680 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1679581782
transform 1 0 80352 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1679581782
transform 1 0 81024 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1679581782
transform 1 0 81696 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1679581782
transform 1 0 82368 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1679581782
transform 1 0 83040 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_126
timestamp 1679581782
transform 1 0 83712 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1679581782
transform 1 0 84384 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_140
timestamp 1679581782
transform 1 0 85056 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1679581782
transform 1 0 85728 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1679581782
transform 1 0 86400 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1679581782
transform 1 0 87072 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_168
timestamp 1679581782
transform 1 0 87744 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_175
timestamp 1679581782
transform 1 0 88416 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_182
timestamp 1679581782
transform 1 0 89088 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_189
timestamp 1679581782
transform 1 0 89760 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_196
timestamp 1679581782
transform 1 0 90432 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_203
timestamp 1679581782
transform 1 0 91104 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_210
timestamp 1679581782
transform 1 0 91776 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_217
timestamp 1679581782
transform 1 0 92448 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_224
timestamp 1679581782
transform 1 0 93120 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_231
timestamp 1679581782
transform 1 0 93792 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_238
timestamp 1679581782
transform 1 0 94464 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1679581782
transform 1 0 95136 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_252
timestamp 1679581782
transform 1 0 95808 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_259
timestamp 1679581782
transform 1 0 96480 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_266
timestamp 1679581782
transform 1 0 97152 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_273
timestamp 1679581782
transform 1 0 97824 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_280
timestamp 1679581782
transform 1 0 98496 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_287
timestamp 1679581782
transform 1 0 99168 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_294
timestamp 1679581782
transform 1 0 99840 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_301
timestamp 1679581782
transform 1 0 100512 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_308
timestamp 1679581782
transform 1 0 101184 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_315
timestamp 1679581782
transform 1 0 101856 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_322
timestamp 1679581782
transform 1 0 102528 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_329
timestamp 1679581782
transform 1 0 103200 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_336
timestamp 1679581782
transform 1 0 103872 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_343
timestamp 1679581782
transform 1 0 104544 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_350
timestamp 1679581782
transform 1 0 105216 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_357
timestamp 1679581782
transform 1 0 105888 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_364
timestamp 1679581782
transform 1 0 106560 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_371
timestamp 1679581782
transform 1 0 107232 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_378
timestamp 1679581782
transform 1 0 107904 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_385
timestamp 1679581782
transform 1 0 108576 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_392
timestamp 1679581782
transform 1 0 109248 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_399
timestamp 1679581782
transform 1 0 109920 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_406
timestamp 1679581782
transform 1 0 110592 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_413
timestamp 1679581782
transform 1 0 111264 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_420
timestamp 1679581782
transform 1 0 111936 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_427
timestamp 1679581782
transform 1 0 112608 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_434
timestamp 1679581782
transform 1 0 113280 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_441
timestamp 1679581782
transform 1 0 113952 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_448
timestamp 1679581782
transform 1 0 114624 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_455
timestamp 1679581782
transform 1 0 115296 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_462
timestamp 1679581782
transform 1 0 115968 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_469
timestamp 1679581782
transform 1 0 116640 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_476
timestamp 1679581782
transform 1 0 117312 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_483
timestamp 1679581782
transform 1 0 117984 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_490
timestamp 1679581782
transform 1 0 118656 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_497
timestamp 1679581782
transform 1 0 119328 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_504
timestamp 1679581782
transform 1 0 120000 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_511
timestamp 1679581782
transform 1 0 120672 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_518
timestamp 1679581782
transform 1 0 121344 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_525
timestamp 1679581782
transform 1 0 122016 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_532
timestamp 1679581782
transform 1 0 122688 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_539
timestamp 1679581782
transform 1 0 123360 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_546
timestamp 1679581782
transform 1 0 124032 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_553
timestamp 1679581782
transform 1 0 124704 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_560
timestamp 1679581782
transform 1 0 125376 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_567
timestamp 1679581782
transform 1 0 126048 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_574
timestamp 1679581782
transform 1 0 126720 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_581
timestamp 1679581782
transform 1 0 127392 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_588
timestamp 1679581782
transform 1 0 128064 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_595
timestamp 1679581782
transform 1 0 128736 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_602
timestamp 1679581782
transform 1 0 129408 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_609
timestamp 1679581782
transform 1 0 130080 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_616
timestamp 1679581782
transform 1 0 130752 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_623
timestamp 1679581782
transform 1 0 131424 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_630
timestamp 1679581782
transform 1 0 132096 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_637
timestamp 1679581782
transform 1 0 132768 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_644
timestamp 1679581782
transform 1 0 133440 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_651
timestamp 1679581782
transform 1 0 134112 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_658
timestamp 1679581782
transform 1 0 134784 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_665
timestamp 1679581782
transform 1 0 135456 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_672
timestamp 1679581782
transform 1 0 136128 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_679
timestamp 1679581782
transform 1 0 136800 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_686
timestamp 1679581782
transform 1 0 137472 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_693
timestamp 1679581782
transform 1 0 138144 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_700
timestamp 1679581782
transform 1 0 138816 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_707
timestamp 1679581782
transform 1 0 139488 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_714
timestamp 1679581782
transform 1 0 140160 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_721
timestamp 1679581782
transform 1 0 140832 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_728
timestamp 1679581782
transform 1 0 141504 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_735
timestamp 1679581782
transform 1 0 142176 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_742
timestamp 1679581782
transform 1 0 142848 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_749
timestamp 1679581782
transform 1 0 143520 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_756
timestamp 1679581782
transform 1 0 144192 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_763
timestamp 1679581782
transform 1 0 144864 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_770
timestamp 1679581782
transform 1 0 145536 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_777
timestamp 1679581782
transform 1 0 146208 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_784
timestamp 1679581782
transform 1 0 146880 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_791
timestamp 1679581782
transform 1 0 147552 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_798
timestamp 1679581782
transform 1 0 148224 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_805
timestamp 1679581782
transform 1 0 148896 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_812
timestamp 1679581782
transform 1 0 149568 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_819
timestamp 1679581782
transform 1 0 150240 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_826
timestamp 1679581782
transform 1 0 150912 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_833
timestamp 1679581782
transform 1 0 151584 0 -1 74844
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_840
timestamp 1677579658
transform 1 0 152256 0 -1 74844
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679581782
transform 1 0 71616 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679581782
transform 1 0 72288 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679581782
transform 1 0 72960 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679581782
transform 1 0 73632 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679581782
transform 1 0 74304 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679581782
transform 1 0 74976 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679581782
transform 1 0 75648 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679581782
transform 1 0 76320 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679581782
transform 1 0 76992 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_63
timestamp 1679581782
transform 1 0 77664 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_70
timestamp 1679581782
transform 1 0 78336 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_77
timestamp 1679581782
transform 1 0 79008 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_84
timestamp 1679581782
transform 1 0 79680 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_91
timestamp 1679581782
transform 1 0 80352 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_98
timestamp 1679581782
transform 1 0 81024 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_105
timestamp 1679581782
transform 1 0 81696 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_112
timestamp 1679581782
transform 1 0 82368 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_119
timestamp 1679581782
transform 1 0 83040 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_126
timestamp 1679581782
transform 1 0 83712 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_133
timestamp 1679581782
transform 1 0 84384 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_140
timestamp 1679581782
transform 1 0 85056 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_147
timestamp 1679581782
transform 1 0 85728 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_154
timestamp 1679581782
transform 1 0 86400 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_161
timestamp 1679581782
transform 1 0 87072 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_168
timestamp 1679581782
transform 1 0 87744 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_175
timestamp 1679581782
transform 1 0 88416 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_182
timestamp 1679581782
transform 1 0 89088 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_189
timestamp 1679581782
transform 1 0 89760 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_196
timestamp 1679581782
transform 1 0 90432 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_203
timestamp 1679581782
transform 1 0 91104 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_210
timestamp 1679581782
transform 1 0 91776 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_217
timestamp 1679581782
transform 1 0 92448 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_224
timestamp 1679581782
transform 1 0 93120 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_231
timestamp 1679581782
transform 1 0 93792 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_238
timestamp 1679581782
transform 1 0 94464 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_245
timestamp 1679581782
transform 1 0 95136 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_252
timestamp 1679581782
transform 1 0 95808 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_259
timestamp 1679581782
transform 1 0 96480 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_266
timestamp 1679581782
transform 1 0 97152 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_273
timestamp 1679581782
transform 1 0 97824 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_280
timestamp 1679581782
transform 1 0 98496 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_287
timestamp 1679581782
transform 1 0 99168 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_294
timestamp 1679581782
transform 1 0 99840 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_301
timestamp 1679581782
transform 1 0 100512 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_308
timestamp 1679581782
transform 1 0 101184 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_315
timestamp 1679581782
transform 1 0 101856 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_322
timestamp 1679581782
transform 1 0 102528 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_329
timestamp 1679581782
transform 1 0 103200 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_336
timestamp 1679581782
transform 1 0 103872 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_343
timestamp 1679581782
transform 1 0 104544 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_350
timestamp 1679581782
transform 1 0 105216 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_357
timestamp 1679581782
transform 1 0 105888 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_364
timestamp 1679581782
transform 1 0 106560 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_371
timestamp 1679581782
transform 1 0 107232 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_378
timestamp 1679581782
transform 1 0 107904 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_385
timestamp 1679581782
transform 1 0 108576 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_392
timestamp 1679581782
transform 1 0 109248 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_399
timestamp 1679581782
transform 1 0 109920 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_406
timestamp 1679581782
transform 1 0 110592 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_413
timestamp 1679581782
transform 1 0 111264 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_420
timestamp 1679581782
transform 1 0 111936 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_427
timestamp 1679581782
transform 1 0 112608 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_434
timestamp 1679581782
transform 1 0 113280 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_441
timestamp 1679581782
transform 1 0 113952 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_448
timestamp 1679581782
transform 1 0 114624 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_455
timestamp 1679581782
transform 1 0 115296 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_462
timestamp 1679581782
transform 1 0 115968 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_469
timestamp 1679581782
transform 1 0 116640 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_476
timestamp 1679581782
transform 1 0 117312 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_483
timestamp 1679581782
transform 1 0 117984 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_490
timestamp 1679581782
transform 1 0 118656 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_497
timestamp 1679581782
transform 1 0 119328 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_504
timestamp 1679581782
transform 1 0 120000 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_511
timestamp 1679581782
transform 1 0 120672 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_518
timestamp 1679581782
transform 1 0 121344 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_525
timestamp 1679581782
transform 1 0 122016 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_532
timestamp 1679581782
transform 1 0 122688 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_539
timestamp 1679581782
transform 1 0 123360 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_546
timestamp 1679581782
transform 1 0 124032 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_553
timestamp 1679581782
transform 1 0 124704 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_560
timestamp 1679581782
transform 1 0 125376 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_567
timestamp 1679581782
transform 1 0 126048 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_574
timestamp 1679581782
transform 1 0 126720 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_581
timestamp 1679581782
transform 1 0 127392 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_588
timestamp 1679581782
transform 1 0 128064 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_595
timestamp 1679581782
transform 1 0 128736 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_602
timestamp 1679581782
transform 1 0 129408 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_609
timestamp 1679581782
transform 1 0 130080 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_616
timestamp 1679581782
transform 1 0 130752 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_623
timestamp 1679581782
transform 1 0 131424 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_630
timestamp 1679581782
transform 1 0 132096 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_637
timestamp 1679581782
transform 1 0 132768 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_644
timestamp 1679581782
transform 1 0 133440 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_651
timestamp 1679581782
transform 1 0 134112 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_658
timestamp 1679581782
transform 1 0 134784 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_665
timestamp 1679581782
transform 1 0 135456 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_672
timestamp 1679581782
transform 1 0 136128 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_679
timestamp 1679581782
transform 1 0 136800 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_686
timestamp 1679581782
transform 1 0 137472 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_693
timestamp 1679581782
transform 1 0 138144 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_700
timestamp 1679581782
transform 1 0 138816 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_707
timestamp 1679581782
transform 1 0 139488 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_714
timestamp 1679581782
transform 1 0 140160 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_721
timestamp 1679581782
transform 1 0 140832 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_728
timestamp 1679581782
transform 1 0 141504 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_735
timestamp 1679581782
transform 1 0 142176 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_742
timestamp 1679581782
transform 1 0 142848 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_749
timestamp 1679581782
transform 1 0 143520 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_756
timestamp 1679581782
transform 1 0 144192 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_763
timestamp 1679581782
transform 1 0 144864 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_770
timestamp 1679581782
transform 1 0 145536 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_777
timestamp 1679581782
transform 1 0 146208 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_784
timestamp 1679581782
transform 1 0 146880 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_791
timestamp 1679581782
transform 1 0 147552 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_798
timestamp 1679581782
transform 1 0 148224 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_805
timestamp 1679581782
transform 1 0 148896 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_812
timestamp 1679581782
transform 1 0 149568 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_819
timestamp 1679581782
transform 1 0 150240 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_826
timestamp 1679581782
transform 1 0 150912 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_833
timestamp 1679581782
transform 1 0 151584 0 1 74844
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_840
timestamp 1677579658
transform 1 0 152256 0 1 74844
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679581782
transform 1 0 71616 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679581782
transform 1 0 72288 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679581782
transform 1 0 72960 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679581782
transform 1 0 73632 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679581782
transform 1 0 74304 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679581782
transform 1 0 74976 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679581782
transform 1 0 75648 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1679581782
transform 1 0 76320 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_56
timestamp 1679581782
transform 1 0 76992 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_63
timestamp 1679581782
transform 1 0 77664 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679581782
transform 1 0 78336 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_77
timestamp 1679581782
transform 1 0 79008 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_84
timestamp 1679581782
transform 1 0 79680 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_91
timestamp 1679581782
transform 1 0 80352 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_98
timestamp 1679581782
transform 1 0 81024 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_105
timestamp 1679581782
transform 1 0 81696 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_112
timestamp 1679581782
transform 1 0 82368 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_119
timestamp 1679581782
transform 1 0 83040 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_126
timestamp 1679581782
transform 1 0 83712 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_133
timestamp 1679581782
transform 1 0 84384 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_140
timestamp 1679581782
transform 1 0 85056 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_147
timestamp 1679581782
transform 1 0 85728 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_154
timestamp 1679581782
transform 1 0 86400 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_161
timestamp 1679581782
transform 1 0 87072 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_168
timestamp 1679581782
transform 1 0 87744 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_175
timestamp 1679581782
transform 1 0 88416 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_182
timestamp 1679581782
transform 1 0 89088 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_189
timestamp 1679581782
transform 1 0 89760 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_196
timestamp 1679581782
transform 1 0 90432 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_203
timestamp 1679581782
transform 1 0 91104 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_210
timestamp 1679581782
transform 1 0 91776 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_217
timestamp 1679581782
transform 1 0 92448 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_224
timestamp 1679581782
transform 1 0 93120 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_231
timestamp 1679581782
transform 1 0 93792 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_238
timestamp 1679581782
transform 1 0 94464 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_245
timestamp 1679581782
transform 1 0 95136 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_252
timestamp 1679581782
transform 1 0 95808 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_259
timestamp 1679581782
transform 1 0 96480 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_266
timestamp 1679581782
transform 1 0 97152 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_273
timestamp 1679581782
transform 1 0 97824 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_280
timestamp 1679581782
transform 1 0 98496 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_287
timestamp 1679581782
transform 1 0 99168 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_294
timestamp 1679581782
transform 1 0 99840 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_301
timestamp 1679581782
transform 1 0 100512 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_308
timestamp 1679581782
transform 1 0 101184 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_315
timestamp 1679581782
transform 1 0 101856 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_322
timestamp 1679581782
transform 1 0 102528 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_329
timestamp 1679581782
transform 1 0 103200 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_336
timestamp 1679581782
transform 1 0 103872 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_343
timestamp 1679581782
transform 1 0 104544 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_350
timestamp 1679581782
transform 1 0 105216 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_357
timestamp 1679581782
transform 1 0 105888 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_364
timestamp 1679581782
transform 1 0 106560 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_371
timestamp 1679581782
transform 1 0 107232 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_378
timestamp 1679581782
transform 1 0 107904 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_385
timestamp 1679581782
transform 1 0 108576 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_392
timestamp 1679581782
transform 1 0 109248 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_399
timestamp 1679581782
transform 1 0 109920 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_406
timestamp 1679581782
transform 1 0 110592 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_413
timestamp 1679581782
transform 1 0 111264 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_420
timestamp 1679581782
transform 1 0 111936 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_427
timestamp 1679581782
transform 1 0 112608 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_434
timestamp 1679581782
transform 1 0 113280 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_441
timestamp 1679581782
transform 1 0 113952 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_448
timestamp 1679581782
transform 1 0 114624 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_455
timestamp 1679581782
transform 1 0 115296 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_462
timestamp 1679581782
transform 1 0 115968 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_469
timestamp 1679581782
transform 1 0 116640 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_476
timestamp 1679581782
transform 1 0 117312 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_483
timestamp 1679581782
transform 1 0 117984 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_490
timestamp 1679581782
transform 1 0 118656 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_497
timestamp 1679581782
transform 1 0 119328 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_504
timestamp 1679581782
transform 1 0 120000 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_511
timestamp 1679581782
transform 1 0 120672 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_518
timestamp 1679581782
transform 1 0 121344 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_525
timestamp 1679581782
transform 1 0 122016 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_532
timestamp 1679581782
transform 1 0 122688 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_539
timestamp 1679581782
transform 1 0 123360 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_546
timestamp 1679581782
transform 1 0 124032 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_553
timestamp 1679581782
transform 1 0 124704 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_560
timestamp 1679581782
transform 1 0 125376 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_567
timestamp 1679581782
transform 1 0 126048 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_574
timestamp 1679581782
transform 1 0 126720 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_581
timestamp 1679581782
transform 1 0 127392 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_588
timestamp 1679581782
transform 1 0 128064 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_595
timestamp 1679581782
transform 1 0 128736 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_602
timestamp 1679581782
transform 1 0 129408 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_609
timestamp 1679581782
transform 1 0 130080 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_616
timestamp 1679581782
transform 1 0 130752 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_623
timestamp 1679581782
transform 1 0 131424 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_630
timestamp 1679581782
transform 1 0 132096 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_637
timestamp 1679581782
transform 1 0 132768 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_644
timestamp 1679581782
transform 1 0 133440 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_651
timestamp 1679581782
transform 1 0 134112 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_658
timestamp 1679581782
transform 1 0 134784 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_665
timestamp 1679581782
transform 1 0 135456 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_672
timestamp 1679581782
transform 1 0 136128 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_679
timestamp 1679581782
transform 1 0 136800 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_686
timestamp 1679581782
transform 1 0 137472 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_693
timestamp 1679581782
transform 1 0 138144 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_700
timestamp 1679581782
transform 1 0 138816 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_707
timestamp 1679581782
transform 1 0 139488 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_714
timestamp 1679581782
transform 1 0 140160 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_721
timestamp 1679581782
transform 1 0 140832 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_728
timestamp 1679581782
transform 1 0 141504 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_735
timestamp 1679581782
transform 1 0 142176 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_742
timestamp 1679581782
transform 1 0 142848 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_749
timestamp 1679581782
transform 1 0 143520 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_756
timestamp 1679581782
transform 1 0 144192 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_763
timestamp 1679581782
transform 1 0 144864 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_770
timestamp 1679581782
transform 1 0 145536 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_777
timestamp 1679581782
transform 1 0 146208 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_784
timestamp 1679581782
transform 1 0 146880 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_791
timestamp 1679581782
transform 1 0 147552 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_798
timestamp 1679581782
transform 1 0 148224 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_805
timestamp 1679581782
transform 1 0 148896 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_812
timestamp 1679581782
transform 1 0 149568 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_819
timestamp 1679581782
transform 1 0 150240 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_826
timestamp 1679581782
transform 1 0 150912 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_833
timestamp 1679581782
transform 1 0 151584 0 -1 76356
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_840
timestamp 1677579658
transform 1 0 152256 0 -1 76356
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679581782
transform 1 0 71616 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679581782
transform 1 0 72288 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679581782
transform 1 0 72960 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679581782
transform 1 0 73632 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679581782
transform 1 0 74304 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679581782
transform 1 0 74976 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679581782
transform 1 0 75648 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679581782
transform 1 0 76320 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679581782
transform 1 0 76992 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679581782
transform 1 0 77664 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679581782
transform 1 0 78336 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679581782
transform 1 0 79008 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679581782
transform 1 0 79680 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_91
timestamp 1679581782
transform 1 0 80352 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679581782
transform 1 0 81024 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679581782
transform 1 0 81696 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_112
timestamp 1679581782
transform 1 0 82368 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_119
timestamp 1679581782
transform 1 0 83040 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_126
timestamp 1679581782
transform 1 0 83712 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_133
timestamp 1679581782
transform 1 0 84384 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_140
timestamp 1679581782
transform 1 0 85056 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_147
timestamp 1679581782
transform 1 0 85728 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_154
timestamp 1679581782
transform 1 0 86400 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_161
timestamp 1679581782
transform 1 0 87072 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_168
timestamp 1679581782
transform 1 0 87744 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_175
timestamp 1679581782
transform 1 0 88416 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_182
timestamp 1679581782
transform 1 0 89088 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_189
timestamp 1679581782
transform 1 0 89760 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_196
timestamp 1679581782
transform 1 0 90432 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_203
timestamp 1679581782
transform 1 0 91104 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_210
timestamp 1679581782
transform 1 0 91776 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_217
timestamp 1679581782
transform 1 0 92448 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_224
timestamp 1679581782
transform 1 0 93120 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_231
timestamp 1679581782
transform 1 0 93792 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_238
timestamp 1679581782
transform 1 0 94464 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_245
timestamp 1679581782
transform 1 0 95136 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_252
timestamp 1679581782
transform 1 0 95808 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_259
timestamp 1679581782
transform 1 0 96480 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_266
timestamp 1679581782
transform 1 0 97152 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_273
timestamp 1679581782
transform 1 0 97824 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_280
timestamp 1679581782
transform 1 0 98496 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_287
timestamp 1679581782
transform 1 0 99168 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_294
timestamp 1679581782
transform 1 0 99840 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_301
timestamp 1679581782
transform 1 0 100512 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_308
timestamp 1679581782
transform 1 0 101184 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_315
timestamp 1679581782
transform 1 0 101856 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_322
timestamp 1679581782
transform 1 0 102528 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_329
timestamp 1679581782
transform 1 0 103200 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_336
timestamp 1679581782
transform 1 0 103872 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_343
timestamp 1679581782
transform 1 0 104544 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_350
timestamp 1679581782
transform 1 0 105216 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_357
timestamp 1679581782
transform 1 0 105888 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_364
timestamp 1679581782
transform 1 0 106560 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_371
timestamp 1679581782
transform 1 0 107232 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_378
timestamp 1679581782
transform 1 0 107904 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_385
timestamp 1679581782
transform 1 0 108576 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_392
timestamp 1679581782
transform 1 0 109248 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_399
timestamp 1679581782
transform 1 0 109920 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_406
timestamp 1679581782
transform 1 0 110592 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_413
timestamp 1679581782
transform 1 0 111264 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_420
timestamp 1679581782
transform 1 0 111936 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_427
timestamp 1679581782
transform 1 0 112608 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_434
timestamp 1679581782
transform 1 0 113280 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_441
timestamp 1679581782
transform 1 0 113952 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_448
timestamp 1679581782
transform 1 0 114624 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_455
timestamp 1679581782
transform 1 0 115296 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_462
timestamp 1679581782
transform 1 0 115968 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_469
timestamp 1679581782
transform 1 0 116640 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_476
timestamp 1679581782
transform 1 0 117312 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_483
timestamp 1679581782
transform 1 0 117984 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_490
timestamp 1679581782
transform 1 0 118656 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_497
timestamp 1679581782
transform 1 0 119328 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_504
timestamp 1679581782
transform 1 0 120000 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_511
timestamp 1679581782
transform 1 0 120672 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_518
timestamp 1679581782
transform 1 0 121344 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_525
timestamp 1679581782
transform 1 0 122016 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_532
timestamp 1679581782
transform 1 0 122688 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_539
timestamp 1679581782
transform 1 0 123360 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_546
timestamp 1679581782
transform 1 0 124032 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_553
timestamp 1679581782
transform 1 0 124704 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_560
timestamp 1679581782
transform 1 0 125376 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_567
timestamp 1679581782
transform 1 0 126048 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_574
timestamp 1679581782
transform 1 0 126720 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_581
timestamp 1679581782
transform 1 0 127392 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_588
timestamp 1679581782
transform 1 0 128064 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_595
timestamp 1679581782
transform 1 0 128736 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_602
timestamp 1679581782
transform 1 0 129408 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_609
timestamp 1679581782
transform 1 0 130080 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_616
timestamp 1679581782
transform 1 0 130752 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_623
timestamp 1679581782
transform 1 0 131424 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_630
timestamp 1679581782
transform 1 0 132096 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_637
timestamp 1679581782
transform 1 0 132768 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_644
timestamp 1679581782
transform 1 0 133440 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_651
timestamp 1679581782
transform 1 0 134112 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_658
timestamp 1679581782
transform 1 0 134784 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_665
timestamp 1679581782
transform 1 0 135456 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_672
timestamp 1679581782
transform 1 0 136128 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_679
timestamp 1679581782
transform 1 0 136800 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_686
timestamp 1679581782
transform 1 0 137472 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_693
timestamp 1679581782
transform 1 0 138144 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_700
timestamp 1679581782
transform 1 0 138816 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_707
timestamp 1679581782
transform 1 0 139488 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_714
timestamp 1679581782
transform 1 0 140160 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_721
timestamp 1679581782
transform 1 0 140832 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_728
timestamp 1679581782
transform 1 0 141504 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_735
timestamp 1679581782
transform 1 0 142176 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_742
timestamp 1679581782
transform 1 0 142848 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_749
timestamp 1679581782
transform 1 0 143520 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_756
timestamp 1679581782
transform 1 0 144192 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_763
timestamp 1679581782
transform 1 0 144864 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_770
timestamp 1679581782
transform 1 0 145536 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_777
timestamp 1679581782
transform 1 0 146208 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_784
timestamp 1679581782
transform 1 0 146880 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_791
timestamp 1679581782
transform 1 0 147552 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_798
timestamp 1679581782
transform 1 0 148224 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_805
timestamp 1679581782
transform 1 0 148896 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_812
timestamp 1679581782
transform 1 0 149568 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_819
timestamp 1679581782
transform 1 0 150240 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_826
timestamp 1679581782
transform 1 0 150912 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_833
timestamp 1679581782
transform 1 0 151584 0 1 76356
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_840
timestamp 1677579658
transform 1 0 152256 0 1 76356
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679581782
transform 1 0 71616 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679581782
transform 1 0 72288 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679581782
transform 1 0 72960 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679581782
transform 1 0 73632 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679581782
transform 1 0 74304 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679581782
transform 1 0 74976 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679581782
transform 1 0 75648 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679581782
transform 1 0 76320 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679581782
transform 1 0 76992 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679581782
transform 1 0 77664 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679581782
transform 1 0 78336 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679581782
transform 1 0 79008 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679581782
transform 1 0 79680 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679581782
transform 1 0 80352 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_98
timestamp 1679581782
transform 1 0 81024 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679581782
transform 1 0 81696 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_112
timestamp 1679581782
transform 1 0 82368 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679581782
transform 1 0 83040 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_126
timestamp 1679581782
transform 1 0 83712 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679581782
transform 1 0 84384 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_140
timestamp 1679581782
transform 1 0 85056 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679581782
transform 1 0 85728 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_154
timestamp 1679581782
transform 1 0 86400 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679581782
transform 1 0 87072 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679581782
transform 1 0 87744 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_175
timestamp 1679581782
transform 1 0 88416 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_182
timestamp 1679581782
transform 1 0 89088 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_189
timestamp 1679581782
transform 1 0 89760 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_196
timestamp 1679581782
transform 1 0 90432 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_203
timestamp 1679581782
transform 1 0 91104 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_210
timestamp 1679581782
transform 1 0 91776 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_217
timestamp 1679581782
transform 1 0 92448 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_224
timestamp 1679581782
transform 1 0 93120 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_231
timestamp 1679581782
transform 1 0 93792 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_238
timestamp 1679581782
transform 1 0 94464 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_245
timestamp 1679581782
transform 1 0 95136 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_252
timestamp 1679581782
transform 1 0 95808 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_259
timestamp 1679581782
transform 1 0 96480 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_266
timestamp 1679581782
transform 1 0 97152 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_273
timestamp 1679581782
transform 1 0 97824 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_280
timestamp 1679581782
transform 1 0 98496 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_287
timestamp 1679581782
transform 1 0 99168 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_294
timestamp 1679581782
transform 1 0 99840 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_301
timestamp 1679581782
transform 1 0 100512 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_308
timestamp 1679581782
transform 1 0 101184 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_315
timestamp 1679581782
transform 1 0 101856 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_322
timestamp 1679581782
transform 1 0 102528 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_329
timestamp 1679581782
transform 1 0 103200 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_336
timestamp 1679581782
transform 1 0 103872 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_343
timestamp 1679581782
transform 1 0 104544 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_350
timestamp 1679581782
transform 1 0 105216 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_357
timestamp 1679581782
transform 1 0 105888 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_364
timestamp 1679581782
transform 1 0 106560 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_371
timestamp 1679581782
transform 1 0 107232 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_378
timestamp 1679581782
transform 1 0 107904 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_385
timestamp 1679581782
transform 1 0 108576 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_392
timestamp 1679581782
transform 1 0 109248 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_399
timestamp 1679581782
transform 1 0 109920 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_406
timestamp 1679581782
transform 1 0 110592 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_413
timestamp 1679581782
transform 1 0 111264 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_420
timestamp 1679581782
transform 1 0 111936 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_427
timestamp 1679581782
transform 1 0 112608 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_434
timestamp 1679581782
transform 1 0 113280 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_441
timestamp 1679581782
transform 1 0 113952 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_448
timestamp 1679581782
transform 1 0 114624 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_455
timestamp 1679581782
transform 1 0 115296 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_462
timestamp 1679581782
transform 1 0 115968 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_469
timestamp 1679581782
transform 1 0 116640 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_476
timestamp 1679581782
transform 1 0 117312 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_483
timestamp 1679581782
transform 1 0 117984 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_490
timestamp 1679581782
transform 1 0 118656 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_497
timestamp 1679581782
transform 1 0 119328 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_504
timestamp 1679581782
transform 1 0 120000 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_511
timestamp 1679581782
transform 1 0 120672 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_518
timestamp 1679581782
transform 1 0 121344 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_525
timestamp 1679581782
transform 1 0 122016 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_532
timestamp 1679581782
transform 1 0 122688 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_539
timestamp 1679581782
transform 1 0 123360 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_546
timestamp 1679581782
transform 1 0 124032 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_553
timestamp 1679581782
transform 1 0 124704 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_560
timestamp 1679581782
transform 1 0 125376 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_567
timestamp 1679581782
transform 1 0 126048 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_574
timestamp 1679581782
transform 1 0 126720 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_581
timestamp 1679581782
transform 1 0 127392 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_588
timestamp 1679581782
transform 1 0 128064 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_595
timestamp 1679581782
transform 1 0 128736 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_602
timestamp 1679581782
transform 1 0 129408 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_609
timestamp 1679581782
transform 1 0 130080 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_616
timestamp 1679581782
transform 1 0 130752 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_623
timestamp 1679581782
transform 1 0 131424 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_630
timestamp 1679581782
transform 1 0 132096 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_637
timestamp 1679581782
transform 1 0 132768 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_644
timestamp 1679581782
transform 1 0 133440 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_651
timestamp 1679581782
transform 1 0 134112 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_658
timestamp 1679581782
transform 1 0 134784 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_665
timestamp 1679581782
transform 1 0 135456 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_672
timestamp 1679581782
transform 1 0 136128 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_679
timestamp 1679581782
transform 1 0 136800 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_686
timestamp 1679581782
transform 1 0 137472 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_693
timestamp 1679581782
transform 1 0 138144 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_700
timestamp 1679581782
transform 1 0 138816 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_707
timestamp 1679581782
transform 1 0 139488 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_714
timestamp 1679581782
transform 1 0 140160 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_721
timestamp 1679581782
transform 1 0 140832 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_728
timestamp 1679581782
transform 1 0 141504 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_735
timestamp 1679581782
transform 1 0 142176 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_742
timestamp 1679581782
transform 1 0 142848 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_749
timestamp 1679581782
transform 1 0 143520 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_756
timestamp 1679581782
transform 1 0 144192 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_763
timestamp 1679581782
transform 1 0 144864 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_770
timestamp 1679581782
transform 1 0 145536 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_777
timestamp 1679581782
transform 1 0 146208 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_784
timestamp 1679581782
transform 1 0 146880 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_791
timestamp 1679581782
transform 1 0 147552 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_798
timestamp 1679581782
transform 1 0 148224 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_805
timestamp 1679581782
transform 1 0 148896 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_812
timestamp 1679581782
transform 1 0 149568 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_819
timestamp 1679581782
transform 1 0 150240 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_826
timestamp 1679581782
transform 1 0 150912 0 -1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_833
timestamp 1679581782
transform 1 0 151584 0 -1 77868
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_840
timestamp 1677579658
transform 1 0 152256 0 -1 77868
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679581782
transform 1 0 71616 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679581782
transform 1 0 72288 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679581782
transform 1 0 72960 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679581782
transform 1 0 73632 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679581782
transform 1 0 74304 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679581782
transform 1 0 74976 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679581782
transform 1 0 75648 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679581782
transform 1 0 76320 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679581782
transform 1 0 76992 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679581782
transform 1 0 77664 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679581782
transform 1 0 78336 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679581782
transform 1 0 79008 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679581782
transform 1 0 79680 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_91
timestamp 1679581782
transform 1 0 80352 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_98
timestamp 1679581782
transform 1 0 81024 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_105
timestamp 1679581782
transform 1 0 81696 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_112
timestamp 1679581782
transform 1 0 82368 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_119
timestamp 1679581782
transform 1 0 83040 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_126
timestamp 1679581782
transform 1 0 83712 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_133
timestamp 1679581782
transform 1 0 84384 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_140
timestamp 1679581782
transform 1 0 85056 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_147
timestamp 1679581782
transform 1 0 85728 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_154
timestamp 1679581782
transform 1 0 86400 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_161
timestamp 1679581782
transform 1 0 87072 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_168
timestamp 1679581782
transform 1 0 87744 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_175
timestamp 1679581782
transform 1 0 88416 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_182
timestamp 1679581782
transform 1 0 89088 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_189
timestamp 1679581782
transform 1 0 89760 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_196
timestamp 1679581782
transform 1 0 90432 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_203
timestamp 1679581782
transform 1 0 91104 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_210
timestamp 1679581782
transform 1 0 91776 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_217
timestamp 1679581782
transform 1 0 92448 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_224
timestamp 1679581782
transform 1 0 93120 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_231
timestamp 1679581782
transform 1 0 93792 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_238
timestamp 1679581782
transform 1 0 94464 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_245
timestamp 1679581782
transform 1 0 95136 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_252
timestamp 1679581782
transform 1 0 95808 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_259
timestamp 1679581782
transform 1 0 96480 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_266
timestamp 1679581782
transform 1 0 97152 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_273
timestamp 1679581782
transform 1 0 97824 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_280
timestamp 1679581782
transform 1 0 98496 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_287
timestamp 1679581782
transform 1 0 99168 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_294
timestamp 1679581782
transform 1 0 99840 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_301
timestamp 1679581782
transform 1 0 100512 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_308
timestamp 1679581782
transform 1 0 101184 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_315
timestamp 1679581782
transform 1 0 101856 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_322
timestamp 1679581782
transform 1 0 102528 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_329
timestamp 1679581782
transform 1 0 103200 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_336
timestamp 1679581782
transform 1 0 103872 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_343
timestamp 1679581782
transform 1 0 104544 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_350
timestamp 1679581782
transform 1 0 105216 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_357
timestamp 1679581782
transform 1 0 105888 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_364
timestamp 1679581782
transform 1 0 106560 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_371
timestamp 1679581782
transform 1 0 107232 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_378
timestamp 1679581782
transform 1 0 107904 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_385
timestamp 1679581782
transform 1 0 108576 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_392
timestamp 1679581782
transform 1 0 109248 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_399
timestamp 1679581782
transform 1 0 109920 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_406
timestamp 1679581782
transform 1 0 110592 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_413
timestamp 1679581782
transform 1 0 111264 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_420
timestamp 1679581782
transform 1 0 111936 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_427
timestamp 1679581782
transform 1 0 112608 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_434
timestamp 1679581782
transform 1 0 113280 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_441
timestamp 1679581782
transform 1 0 113952 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_448
timestamp 1679581782
transform 1 0 114624 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_455
timestamp 1679581782
transform 1 0 115296 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_462
timestamp 1679581782
transform 1 0 115968 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_469
timestamp 1679581782
transform 1 0 116640 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_476
timestamp 1679581782
transform 1 0 117312 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_483
timestamp 1679581782
transform 1 0 117984 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_490
timestamp 1679581782
transform 1 0 118656 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_497
timestamp 1679581782
transform 1 0 119328 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_504
timestamp 1679581782
transform 1 0 120000 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_511
timestamp 1679581782
transform 1 0 120672 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_518
timestamp 1679581782
transform 1 0 121344 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_525
timestamp 1679581782
transform 1 0 122016 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_532
timestamp 1679581782
transform 1 0 122688 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_539
timestamp 1679581782
transform 1 0 123360 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_546
timestamp 1679581782
transform 1 0 124032 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_553
timestamp 1679581782
transform 1 0 124704 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_560
timestamp 1679581782
transform 1 0 125376 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_567
timestamp 1679581782
transform 1 0 126048 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_574
timestamp 1679581782
transform 1 0 126720 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_581
timestamp 1679581782
transform 1 0 127392 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_588
timestamp 1679581782
transform 1 0 128064 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_595
timestamp 1679581782
transform 1 0 128736 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_602
timestamp 1679581782
transform 1 0 129408 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_609
timestamp 1679581782
transform 1 0 130080 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_616
timestamp 1679581782
transform 1 0 130752 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_623
timestamp 1679581782
transform 1 0 131424 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_630
timestamp 1679581782
transform 1 0 132096 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_637
timestamp 1679581782
transform 1 0 132768 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_644
timestamp 1679581782
transform 1 0 133440 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_651
timestamp 1679581782
transform 1 0 134112 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_658
timestamp 1679581782
transform 1 0 134784 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_665
timestamp 1679581782
transform 1 0 135456 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_672
timestamp 1679581782
transform 1 0 136128 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_679
timestamp 1679581782
transform 1 0 136800 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_686
timestamp 1679581782
transform 1 0 137472 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_693
timestamp 1679581782
transform 1 0 138144 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_700
timestamp 1679581782
transform 1 0 138816 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_707
timestamp 1679581782
transform 1 0 139488 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_714
timestamp 1679581782
transform 1 0 140160 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_721
timestamp 1679581782
transform 1 0 140832 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_728
timestamp 1679581782
transform 1 0 141504 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_735
timestamp 1679581782
transform 1 0 142176 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_742
timestamp 1679581782
transform 1 0 142848 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_749
timestamp 1679581782
transform 1 0 143520 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_756
timestamp 1679581782
transform 1 0 144192 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_763
timestamp 1679581782
transform 1 0 144864 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_770
timestamp 1679581782
transform 1 0 145536 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_777
timestamp 1679581782
transform 1 0 146208 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_784
timestamp 1679581782
transform 1 0 146880 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_791
timestamp 1679581782
transform 1 0 147552 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_798
timestamp 1679581782
transform 1 0 148224 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_805
timestamp 1679581782
transform 1 0 148896 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_812
timestamp 1679581782
transform 1 0 149568 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_819
timestamp 1679581782
transform 1 0 150240 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_826
timestamp 1679581782
transform 1 0 150912 0 1 77868
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_833
timestamp 1679581782
transform 1 0 151584 0 1 77868
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_840
timestamp 1677579658
transform 1 0 152256 0 1 77868
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 71616 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679581782
transform 1 0 72288 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679581782
transform 1 0 72960 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679581782
transform 1 0 73632 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679581782
transform 1 0 74304 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679581782
transform 1 0 74976 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679581782
transform 1 0 75648 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_49
timestamp 1679581782
transform 1 0 76320 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_56
timestamp 1679581782
transform 1 0 76992 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_63
timestamp 1679581782
transform 1 0 77664 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_70
timestamp 1679581782
transform 1 0 78336 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1679581782
transform 1 0 79008 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1679581782
transform 1 0 79680 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_91
timestamp 1679581782
transform 1 0 80352 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_98
timestamp 1679581782
transform 1 0 81024 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_105
timestamp 1679581782
transform 1 0 81696 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_112
timestamp 1679581782
transform 1 0 82368 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_119
timestamp 1679581782
transform 1 0 83040 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_126
timestamp 1679581782
transform 1 0 83712 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_133
timestamp 1679581782
transform 1 0 84384 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_140
timestamp 1679581782
transform 1 0 85056 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_147
timestamp 1679581782
transform 1 0 85728 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_154
timestamp 1679581782
transform 1 0 86400 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_161
timestamp 1679581782
transform 1 0 87072 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_168
timestamp 1679581782
transform 1 0 87744 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_175
timestamp 1679581782
transform 1 0 88416 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_182
timestamp 1679581782
transform 1 0 89088 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_189
timestamp 1679581782
transform 1 0 89760 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_196
timestamp 1679581782
transform 1 0 90432 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_203
timestamp 1679581782
transform 1 0 91104 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_210
timestamp 1679581782
transform 1 0 91776 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_217
timestamp 1679581782
transform 1 0 92448 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_224
timestamp 1679581782
transform 1 0 93120 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_231
timestamp 1679581782
transform 1 0 93792 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_238
timestamp 1679581782
transform 1 0 94464 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_245
timestamp 1679581782
transform 1 0 95136 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_252
timestamp 1679581782
transform 1 0 95808 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_259
timestamp 1679581782
transform 1 0 96480 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_266
timestamp 1679581782
transform 1 0 97152 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_273
timestamp 1679581782
transform 1 0 97824 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_280
timestamp 1679581782
transform 1 0 98496 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_287
timestamp 1679581782
transform 1 0 99168 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_294
timestamp 1679581782
transform 1 0 99840 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_301
timestamp 1679581782
transform 1 0 100512 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_308
timestamp 1679581782
transform 1 0 101184 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_315
timestamp 1679581782
transform 1 0 101856 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_322
timestamp 1679581782
transform 1 0 102528 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_329
timestamp 1679581782
transform 1 0 103200 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_336
timestamp 1679581782
transform 1 0 103872 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_343
timestamp 1679581782
transform 1 0 104544 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_350
timestamp 1679581782
transform 1 0 105216 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_357
timestamp 1679581782
transform 1 0 105888 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_364
timestamp 1679581782
transform 1 0 106560 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_371
timestamp 1679581782
transform 1 0 107232 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_378
timestamp 1679581782
transform 1 0 107904 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_385
timestamp 1679581782
transform 1 0 108576 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_392
timestamp 1679581782
transform 1 0 109248 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_399
timestamp 1679581782
transform 1 0 109920 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_406
timestamp 1679581782
transform 1 0 110592 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_413
timestamp 1679581782
transform 1 0 111264 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_420
timestamp 1679581782
transform 1 0 111936 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_427
timestamp 1679581782
transform 1 0 112608 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_434
timestamp 1679581782
transform 1 0 113280 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_441
timestamp 1679581782
transform 1 0 113952 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_448
timestamp 1679581782
transform 1 0 114624 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_455
timestamp 1679581782
transform 1 0 115296 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_462
timestamp 1679581782
transform 1 0 115968 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_469
timestamp 1679581782
transform 1 0 116640 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_476
timestamp 1679581782
transform 1 0 117312 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_483
timestamp 1679581782
transform 1 0 117984 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_490
timestamp 1679581782
transform 1 0 118656 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_497
timestamp 1679581782
transform 1 0 119328 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_504
timestamp 1679581782
transform 1 0 120000 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_511
timestamp 1679581782
transform 1 0 120672 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_518
timestamp 1679581782
transform 1 0 121344 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_525
timestamp 1679581782
transform 1 0 122016 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_532
timestamp 1679581782
transform 1 0 122688 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_539
timestamp 1679581782
transform 1 0 123360 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_546
timestamp 1679581782
transform 1 0 124032 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_553
timestamp 1679581782
transform 1 0 124704 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_560
timestamp 1679581782
transform 1 0 125376 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_567
timestamp 1679581782
transform 1 0 126048 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_574
timestamp 1679581782
transform 1 0 126720 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_581
timestamp 1679581782
transform 1 0 127392 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_588
timestamp 1679581782
transform 1 0 128064 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_595
timestamp 1679581782
transform 1 0 128736 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_602
timestamp 1679581782
transform 1 0 129408 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_609
timestamp 1679581782
transform 1 0 130080 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_616
timestamp 1679581782
transform 1 0 130752 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_623
timestamp 1679581782
transform 1 0 131424 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_630
timestamp 1679581782
transform 1 0 132096 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_637
timestamp 1679581782
transform 1 0 132768 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_644
timestamp 1679581782
transform 1 0 133440 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_651
timestamp 1679581782
transform 1 0 134112 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_658
timestamp 1679581782
transform 1 0 134784 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_665
timestamp 1679581782
transform 1 0 135456 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_672
timestamp 1679581782
transform 1 0 136128 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_679
timestamp 1679581782
transform 1 0 136800 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_686
timestamp 1679581782
transform 1 0 137472 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_693
timestamp 1679581782
transform 1 0 138144 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_700
timestamp 1679581782
transform 1 0 138816 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_707
timestamp 1679581782
transform 1 0 139488 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_714
timestamp 1679581782
transform 1 0 140160 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_721
timestamp 1679581782
transform 1 0 140832 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_728
timestamp 1679581782
transform 1 0 141504 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_735
timestamp 1679581782
transform 1 0 142176 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_742
timestamp 1679581782
transform 1 0 142848 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_749
timestamp 1679581782
transform 1 0 143520 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_756
timestamp 1679581782
transform 1 0 144192 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_763
timestamp 1679581782
transform 1 0 144864 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_770
timestamp 1679581782
transform 1 0 145536 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_777
timestamp 1679581782
transform 1 0 146208 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_784
timestamp 1679581782
transform 1 0 146880 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_791
timestamp 1679581782
transform 1 0 147552 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_798
timestamp 1679581782
transform 1 0 148224 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_805
timestamp 1679581782
transform 1 0 148896 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_812
timestamp 1679581782
transform 1 0 149568 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_819
timestamp 1679581782
transform 1 0 150240 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_826
timestamp 1679581782
transform 1 0 150912 0 -1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_833
timestamp 1679581782
transform 1 0 151584 0 -1 79380
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_840
timestamp 1677579658
transform 1 0 152256 0 -1 79380
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679581782
transform 1 0 71616 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679581782
transform 1 0 72288 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1679581782
transform 1 0 72960 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_21
timestamp 1679581782
transform 1 0 73632 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_28
timestamp 1679581782
transform 1 0 74304 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_35
timestamp 1679581782
transform 1 0 74976 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_42
timestamp 1679581782
transform 1 0 75648 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_49
timestamp 1679581782
transform 1 0 76320 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_56
timestamp 1679581782
transform 1 0 76992 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_63
timestamp 1679581782
transform 1 0 77664 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_70
timestamp 1679581782
transform 1 0 78336 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_77
timestamp 1679581782
transform 1 0 79008 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_84
timestamp 1679581782
transform 1 0 79680 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_91
timestamp 1679581782
transform 1 0 80352 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_98
timestamp 1679581782
transform 1 0 81024 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_105
timestamp 1679581782
transform 1 0 81696 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_112
timestamp 1679581782
transform 1 0 82368 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_119
timestamp 1679581782
transform 1 0 83040 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_126
timestamp 1679581782
transform 1 0 83712 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_133
timestamp 1679581782
transform 1 0 84384 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_140
timestamp 1679581782
transform 1 0 85056 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_147
timestamp 1679581782
transform 1 0 85728 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_154
timestamp 1679581782
transform 1 0 86400 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_161
timestamp 1679581782
transform 1 0 87072 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_168
timestamp 1679581782
transform 1 0 87744 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_175
timestamp 1679581782
transform 1 0 88416 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_182
timestamp 1679581782
transform 1 0 89088 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_189
timestamp 1679581782
transform 1 0 89760 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_196
timestamp 1679581782
transform 1 0 90432 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_203
timestamp 1679581782
transform 1 0 91104 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_210
timestamp 1679581782
transform 1 0 91776 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_217
timestamp 1679581782
transform 1 0 92448 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_224
timestamp 1679581782
transform 1 0 93120 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_231
timestamp 1679581782
transform 1 0 93792 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_238
timestamp 1679581782
transform 1 0 94464 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_245
timestamp 1679581782
transform 1 0 95136 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_252
timestamp 1679581782
transform 1 0 95808 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_259
timestamp 1679581782
transform 1 0 96480 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_266
timestamp 1679581782
transform 1 0 97152 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_273
timestamp 1679581782
transform 1 0 97824 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_280
timestamp 1679581782
transform 1 0 98496 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_287
timestamp 1679581782
transform 1 0 99168 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_294
timestamp 1679581782
transform 1 0 99840 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_301
timestamp 1679581782
transform 1 0 100512 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_308
timestamp 1679581782
transform 1 0 101184 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_315
timestamp 1679581782
transform 1 0 101856 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_322
timestamp 1679581782
transform 1 0 102528 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_329
timestamp 1679581782
transform 1 0 103200 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_336
timestamp 1679581782
transform 1 0 103872 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_343
timestamp 1679581782
transform 1 0 104544 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_350
timestamp 1679581782
transform 1 0 105216 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_357
timestamp 1679581782
transform 1 0 105888 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_364
timestamp 1679581782
transform 1 0 106560 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_371
timestamp 1679581782
transform 1 0 107232 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_378
timestamp 1679581782
transform 1 0 107904 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_385
timestamp 1679581782
transform 1 0 108576 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_392
timestamp 1679581782
transform 1 0 109248 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_399
timestamp 1679581782
transform 1 0 109920 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_406
timestamp 1679581782
transform 1 0 110592 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_413
timestamp 1679581782
transform 1 0 111264 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_420
timestamp 1679581782
transform 1 0 111936 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_427
timestamp 1679581782
transform 1 0 112608 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_434
timestamp 1679581782
transform 1 0 113280 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_441
timestamp 1679581782
transform 1 0 113952 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_448
timestamp 1679581782
transform 1 0 114624 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_455
timestamp 1679581782
transform 1 0 115296 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_462
timestamp 1679581782
transform 1 0 115968 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_469
timestamp 1679581782
transform 1 0 116640 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_476
timestamp 1679581782
transform 1 0 117312 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_483
timestamp 1679581782
transform 1 0 117984 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_490
timestamp 1679581782
transform 1 0 118656 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_497
timestamp 1679581782
transform 1 0 119328 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_504
timestamp 1679581782
transform 1 0 120000 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_511
timestamp 1679581782
transform 1 0 120672 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_518
timestamp 1679581782
transform 1 0 121344 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_525
timestamp 1679581782
transform 1 0 122016 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_532
timestamp 1679581782
transform 1 0 122688 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_539
timestamp 1679581782
transform 1 0 123360 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_546
timestamp 1679581782
transform 1 0 124032 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_553
timestamp 1679581782
transform 1 0 124704 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_560
timestamp 1679581782
transform 1 0 125376 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_567
timestamp 1679581782
transform 1 0 126048 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_574
timestamp 1679581782
transform 1 0 126720 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_581
timestamp 1679581782
transform 1 0 127392 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_588
timestamp 1679581782
transform 1 0 128064 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_595
timestamp 1679581782
transform 1 0 128736 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_602
timestamp 1679581782
transform 1 0 129408 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_609
timestamp 1679581782
transform 1 0 130080 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_616
timestamp 1679581782
transform 1 0 130752 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_623
timestamp 1679581782
transform 1 0 131424 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_630
timestamp 1679581782
transform 1 0 132096 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_637
timestamp 1679581782
transform 1 0 132768 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_644
timestamp 1679581782
transform 1 0 133440 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_651
timestamp 1679581782
transform 1 0 134112 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_658
timestamp 1679581782
transform 1 0 134784 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_665
timestamp 1679581782
transform 1 0 135456 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_672
timestamp 1679581782
transform 1 0 136128 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_679
timestamp 1679581782
transform 1 0 136800 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_686
timestamp 1679581782
transform 1 0 137472 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_693
timestamp 1679581782
transform 1 0 138144 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_700
timestamp 1679581782
transform 1 0 138816 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_707
timestamp 1679581782
transform 1 0 139488 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_714
timestamp 1679581782
transform 1 0 140160 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_721
timestamp 1679581782
transform 1 0 140832 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_728
timestamp 1679581782
transform 1 0 141504 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_735
timestamp 1679581782
transform 1 0 142176 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_742
timestamp 1679581782
transform 1 0 142848 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_749
timestamp 1679581782
transform 1 0 143520 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_756
timestamp 1679581782
transform 1 0 144192 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_763
timestamp 1679581782
transform 1 0 144864 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_770
timestamp 1679581782
transform 1 0 145536 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_777
timestamp 1679581782
transform 1 0 146208 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_784
timestamp 1679581782
transform 1 0 146880 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_791
timestamp 1679581782
transform 1 0 147552 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_798
timestamp 1679581782
transform 1 0 148224 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_805
timestamp 1679581782
transform 1 0 148896 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_812
timestamp 1679581782
transform 1 0 149568 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_819
timestamp 1679581782
transform 1 0 150240 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_826
timestamp 1679581782
transform 1 0 150912 0 1 79380
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_833
timestamp 1679581782
transform 1 0 151584 0 1 79380
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_840
timestamp 1677579658
transform 1 0 152256 0 1 79380
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1679581782
transform 1 0 71616 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_7
timestamp 1679581782
transform 1 0 72288 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_14
timestamp 1679581782
transform 1 0 72960 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_21
timestamp 1679581782
transform 1 0 73632 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_28
timestamp 1679581782
transform 1 0 74304 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_35
timestamp 1679581782
transform 1 0 74976 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_42
timestamp 1679581782
transform 1 0 75648 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_49
timestamp 1679581782
transform 1 0 76320 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_56
timestamp 1679581782
transform 1 0 76992 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_63
timestamp 1679581782
transform 1 0 77664 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_70
timestamp 1679581782
transform 1 0 78336 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_77
timestamp 1679581782
transform 1 0 79008 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_84
timestamp 1679581782
transform 1 0 79680 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_91
timestamp 1679581782
transform 1 0 80352 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_98
timestamp 1679581782
transform 1 0 81024 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_105
timestamp 1679581782
transform 1 0 81696 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_112
timestamp 1679581782
transform 1 0 82368 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_119
timestamp 1679581782
transform 1 0 83040 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_126
timestamp 1679581782
transform 1 0 83712 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_133
timestamp 1679581782
transform 1 0 84384 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_140
timestamp 1679581782
transform 1 0 85056 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_147
timestamp 1679581782
transform 1 0 85728 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_154
timestamp 1679581782
transform 1 0 86400 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_161
timestamp 1679581782
transform 1 0 87072 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_168
timestamp 1679581782
transform 1 0 87744 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_175
timestamp 1679581782
transform 1 0 88416 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_182
timestamp 1679581782
transform 1 0 89088 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_189
timestamp 1679581782
transform 1 0 89760 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_196
timestamp 1679581782
transform 1 0 90432 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_203
timestamp 1679581782
transform 1 0 91104 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_210
timestamp 1679581782
transform 1 0 91776 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_217
timestamp 1679581782
transform 1 0 92448 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_224
timestamp 1679581782
transform 1 0 93120 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_231
timestamp 1679581782
transform 1 0 93792 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_238
timestamp 1679581782
transform 1 0 94464 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_245
timestamp 1679581782
transform 1 0 95136 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_252
timestamp 1679581782
transform 1 0 95808 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_259
timestamp 1679581782
transform 1 0 96480 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_266
timestamp 1679581782
transform 1 0 97152 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_273
timestamp 1679581782
transform 1 0 97824 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_280
timestamp 1679581782
transform 1 0 98496 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_287
timestamp 1679581782
transform 1 0 99168 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_294
timestamp 1679581782
transform 1 0 99840 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_301
timestamp 1679581782
transform 1 0 100512 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_308
timestamp 1679581782
transform 1 0 101184 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_315
timestamp 1679581782
transform 1 0 101856 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_322
timestamp 1679581782
transform 1 0 102528 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_329
timestamp 1679581782
transform 1 0 103200 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_336
timestamp 1679581782
transform 1 0 103872 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_343
timestamp 1679581782
transform 1 0 104544 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_350
timestamp 1679581782
transform 1 0 105216 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_357
timestamp 1679581782
transform 1 0 105888 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_364
timestamp 1679581782
transform 1 0 106560 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_371
timestamp 1679581782
transform 1 0 107232 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_378
timestamp 1679581782
transform 1 0 107904 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_385
timestamp 1679581782
transform 1 0 108576 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_392
timestamp 1679581782
transform 1 0 109248 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_399
timestamp 1679581782
transform 1 0 109920 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_406
timestamp 1679581782
transform 1 0 110592 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_413
timestamp 1679581782
transform 1 0 111264 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_420
timestamp 1679581782
transform 1 0 111936 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_427
timestamp 1679581782
transform 1 0 112608 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_434
timestamp 1679581782
transform 1 0 113280 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_441
timestamp 1679581782
transform 1 0 113952 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_448
timestamp 1679581782
transform 1 0 114624 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_455
timestamp 1679581782
transform 1 0 115296 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_462
timestamp 1679581782
transform 1 0 115968 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_469
timestamp 1679581782
transform 1 0 116640 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_476
timestamp 1679581782
transform 1 0 117312 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_483
timestamp 1679581782
transform 1 0 117984 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_490
timestamp 1679581782
transform 1 0 118656 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_497
timestamp 1679581782
transform 1 0 119328 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_504
timestamp 1679581782
transform 1 0 120000 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_511
timestamp 1679581782
transform 1 0 120672 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_518
timestamp 1679581782
transform 1 0 121344 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_525
timestamp 1679581782
transform 1 0 122016 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_532
timestamp 1679581782
transform 1 0 122688 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_539
timestamp 1679581782
transform 1 0 123360 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_546
timestamp 1679581782
transform 1 0 124032 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_553
timestamp 1679581782
transform 1 0 124704 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_560
timestamp 1679581782
transform 1 0 125376 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_567
timestamp 1679581782
transform 1 0 126048 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_574
timestamp 1679581782
transform 1 0 126720 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_581
timestamp 1679581782
transform 1 0 127392 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_588
timestamp 1679581782
transform 1 0 128064 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_595
timestamp 1679581782
transform 1 0 128736 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_602
timestamp 1679581782
transform 1 0 129408 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_609
timestamp 1679581782
transform 1 0 130080 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_616
timestamp 1679581782
transform 1 0 130752 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_623
timestamp 1679581782
transform 1 0 131424 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_630
timestamp 1679581782
transform 1 0 132096 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_637
timestamp 1679581782
transform 1 0 132768 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_644
timestamp 1679581782
transform 1 0 133440 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_651
timestamp 1679581782
transform 1 0 134112 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_658
timestamp 1679581782
transform 1 0 134784 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_665
timestamp 1679581782
transform 1 0 135456 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_672
timestamp 1679581782
transform 1 0 136128 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_679
timestamp 1679581782
transform 1 0 136800 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_686
timestamp 1679581782
transform 1 0 137472 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_693
timestamp 1679581782
transform 1 0 138144 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_700
timestamp 1679581782
transform 1 0 138816 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_707
timestamp 1679581782
transform 1 0 139488 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_714
timestamp 1679581782
transform 1 0 140160 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_721
timestamp 1679581782
transform 1 0 140832 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_728
timestamp 1679581782
transform 1 0 141504 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_735
timestamp 1679581782
transform 1 0 142176 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_742
timestamp 1679581782
transform 1 0 142848 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_749
timestamp 1679581782
transform 1 0 143520 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_756
timestamp 1679581782
transform 1 0 144192 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_763
timestamp 1679581782
transform 1 0 144864 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_770
timestamp 1679581782
transform 1 0 145536 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_777
timestamp 1679581782
transform 1 0 146208 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_784
timestamp 1679581782
transform 1 0 146880 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_791
timestamp 1679581782
transform 1 0 147552 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_798
timestamp 1679581782
transform 1 0 148224 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_805
timestamp 1679581782
transform 1 0 148896 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_812
timestamp 1679581782
transform 1 0 149568 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_819
timestamp 1679581782
transform 1 0 150240 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_826
timestamp 1679581782
transform 1 0 150912 0 -1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_833
timestamp 1679581782
transform 1 0 151584 0 -1 80892
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_840
timestamp 1677579658
transform 1 0 152256 0 -1 80892
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_0
timestamp 1679581782
transform 1 0 71616 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_7
timestamp 1679581782
transform 1 0 72288 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_14
timestamp 1679581782
transform 1 0 72960 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_21
timestamp 1679581782
transform 1 0 73632 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_28
timestamp 1679581782
transform 1 0 74304 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_35
timestamp 1679581782
transform 1 0 74976 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_42
timestamp 1679581782
transform 1 0 75648 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_49
timestamp 1679581782
transform 1 0 76320 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_56
timestamp 1679581782
transform 1 0 76992 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_63
timestamp 1679581782
transform 1 0 77664 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_70
timestamp 1679581782
transform 1 0 78336 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_77
timestamp 1679581782
transform 1 0 79008 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_84
timestamp 1679581782
transform 1 0 79680 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_91
timestamp 1679581782
transform 1 0 80352 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_98
timestamp 1679581782
transform 1 0 81024 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_105
timestamp 1679581782
transform 1 0 81696 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_112
timestamp 1679581782
transform 1 0 82368 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_119
timestamp 1679581782
transform 1 0 83040 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_126
timestamp 1679581782
transform 1 0 83712 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_133
timestamp 1679581782
transform 1 0 84384 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_140
timestamp 1679581782
transform 1 0 85056 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_147
timestamp 1679581782
transform 1 0 85728 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_154
timestamp 1679581782
transform 1 0 86400 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_161
timestamp 1679581782
transform 1 0 87072 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_168
timestamp 1679581782
transform 1 0 87744 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_175
timestamp 1679581782
transform 1 0 88416 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_182
timestamp 1679581782
transform 1 0 89088 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_189
timestamp 1679581782
transform 1 0 89760 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_196
timestamp 1679581782
transform 1 0 90432 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_203
timestamp 1679581782
transform 1 0 91104 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_210
timestamp 1679581782
transform 1 0 91776 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_217
timestamp 1679581782
transform 1 0 92448 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_224
timestamp 1679581782
transform 1 0 93120 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_231
timestamp 1679581782
transform 1 0 93792 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_238
timestamp 1679581782
transform 1 0 94464 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_245
timestamp 1679581782
transform 1 0 95136 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_252
timestamp 1679581782
transform 1 0 95808 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_259
timestamp 1679581782
transform 1 0 96480 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_266
timestamp 1679581782
transform 1 0 97152 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_273
timestamp 1679581782
transform 1 0 97824 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_280
timestamp 1679581782
transform 1 0 98496 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_287
timestamp 1679581782
transform 1 0 99168 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_294
timestamp 1679581782
transform 1 0 99840 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_301
timestamp 1679581782
transform 1 0 100512 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_308
timestamp 1679581782
transform 1 0 101184 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_315
timestamp 1679581782
transform 1 0 101856 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_322
timestamp 1679581782
transform 1 0 102528 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_329
timestamp 1679581782
transform 1 0 103200 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_336
timestamp 1679581782
transform 1 0 103872 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_343
timestamp 1679581782
transform 1 0 104544 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_350
timestamp 1679581782
transform 1 0 105216 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_357
timestamp 1679581782
transform 1 0 105888 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_364
timestamp 1679581782
transform 1 0 106560 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_371
timestamp 1679581782
transform 1 0 107232 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_378
timestamp 1679581782
transform 1 0 107904 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_385
timestamp 1679581782
transform 1 0 108576 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_392
timestamp 1679581782
transform 1 0 109248 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_399
timestamp 1679581782
transform 1 0 109920 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_406
timestamp 1679581782
transform 1 0 110592 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_413
timestamp 1679581782
transform 1 0 111264 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_420
timestamp 1679581782
transform 1 0 111936 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_427
timestamp 1679581782
transform 1 0 112608 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_434
timestamp 1679581782
transform 1 0 113280 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_441
timestamp 1679581782
transform 1 0 113952 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_448
timestamp 1679581782
transform 1 0 114624 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_455
timestamp 1679581782
transform 1 0 115296 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_462
timestamp 1679581782
transform 1 0 115968 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_469
timestamp 1679581782
transform 1 0 116640 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_476
timestamp 1679581782
transform 1 0 117312 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_483
timestamp 1679581782
transform 1 0 117984 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_490
timestamp 1679581782
transform 1 0 118656 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_497
timestamp 1679581782
transform 1 0 119328 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_504
timestamp 1679581782
transform 1 0 120000 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_511
timestamp 1679581782
transform 1 0 120672 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_518
timestamp 1679581782
transform 1 0 121344 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_525
timestamp 1679581782
transform 1 0 122016 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_532
timestamp 1679581782
transform 1 0 122688 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_539
timestamp 1679581782
transform 1 0 123360 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_546
timestamp 1679581782
transform 1 0 124032 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_553
timestamp 1679581782
transform 1 0 124704 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_560
timestamp 1679581782
transform 1 0 125376 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_567
timestamp 1679581782
transform 1 0 126048 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_574
timestamp 1679581782
transform 1 0 126720 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_581
timestamp 1679581782
transform 1 0 127392 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_588
timestamp 1679581782
transform 1 0 128064 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_595
timestamp 1679581782
transform 1 0 128736 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_602
timestamp 1679581782
transform 1 0 129408 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_609
timestamp 1679581782
transform 1 0 130080 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_616
timestamp 1679581782
transform 1 0 130752 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_623
timestamp 1679581782
transform 1 0 131424 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_630
timestamp 1679581782
transform 1 0 132096 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_637
timestamp 1679581782
transform 1 0 132768 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_644
timestamp 1679581782
transform 1 0 133440 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_651
timestamp 1679581782
transform 1 0 134112 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_658
timestamp 1679581782
transform 1 0 134784 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_665
timestamp 1679581782
transform 1 0 135456 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_672
timestamp 1679581782
transform 1 0 136128 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_679
timestamp 1679581782
transform 1 0 136800 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_686
timestamp 1679581782
transform 1 0 137472 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_693
timestamp 1679581782
transform 1 0 138144 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_700
timestamp 1679581782
transform 1 0 138816 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_707
timestamp 1679581782
transform 1 0 139488 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_714
timestamp 1679581782
transform 1 0 140160 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_721
timestamp 1679581782
transform 1 0 140832 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_728
timestamp 1679581782
transform 1 0 141504 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_735
timestamp 1679581782
transform 1 0 142176 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_742
timestamp 1679581782
transform 1 0 142848 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_749
timestamp 1679581782
transform 1 0 143520 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_756
timestamp 1679581782
transform 1 0 144192 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_763
timestamp 1679581782
transform 1 0 144864 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_770
timestamp 1679581782
transform 1 0 145536 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_777
timestamp 1679581782
transform 1 0 146208 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_784
timestamp 1679581782
transform 1 0 146880 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_791
timestamp 1679581782
transform 1 0 147552 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_798
timestamp 1679581782
transform 1 0 148224 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_805
timestamp 1679581782
transform 1 0 148896 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_812
timestamp 1679581782
transform 1 0 149568 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_819
timestamp 1679581782
transform 1 0 150240 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_826
timestamp 1679581782
transform 1 0 150912 0 1 80892
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_833
timestamp 1679581782
transform 1 0 151584 0 1 80892
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_840
timestamp 1677579658
transform 1 0 152256 0 1 80892
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_0
timestamp 1679581782
transform 1 0 71616 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_7
timestamp 1679581782
transform 1 0 72288 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_14
timestamp 1679581782
transform 1 0 72960 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_21
timestamp 1679581782
transform 1 0 73632 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_28
timestamp 1679581782
transform 1 0 74304 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_35
timestamp 1679581782
transform 1 0 74976 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_42
timestamp 1679581782
transform 1 0 75648 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_49
timestamp 1679581782
transform 1 0 76320 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_56
timestamp 1679581782
transform 1 0 76992 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_63
timestamp 1679581782
transform 1 0 77664 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_70
timestamp 1679581782
transform 1 0 78336 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_77
timestamp 1679581782
transform 1 0 79008 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_84
timestamp 1679581782
transform 1 0 79680 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_91
timestamp 1679581782
transform 1 0 80352 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_98
timestamp 1679581782
transform 1 0 81024 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_105
timestamp 1679581782
transform 1 0 81696 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_112
timestamp 1679581782
transform 1 0 82368 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_119
timestamp 1679581782
transform 1 0 83040 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_126
timestamp 1679581782
transform 1 0 83712 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_133
timestamp 1679581782
transform 1 0 84384 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_140
timestamp 1679581782
transform 1 0 85056 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_147
timestamp 1679581782
transform 1 0 85728 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_154
timestamp 1679581782
transform 1 0 86400 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_161
timestamp 1679581782
transform 1 0 87072 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_168
timestamp 1679581782
transform 1 0 87744 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_175
timestamp 1679581782
transform 1 0 88416 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_182
timestamp 1679581782
transform 1 0 89088 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_189
timestamp 1679581782
transform 1 0 89760 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_196
timestamp 1679581782
transform 1 0 90432 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_203
timestamp 1679581782
transform 1 0 91104 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_210
timestamp 1679581782
transform 1 0 91776 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_217
timestamp 1679581782
transform 1 0 92448 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_224
timestamp 1679581782
transform 1 0 93120 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_231
timestamp 1679581782
transform 1 0 93792 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_238
timestamp 1679581782
transform 1 0 94464 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_245
timestamp 1679581782
transform 1 0 95136 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_252
timestamp 1679581782
transform 1 0 95808 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_259
timestamp 1679581782
transform 1 0 96480 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_266
timestamp 1679581782
transform 1 0 97152 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_273
timestamp 1679581782
transform 1 0 97824 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_280
timestamp 1679581782
transform 1 0 98496 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_287
timestamp 1679581782
transform 1 0 99168 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_294
timestamp 1679581782
transform 1 0 99840 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_301
timestamp 1679581782
transform 1 0 100512 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_308
timestamp 1679581782
transform 1 0 101184 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_315
timestamp 1679581782
transform 1 0 101856 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_322
timestamp 1679581782
transform 1 0 102528 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_329
timestamp 1679581782
transform 1 0 103200 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_336
timestamp 1679581782
transform 1 0 103872 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_343
timestamp 1679581782
transform 1 0 104544 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_350
timestamp 1679581782
transform 1 0 105216 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_357
timestamp 1679581782
transform 1 0 105888 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_364
timestamp 1679581782
transform 1 0 106560 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_371
timestamp 1679581782
transform 1 0 107232 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_378
timestamp 1679581782
transform 1 0 107904 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_385
timestamp 1679581782
transform 1 0 108576 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_392
timestamp 1679581782
transform 1 0 109248 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_399
timestamp 1679581782
transform 1 0 109920 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_406
timestamp 1679581782
transform 1 0 110592 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_413
timestamp 1679581782
transform 1 0 111264 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_420
timestamp 1679581782
transform 1 0 111936 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_427
timestamp 1679581782
transform 1 0 112608 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_434
timestamp 1679581782
transform 1 0 113280 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_441
timestamp 1679581782
transform 1 0 113952 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_448
timestamp 1679581782
transform 1 0 114624 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_455
timestamp 1679581782
transform 1 0 115296 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_462
timestamp 1679581782
transform 1 0 115968 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_469
timestamp 1679581782
transform 1 0 116640 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_476
timestamp 1679581782
transform 1 0 117312 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_483
timestamp 1679581782
transform 1 0 117984 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_490
timestamp 1679581782
transform 1 0 118656 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_497
timestamp 1679581782
transform 1 0 119328 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_504
timestamp 1679581782
transform 1 0 120000 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_511
timestamp 1679581782
transform 1 0 120672 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_518
timestamp 1679581782
transform 1 0 121344 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_525
timestamp 1679581782
transform 1 0 122016 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_532
timestamp 1679581782
transform 1 0 122688 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_539
timestamp 1679581782
transform 1 0 123360 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_546
timestamp 1679581782
transform 1 0 124032 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_553
timestamp 1679581782
transform 1 0 124704 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_560
timestamp 1679581782
transform 1 0 125376 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_567
timestamp 1679581782
transform 1 0 126048 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_574
timestamp 1679581782
transform 1 0 126720 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_581
timestamp 1679581782
transform 1 0 127392 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_588
timestamp 1679581782
transform 1 0 128064 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_595
timestamp 1679581782
transform 1 0 128736 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_602
timestamp 1679581782
transform 1 0 129408 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_609
timestamp 1679581782
transform 1 0 130080 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_616
timestamp 1679581782
transform 1 0 130752 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_623
timestamp 1679581782
transform 1 0 131424 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_630
timestamp 1679581782
transform 1 0 132096 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_637
timestamp 1679581782
transform 1 0 132768 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_644
timestamp 1679581782
transform 1 0 133440 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_651
timestamp 1679581782
transform 1 0 134112 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_658
timestamp 1679581782
transform 1 0 134784 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_665
timestamp 1679581782
transform 1 0 135456 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_672
timestamp 1679581782
transform 1 0 136128 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_679
timestamp 1679581782
transform 1 0 136800 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_686
timestamp 1679581782
transform 1 0 137472 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_693
timestamp 1679581782
transform 1 0 138144 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_700
timestamp 1679581782
transform 1 0 138816 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_707
timestamp 1679581782
transform 1 0 139488 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_714
timestamp 1679581782
transform 1 0 140160 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_721
timestamp 1679581782
transform 1 0 140832 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_728
timestamp 1679581782
transform 1 0 141504 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_735
timestamp 1679581782
transform 1 0 142176 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_742
timestamp 1679581782
transform 1 0 142848 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_749
timestamp 1679581782
transform 1 0 143520 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_756
timestamp 1679581782
transform 1 0 144192 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_763
timestamp 1679581782
transform 1 0 144864 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_770
timestamp 1679581782
transform 1 0 145536 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_777
timestamp 1679581782
transform 1 0 146208 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_784
timestamp 1679581782
transform 1 0 146880 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_791
timestamp 1679581782
transform 1 0 147552 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_798
timestamp 1679581782
transform 1 0 148224 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_805
timestamp 1679581782
transform 1 0 148896 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_812
timestamp 1679581782
transform 1 0 149568 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_819
timestamp 1679581782
transform 1 0 150240 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_826
timestamp 1679581782
transform 1 0 150912 0 -1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_833
timestamp 1679581782
transform 1 0 151584 0 -1 82404
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_840
timestamp 1677579658
transform 1 0 152256 0 -1 82404
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_0
timestamp 1679581782
transform 1 0 71616 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_7
timestamp 1679581782
transform 1 0 72288 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_14
timestamp 1679581782
transform 1 0 72960 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_21
timestamp 1679581782
transform 1 0 73632 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_28
timestamp 1679581782
transform 1 0 74304 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_35
timestamp 1679581782
transform 1 0 74976 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_42
timestamp 1679581782
transform 1 0 75648 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_49
timestamp 1679581782
transform 1 0 76320 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_56
timestamp 1679581782
transform 1 0 76992 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_63
timestamp 1679581782
transform 1 0 77664 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_70
timestamp 1679581782
transform 1 0 78336 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_77
timestamp 1679581782
transform 1 0 79008 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_84
timestamp 1679581782
transform 1 0 79680 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_91
timestamp 1679581782
transform 1 0 80352 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_98
timestamp 1679581782
transform 1 0 81024 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_105
timestamp 1679581782
transform 1 0 81696 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_112
timestamp 1679581782
transform 1 0 82368 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_119
timestamp 1679581782
transform 1 0 83040 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_126
timestamp 1679581782
transform 1 0 83712 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_133
timestamp 1679581782
transform 1 0 84384 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_140
timestamp 1679581782
transform 1 0 85056 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_147
timestamp 1679581782
transform 1 0 85728 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_154
timestamp 1679581782
transform 1 0 86400 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_161
timestamp 1679581782
transform 1 0 87072 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_168
timestamp 1679581782
transform 1 0 87744 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_175
timestamp 1679581782
transform 1 0 88416 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_182
timestamp 1679581782
transform 1 0 89088 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_189
timestamp 1679581782
transform 1 0 89760 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_196
timestamp 1679581782
transform 1 0 90432 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_203
timestamp 1679581782
transform 1 0 91104 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_210
timestamp 1679581782
transform 1 0 91776 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_217
timestamp 1679581782
transform 1 0 92448 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_224
timestamp 1679581782
transform 1 0 93120 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_231
timestamp 1679581782
transform 1 0 93792 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_238
timestamp 1679581782
transform 1 0 94464 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_245
timestamp 1679581782
transform 1 0 95136 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_252
timestamp 1679581782
transform 1 0 95808 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_259
timestamp 1679581782
transform 1 0 96480 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_266
timestamp 1679581782
transform 1 0 97152 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_273
timestamp 1679581782
transform 1 0 97824 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_280
timestamp 1679581782
transform 1 0 98496 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_287
timestamp 1679581782
transform 1 0 99168 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_294
timestamp 1679581782
transform 1 0 99840 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_301
timestamp 1679581782
transform 1 0 100512 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_308
timestamp 1679581782
transform 1 0 101184 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_315
timestamp 1679581782
transform 1 0 101856 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_322
timestamp 1679581782
transform 1 0 102528 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_329
timestamp 1679581782
transform 1 0 103200 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_336
timestamp 1679581782
transform 1 0 103872 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_343
timestamp 1679581782
transform 1 0 104544 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_350
timestamp 1679581782
transform 1 0 105216 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_357
timestamp 1679581782
transform 1 0 105888 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_364
timestamp 1679581782
transform 1 0 106560 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_371
timestamp 1679581782
transform 1 0 107232 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_378
timestamp 1679581782
transform 1 0 107904 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_385
timestamp 1679581782
transform 1 0 108576 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_392
timestamp 1679581782
transform 1 0 109248 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_399
timestamp 1679581782
transform 1 0 109920 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_406
timestamp 1679581782
transform 1 0 110592 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_413
timestamp 1679581782
transform 1 0 111264 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_420
timestamp 1679581782
transform 1 0 111936 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_427
timestamp 1679581782
transform 1 0 112608 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_434
timestamp 1679581782
transform 1 0 113280 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_441
timestamp 1679581782
transform 1 0 113952 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_448
timestamp 1679581782
transform 1 0 114624 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_455
timestamp 1679581782
transform 1 0 115296 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_462
timestamp 1679581782
transform 1 0 115968 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_469
timestamp 1679581782
transform 1 0 116640 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_476
timestamp 1679581782
transform 1 0 117312 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_483
timestamp 1679581782
transform 1 0 117984 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_490
timestamp 1679581782
transform 1 0 118656 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_497
timestamp 1679581782
transform 1 0 119328 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_504
timestamp 1679581782
transform 1 0 120000 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_511
timestamp 1679581782
transform 1 0 120672 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_518
timestamp 1679581782
transform 1 0 121344 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_525
timestamp 1679581782
transform 1 0 122016 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_532
timestamp 1679581782
transform 1 0 122688 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_539
timestamp 1679581782
transform 1 0 123360 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_546
timestamp 1679581782
transform 1 0 124032 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_553
timestamp 1679581782
transform 1 0 124704 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_560
timestamp 1679581782
transform 1 0 125376 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_567
timestamp 1679581782
transform 1 0 126048 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_574
timestamp 1679581782
transform 1 0 126720 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_581
timestamp 1679581782
transform 1 0 127392 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_588
timestamp 1679581782
transform 1 0 128064 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_595
timestamp 1679581782
transform 1 0 128736 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_602
timestamp 1679581782
transform 1 0 129408 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_609
timestamp 1679581782
transform 1 0 130080 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_616
timestamp 1679581782
transform 1 0 130752 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_623
timestamp 1679581782
transform 1 0 131424 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_630
timestamp 1679581782
transform 1 0 132096 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_637
timestamp 1679581782
transform 1 0 132768 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_644
timestamp 1679581782
transform 1 0 133440 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_651
timestamp 1679581782
transform 1 0 134112 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_658
timestamp 1679581782
transform 1 0 134784 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_665
timestamp 1679581782
transform 1 0 135456 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_672
timestamp 1679581782
transform 1 0 136128 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_679
timestamp 1679581782
transform 1 0 136800 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_686
timestamp 1679581782
transform 1 0 137472 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_693
timestamp 1679581782
transform 1 0 138144 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_700
timestamp 1679581782
transform 1 0 138816 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_707
timestamp 1679581782
transform 1 0 139488 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_714
timestamp 1679581782
transform 1 0 140160 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_721
timestamp 1679581782
transform 1 0 140832 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_728
timestamp 1679581782
transform 1 0 141504 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_735
timestamp 1679581782
transform 1 0 142176 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_742
timestamp 1679581782
transform 1 0 142848 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_749
timestamp 1679581782
transform 1 0 143520 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_756
timestamp 1679581782
transform 1 0 144192 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_763
timestamp 1679581782
transform 1 0 144864 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_770
timestamp 1679581782
transform 1 0 145536 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_777
timestamp 1679581782
transform 1 0 146208 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_784
timestamp 1679581782
transform 1 0 146880 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_791
timestamp 1679581782
transform 1 0 147552 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_798
timestamp 1679581782
transform 1 0 148224 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_805
timestamp 1679581782
transform 1 0 148896 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_812
timestamp 1679581782
transform 1 0 149568 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_819
timestamp 1679581782
transform 1 0 150240 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_826
timestamp 1679581782
transform 1 0 150912 0 1 82404
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_833
timestamp 1679581782
transform 1 0 151584 0 1 82404
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_840
timestamp 1677579658
transform 1 0 152256 0 1 82404
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_0
timestamp 1679581782
transform 1 0 71616 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_7
timestamp 1679581782
transform 1 0 72288 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_14
timestamp 1679581782
transform 1 0 72960 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_21
timestamp 1679581782
transform 1 0 73632 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_28
timestamp 1679581782
transform 1 0 74304 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_35
timestamp 1679581782
transform 1 0 74976 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_42
timestamp 1679581782
transform 1 0 75648 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_49
timestamp 1679581782
transform 1 0 76320 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_56
timestamp 1679581782
transform 1 0 76992 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_63
timestamp 1679581782
transform 1 0 77664 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_70
timestamp 1679581782
transform 1 0 78336 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_77
timestamp 1679581782
transform 1 0 79008 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_84
timestamp 1679581782
transform 1 0 79680 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_91
timestamp 1679581782
transform 1 0 80352 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_98
timestamp 1679581782
transform 1 0 81024 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_105
timestamp 1679581782
transform 1 0 81696 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_112
timestamp 1679581782
transform 1 0 82368 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_119
timestamp 1679581782
transform 1 0 83040 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_126
timestamp 1679581782
transform 1 0 83712 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_133
timestamp 1679581782
transform 1 0 84384 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_140
timestamp 1679581782
transform 1 0 85056 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_147
timestamp 1679581782
transform 1 0 85728 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_154
timestamp 1679581782
transform 1 0 86400 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_161
timestamp 1679581782
transform 1 0 87072 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_168
timestamp 1679581782
transform 1 0 87744 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_175
timestamp 1679581782
transform 1 0 88416 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_182
timestamp 1679581782
transform 1 0 89088 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_189
timestamp 1679581782
transform 1 0 89760 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_196
timestamp 1679581782
transform 1 0 90432 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_203
timestamp 1679581782
transform 1 0 91104 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_210
timestamp 1679581782
transform 1 0 91776 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_217
timestamp 1679581782
transform 1 0 92448 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_224
timestamp 1679581782
transform 1 0 93120 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_231
timestamp 1679581782
transform 1 0 93792 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_238
timestamp 1679581782
transform 1 0 94464 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_245
timestamp 1679581782
transform 1 0 95136 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_252
timestamp 1679581782
transform 1 0 95808 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_259
timestamp 1679581782
transform 1 0 96480 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_266
timestamp 1679581782
transform 1 0 97152 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_273
timestamp 1679581782
transform 1 0 97824 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_280
timestamp 1679581782
transform 1 0 98496 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_287
timestamp 1679581782
transform 1 0 99168 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_294
timestamp 1679581782
transform 1 0 99840 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_301
timestamp 1679581782
transform 1 0 100512 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_308
timestamp 1679581782
transform 1 0 101184 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_315
timestamp 1679581782
transform 1 0 101856 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_322
timestamp 1679581782
transform 1 0 102528 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_329
timestamp 1679581782
transform 1 0 103200 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_336
timestamp 1679581782
transform 1 0 103872 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_343
timestamp 1679581782
transform 1 0 104544 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_350
timestamp 1679581782
transform 1 0 105216 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_357
timestamp 1679581782
transform 1 0 105888 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_364
timestamp 1679581782
transform 1 0 106560 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_371
timestamp 1679581782
transform 1 0 107232 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_378
timestamp 1679581782
transform 1 0 107904 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_385
timestamp 1679581782
transform 1 0 108576 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_392
timestamp 1679581782
transform 1 0 109248 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_399
timestamp 1679581782
transform 1 0 109920 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_406
timestamp 1679581782
transform 1 0 110592 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_413
timestamp 1679581782
transform 1 0 111264 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_420
timestamp 1679581782
transform 1 0 111936 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_427
timestamp 1679581782
transform 1 0 112608 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_434
timestamp 1679581782
transform 1 0 113280 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_441
timestamp 1679581782
transform 1 0 113952 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_448
timestamp 1679581782
transform 1 0 114624 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_455
timestamp 1679581782
transform 1 0 115296 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_462
timestamp 1679581782
transform 1 0 115968 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_469
timestamp 1679581782
transform 1 0 116640 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_476
timestamp 1679581782
transform 1 0 117312 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_483
timestamp 1679581782
transform 1 0 117984 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_490
timestamp 1679581782
transform 1 0 118656 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_497
timestamp 1679581782
transform 1 0 119328 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_504
timestamp 1679581782
transform 1 0 120000 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_511
timestamp 1679581782
transform 1 0 120672 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_518
timestamp 1679581782
transform 1 0 121344 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_525
timestamp 1679581782
transform 1 0 122016 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_532
timestamp 1679581782
transform 1 0 122688 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_539
timestamp 1679581782
transform 1 0 123360 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_546
timestamp 1679581782
transform 1 0 124032 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_553
timestamp 1679581782
transform 1 0 124704 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_560
timestamp 1679581782
transform 1 0 125376 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_567
timestamp 1679581782
transform 1 0 126048 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_574
timestamp 1679581782
transform 1 0 126720 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_581
timestamp 1679581782
transform 1 0 127392 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_588
timestamp 1679581782
transform 1 0 128064 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_595
timestamp 1679581782
transform 1 0 128736 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_602
timestamp 1679581782
transform 1 0 129408 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_609
timestamp 1679581782
transform 1 0 130080 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_616
timestamp 1679581782
transform 1 0 130752 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_623
timestamp 1679581782
transform 1 0 131424 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_630
timestamp 1679581782
transform 1 0 132096 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_637
timestamp 1679581782
transform 1 0 132768 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_644
timestamp 1679581782
transform 1 0 133440 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_651
timestamp 1679581782
transform 1 0 134112 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_658
timestamp 1679581782
transform 1 0 134784 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_665
timestamp 1679581782
transform 1 0 135456 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_672
timestamp 1679581782
transform 1 0 136128 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_679
timestamp 1679581782
transform 1 0 136800 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_686
timestamp 1679581782
transform 1 0 137472 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_693
timestamp 1679581782
transform 1 0 138144 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_700
timestamp 1679581782
transform 1 0 138816 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_707
timestamp 1679581782
transform 1 0 139488 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_714
timestamp 1679581782
transform 1 0 140160 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_721
timestamp 1679581782
transform 1 0 140832 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_728
timestamp 1679581782
transform 1 0 141504 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_735
timestamp 1679581782
transform 1 0 142176 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_742
timestamp 1679581782
transform 1 0 142848 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_749
timestamp 1679581782
transform 1 0 143520 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_756
timestamp 1679581782
transform 1 0 144192 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_763
timestamp 1679581782
transform 1 0 144864 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_770
timestamp 1679581782
transform 1 0 145536 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_777
timestamp 1679581782
transform 1 0 146208 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_784
timestamp 1679581782
transform 1 0 146880 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_791
timestamp 1679581782
transform 1 0 147552 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_798
timestamp 1679581782
transform 1 0 148224 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_805
timestamp 1679581782
transform 1 0 148896 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_812
timestamp 1679581782
transform 1 0 149568 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_819
timestamp 1679581782
transform 1 0 150240 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_826
timestamp 1679581782
transform 1 0 150912 0 -1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_833
timestamp 1679581782
transform 1 0 151584 0 -1 83916
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_840
timestamp 1677579658
transform 1 0 152256 0 -1 83916
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_0
timestamp 1679581782
transform 1 0 71616 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_7
timestamp 1679581782
transform 1 0 72288 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_14
timestamp 1679581782
transform 1 0 72960 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_21
timestamp 1679581782
transform 1 0 73632 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_28
timestamp 1679581782
transform 1 0 74304 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_35
timestamp 1679581782
transform 1 0 74976 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_42
timestamp 1679581782
transform 1 0 75648 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_49
timestamp 1679581782
transform 1 0 76320 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_56
timestamp 1679581782
transform 1 0 76992 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_63
timestamp 1679581782
transform 1 0 77664 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_70
timestamp 1679581782
transform 1 0 78336 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_77
timestamp 1679581782
transform 1 0 79008 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_84
timestamp 1679581782
transform 1 0 79680 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_91
timestamp 1679581782
transform 1 0 80352 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_98
timestamp 1679581782
transform 1 0 81024 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_105
timestamp 1679581782
transform 1 0 81696 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_112
timestamp 1679581782
transform 1 0 82368 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_119
timestamp 1679581782
transform 1 0 83040 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_126
timestamp 1679581782
transform 1 0 83712 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_133
timestamp 1679581782
transform 1 0 84384 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_140
timestamp 1679581782
transform 1 0 85056 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_147
timestamp 1679581782
transform 1 0 85728 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_154
timestamp 1679581782
transform 1 0 86400 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_161
timestamp 1679581782
transform 1 0 87072 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_168
timestamp 1679581782
transform 1 0 87744 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_175
timestamp 1679581782
transform 1 0 88416 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_182
timestamp 1679581782
transform 1 0 89088 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_189
timestamp 1679581782
transform 1 0 89760 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_196
timestamp 1679581782
transform 1 0 90432 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_203
timestamp 1679581782
transform 1 0 91104 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_210
timestamp 1679581782
transform 1 0 91776 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_217
timestamp 1679581782
transform 1 0 92448 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_224
timestamp 1679581782
transform 1 0 93120 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_231
timestamp 1679581782
transform 1 0 93792 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_238
timestamp 1679581782
transform 1 0 94464 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_245
timestamp 1679581782
transform 1 0 95136 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_252
timestamp 1679581782
transform 1 0 95808 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_259
timestamp 1679581782
transform 1 0 96480 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_266
timestamp 1679581782
transform 1 0 97152 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_273
timestamp 1679581782
transform 1 0 97824 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_280
timestamp 1679581782
transform 1 0 98496 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_287
timestamp 1679581782
transform 1 0 99168 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_294
timestamp 1679581782
transform 1 0 99840 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_301
timestamp 1679581782
transform 1 0 100512 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_308
timestamp 1679581782
transform 1 0 101184 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_315
timestamp 1679581782
transform 1 0 101856 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_322
timestamp 1679581782
transform 1 0 102528 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_329
timestamp 1679581782
transform 1 0 103200 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_336
timestamp 1679581782
transform 1 0 103872 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_343
timestamp 1679581782
transform 1 0 104544 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_350
timestamp 1679581782
transform 1 0 105216 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_357
timestamp 1679581782
transform 1 0 105888 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_364
timestamp 1679581782
transform 1 0 106560 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_371
timestamp 1679581782
transform 1 0 107232 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_378
timestamp 1679581782
transform 1 0 107904 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_385
timestamp 1679581782
transform 1 0 108576 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_392
timestamp 1679581782
transform 1 0 109248 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_399
timestamp 1679581782
transform 1 0 109920 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_406
timestamp 1679581782
transform 1 0 110592 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_413
timestamp 1679581782
transform 1 0 111264 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_420
timestamp 1679581782
transform 1 0 111936 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_427
timestamp 1679581782
transform 1 0 112608 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_434
timestamp 1679581782
transform 1 0 113280 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_441
timestamp 1679581782
transform 1 0 113952 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_448
timestamp 1679581782
transform 1 0 114624 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_455
timestamp 1679581782
transform 1 0 115296 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_462
timestamp 1679581782
transform 1 0 115968 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_469
timestamp 1679581782
transform 1 0 116640 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_476
timestamp 1679581782
transform 1 0 117312 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_483
timestamp 1679581782
transform 1 0 117984 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_490
timestamp 1679581782
transform 1 0 118656 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_497
timestamp 1679581782
transform 1 0 119328 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_504
timestamp 1679581782
transform 1 0 120000 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_511
timestamp 1679581782
transform 1 0 120672 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_518
timestamp 1679581782
transform 1 0 121344 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_525
timestamp 1679581782
transform 1 0 122016 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_532
timestamp 1679581782
transform 1 0 122688 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_539
timestamp 1679581782
transform 1 0 123360 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_546
timestamp 1679581782
transform 1 0 124032 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_553
timestamp 1679581782
transform 1 0 124704 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_560
timestamp 1679581782
transform 1 0 125376 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_567
timestamp 1679581782
transform 1 0 126048 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_574
timestamp 1679581782
transform 1 0 126720 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_581
timestamp 1679581782
transform 1 0 127392 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_588
timestamp 1679581782
transform 1 0 128064 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_595
timestamp 1679581782
transform 1 0 128736 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_602
timestamp 1679581782
transform 1 0 129408 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_609
timestamp 1679581782
transform 1 0 130080 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_616
timestamp 1679581782
transform 1 0 130752 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_623
timestamp 1679581782
transform 1 0 131424 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_630
timestamp 1679581782
transform 1 0 132096 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_637
timestamp 1679581782
transform 1 0 132768 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_644
timestamp 1679581782
transform 1 0 133440 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_651
timestamp 1679581782
transform 1 0 134112 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_658
timestamp 1679581782
transform 1 0 134784 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_665
timestamp 1679581782
transform 1 0 135456 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_672
timestamp 1679581782
transform 1 0 136128 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_679
timestamp 1679581782
transform 1 0 136800 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_686
timestamp 1679581782
transform 1 0 137472 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_693
timestamp 1679581782
transform 1 0 138144 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_700
timestamp 1679581782
transform 1 0 138816 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_707
timestamp 1679581782
transform 1 0 139488 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_714
timestamp 1679581782
transform 1 0 140160 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_721
timestamp 1679581782
transform 1 0 140832 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_728
timestamp 1679581782
transform 1 0 141504 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_735
timestamp 1679581782
transform 1 0 142176 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_742
timestamp 1679581782
transform 1 0 142848 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_749
timestamp 1679581782
transform 1 0 143520 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_756
timestamp 1679581782
transform 1 0 144192 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_763
timestamp 1679581782
transform 1 0 144864 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_770
timestamp 1679581782
transform 1 0 145536 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_777
timestamp 1679581782
transform 1 0 146208 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_784
timestamp 1679581782
transform 1 0 146880 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_791
timestamp 1679581782
transform 1 0 147552 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_798
timestamp 1679581782
transform 1 0 148224 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_805
timestamp 1679581782
transform 1 0 148896 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_812
timestamp 1679581782
transform 1 0 149568 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_819
timestamp 1679581782
transform 1 0 150240 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_826
timestamp 1679581782
transform 1 0 150912 0 1 83916
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_833
timestamp 1679581782
transform 1 0 151584 0 1 83916
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_840
timestamp 1677579658
transform 1 0 152256 0 1 83916
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679581782
transform 1 0 71616 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_7
timestamp 1679581782
transform 1 0 72288 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_14
timestamp 1679581782
transform 1 0 72960 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_21
timestamp 1679581782
transform 1 0 73632 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_28
timestamp 1679581782
transform 1 0 74304 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_35
timestamp 1679581782
transform 1 0 74976 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_42
timestamp 1679581782
transform 1 0 75648 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_49
timestamp 1679581782
transform 1 0 76320 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_56
timestamp 1679581782
transform 1 0 76992 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_63
timestamp 1679581782
transform 1 0 77664 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_70
timestamp 1679581782
transform 1 0 78336 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_77
timestamp 1679581782
transform 1 0 79008 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_84
timestamp 1679581782
transform 1 0 79680 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_91
timestamp 1679581782
transform 1 0 80352 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_98
timestamp 1679581782
transform 1 0 81024 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_105
timestamp 1679581782
transform 1 0 81696 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_112
timestamp 1679581782
transform 1 0 82368 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_119
timestamp 1679581782
transform 1 0 83040 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_126
timestamp 1679581782
transform 1 0 83712 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_133
timestamp 1679581782
transform 1 0 84384 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_140
timestamp 1679581782
transform 1 0 85056 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_147
timestamp 1679581782
transform 1 0 85728 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_154
timestamp 1679581782
transform 1 0 86400 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_161
timestamp 1679581782
transform 1 0 87072 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_168
timestamp 1679581782
transform 1 0 87744 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_175
timestamp 1679581782
transform 1 0 88416 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_182
timestamp 1679581782
transform 1 0 89088 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_189
timestamp 1679581782
transform 1 0 89760 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_196
timestamp 1679581782
transform 1 0 90432 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_203
timestamp 1679581782
transform 1 0 91104 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_210
timestamp 1679581782
transform 1 0 91776 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_217
timestamp 1679581782
transform 1 0 92448 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_224
timestamp 1679581782
transform 1 0 93120 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_231
timestamp 1679581782
transform 1 0 93792 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_238
timestamp 1679581782
transform 1 0 94464 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_245
timestamp 1679581782
transform 1 0 95136 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_252
timestamp 1679581782
transform 1 0 95808 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_259
timestamp 1679581782
transform 1 0 96480 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_266
timestamp 1679581782
transform 1 0 97152 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_273
timestamp 1679581782
transform 1 0 97824 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_280
timestamp 1679581782
transform 1 0 98496 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_287
timestamp 1679581782
transform 1 0 99168 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_294
timestamp 1679581782
transform 1 0 99840 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_301
timestamp 1679581782
transform 1 0 100512 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_308
timestamp 1679581782
transform 1 0 101184 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_315
timestamp 1679581782
transform 1 0 101856 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_322
timestamp 1679581782
transform 1 0 102528 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_329
timestamp 1679581782
transform 1 0 103200 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_336
timestamp 1679581782
transform 1 0 103872 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_343
timestamp 1679581782
transform 1 0 104544 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_350
timestamp 1679581782
transform 1 0 105216 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_357
timestamp 1679581782
transform 1 0 105888 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_364
timestamp 1679581782
transform 1 0 106560 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_371
timestamp 1679581782
transform 1 0 107232 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_378
timestamp 1679581782
transform 1 0 107904 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_385
timestamp 1679581782
transform 1 0 108576 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_392
timestamp 1679581782
transform 1 0 109248 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_399
timestamp 1679581782
transform 1 0 109920 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_406
timestamp 1679581782
transform 1 0 110592 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_413
timestamp 1679581782
transform 1 0 111264 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_420
timestamp 1679581782
transform 1 0 111936 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_427
timestamp 1679581782
transform 1 0 112608 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_434
timestamp 1679581782
transform 1 0 113280 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_441
timestamp 1679581782
transform 1 0 113952 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_448
timestamp 1679581782
transform 1 0 114624 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_455
timestamp 1679581782
transform 1 0 115296 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_462
timestamp 1679581782
transform 1 0 115968 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_469
timestamp 1679581782
transform 1 0 116640 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_476
timestamp 1679581782
transform 1 0 117312 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_483
timestamp 1679581782
transform 1 0 117984 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_490
timestamp 1679581782
transform 1 0 118656 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_497
timestamp 1679581782
transform 1 0 119328 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_504
timestamp 1679581782
transform 1 0 120000 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_511
timestamp 1679581782
transform 1 0 120672 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_518
timestamp 1679581782
transform 1 0 121344 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_525
timestamp 1679581782
transform 1 0 122016 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_532
timestamp 1679581782
transform 1 0 122688 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_539
timestamp 1679581782
transform 1 0 123360 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_546
timestamp 1679581782
transform 1 0 124032 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_553
timestamp 1679581782
transform 1 0 124704 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_560
timestamp 1679581782
transform 1 0 125376 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_567
timestamp 1679581782
transform 1 0 126048 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_574
timestamp 1679581782
transform 1 0 126720 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_581
timestamp 1679581782
transform 1 0 127392 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_588
timestamp 1679581782
transform 1 0 128064 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_595
timestamp 1679581782
transform 1 0 128736 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_602
timestamp 1679581782
transform 1 0 129408 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_609
timestamp 1679581782
transform 1 0 130080 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_616
timestamp 1679581782
transform 1 0 130752 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_623
timestamp 1679581782
transform 1 0 131424 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_630
timestamp 1679581782
transform 1 0 132096 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_637
timestamp 1679581782
transform 1 0 132768 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_644
timestamp 1679581782
transform 1 0 133440 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_651
timestamp 1679581782
transform 1 0 134112 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_658
timestamp 1679581782
transform 1 0 134784 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_665
timestamp 1679581782
transform 1 0 135456 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_672
timestamp 1679581782
transform 1 0 136128 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_679
timestamp 1679581782
transform 1 0 136800 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_686
timestamp 1679581782
transform 1 0 137472 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_693
timestamp 1679581782
transform 1 0 138144 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_700
timestamp 1679581782
transform 1 0 138816 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_707
timestamp 1679581782
transform 1 0 139488 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_714
timestamp 1679581782
transform 1 0 140160 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_721
timestamp 1679581782
transform 1 0 140832 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_728
timestamp 1679581782
transform 1 0 141504 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_735
timestamp 1679581782
transform 1 0 142176 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_742
timestamp 1679581782
transform 1 0 142848 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_749
timestamp 1679581782
transform 1 0 143520 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_756
timestamp 1679581782
transform 1 0 144192 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_763
timestamp 1679581782
transform 1 0 144864 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_770
timestamp 1679581782
transform 1 0 145536 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_777
timestamp 1679581782
transform 1 0 146208 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_784
timestamp 1679581782
transform 1 0 146880 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_791
timestamp 1679581782
transform 1 0 147552 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_798
timestamp 1679581782
transform 1 0 148224 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_805
timestamp 1679581782
transform 1 0 148896 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_812
timestamp 1679581782
transform 1 0 149568 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_819
timestamp 1679581782
transform 1 0 150240 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_826
timestamp 1679581782
transform 1 0 150912 0 -1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_833
timestamp 1679581782
transform 1 0 151584 0 -1 85428
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_840
timestamp 1677579658
transform 1 0 152256 0 -1 85428
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_0
timestamp 1679581782
transform 1 0 71616 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_7
timestamp 1679581782
transform 1 0 72288 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_14
timestamp 1679581782
transform 1 0 72960 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_21
timestamp 1679581782
transform 1 0 73632 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_28
timestamp 1679581782
transform 1 0 74304 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_35
timestamp 1679581782
transform 1 0 74976 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_42
timestamp 1679581782
transform 1 0 75648 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_49
timestamp 1679581782
transform 1 0 76320 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_56
timestamp 1679581782
transform 1 0 76992 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_63
timestamp 1679581782
transform 1 0 77664 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_70
timestamp 1679581782
transform 1 0 78336 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_77
timestamp 1679581782
transform 1 0 79008 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_84
timestamp 1679581782
transform 1 0 79680 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_91
timestamp 1679581782
transform 1 0 80352 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_98
timestamp 1679581782
transform 1 0 81024 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_105
timestamp 1679581782
transform 1 0 81696 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_112
timestamp 1679581782
transform 1 0 82368 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_119
timestamp 1679581782
transform 1 0 83040 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_126
timestamp 1679581782
transform 1 0 83712 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_133
timestamp 1679581782
transform 1 0 84384 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_140
timestamp 1679581782
transform 1 0 85056 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_147
timestamp 1679581782
transform 1 0 85728 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_154
timestamp 1679581782
transform 1 0 86400 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_161
timestamp 1679581782
transform 1 0 87072 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_168
timestamp 1679581782
transform 1 0 87744 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_175
timestamp 1679581782
transform 1 0 88416 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_182
timestamp 1679581782
transform 1 0 89088 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_189
timestamp 1679581782
transform 1 0 89760 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_196
timestamp 1679581782
transform 1 0 90432 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_203
timestamp 1679581782
transform 1 0 91104 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_210
timestamp 1679581782
transform 1 0 91776 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_217
timestamp 1679581782
transform 1 0 92448 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_224
timestamp 1679581782
transform 1 0 93120 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_231
timestamp 1679581782
transform 1 0 93792 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_238
timestamp 1679581782
transform 1 0 94464 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_245
timestamp 1679581782
transform 1 0 95136 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_252
timestamp 1679581782
transform 1 0 95808 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_259
timestamp 1679581782
transform 1 0 96480 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_266
timestamp 1679581782
transform 1 0 97152 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_273
timestamp 1679581782
transform 1 0 97824 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_280
timestamp 1679581782
transform 1 0 98496 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_287
timestamp 1679581782
transform 1 0 99168 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_294
timestamp 1679581782
transform 1 0 99840 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_301
timestamp 1679581782
transform 1 0 100512 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_308
timestamp 1679581782
transform 1 0 101184 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_315
timestamp 1679581782
transform 1 0 101856 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_322
timestamp 1679581782
transform 1 0 102528 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_329
timestamp 1679581782
transform 1 0 103200 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_336
timestamp 1679581782
transform 1 0 103872 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_343
timestamp 1679581782
transform 1 0 104544 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_350
timestamp 1679581782
transform 1 0 105216 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_357
timestamp 1679581782
transform 1 0 105888 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_364
timestamp 1679581782
transform 1 0 106560 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_371
timestamp 1679581782
transform 1 0 107232 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_378
timestamp 1679581782
transform 1 0 107904 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_385
timestamp 1679581782
transform 1 0 108576 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_392
timestamp 1679581782
transform 1 0 109248 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_399
timestamp 1679581782
transform 1 0 109920 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_406
timestamp 1679581782
transform 1 0 110592 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_413
timestamp 1679581782
transform 1 0 111264 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_420
timestamp 1679581782
transform 1 0 111936 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_427
timestamp 1679581782
transform 1 0 112608 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_434
timestamp 1679581782
transform 1 0 113280 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_441
timestamp 1679581782
transform 1 0 113952 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_448
timestamp 1679581782
transform 1 0 114624 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_455
timestamp 1679581782
transform 1 0 115296 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_462
timestamp 1679581782
transform 1 0 115968 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_469
timestamp 1679581782
transform 1 0 116640 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_476
timestamp 1679581782
transform 1 0 117312 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_483
timestamp 1679581782
transform 1 0 117984 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_490
timestamp 1679581782
transform 1 0 118656 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_497
timestamp 1679581782
transform 1 0 119328 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_504
timestamp 1679581782
transform 1 0 120000 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_511
timestamp 1679581782
transform 1 0 120672 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_518
timestamp 1679581782
transform 1 0 121344 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_525
timestamp 1679581782
transform 1 0 122016 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_532
timestamp 1679581782
transform 1 0 122688 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_539
timestamp 1679581782
transform 1 0 123360 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_546
timestamp 1679581782
transform 1 0 124032 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_553
timestamp 1679581782
transform 1 0 124704 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_560
timestamp 1679581782
transform 1 0 125376 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_567
timestamp 1679581782
transform 1 0 126048 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_574
timestamp 1679581782
transform 1 0 126720 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_581
timestamp 1679581782
transform 1 0 127392 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_588
timestamp 1679581782
transform 1 0 128064 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_595
timestamp 1679581782
transform 1 0 128736 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_602
timestamp 1679581782
transform 1 0 129408 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_609
timestamp 1679581782
transform 1 0 130080 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_616
timestamp 1679581782
transform 1 0 130752 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_623
timestamp 1679581782
transform 1 0 131424 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_630
timestamp 1679581782
transform 1 0 132096 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_637
timestamp 1679581782
transform 1 0 132768 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_644
timestamp 1679581782
transform 1 0 133440 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_651
timestamp 1679581782
transform 1 0 134112 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_658
timestamp 1679581782
transform 1 0 134784 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_665
timestamp 1679581782
transform 1 0 135456 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_672
timestamp 1679581782
transform 1 0 136128 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_679
timestamp 1679581782
transform 1 0 136800 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_686
timestamp 1679581782
transform 1 0 137472 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_693
timestamp 1679581782
transform 1 0 138144 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_700
timestamp 1679581782
transform 1 0 138816 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_707
timestamp 1679581782
transform 1 0 139488 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_714
timestamp 1679581782
transform 1 0 140160 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_721
timestamp 1679581782
transform 1 0 140832 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_728
timestamp 1679581782
transform 1 0 141504 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_735
timestamp 1679581782
transform 1 0 142176 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_742
timestamp 1679581782
transform 1 0 142848 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_749
timestamp 1679581782
transform 1 0 143520 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_756
timestamp 1679581782
transform 1 0 144192 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_763
timestamp 1679581782
transform 1 0 144864 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_770
timestamp 1679581782
transform 1 0 145536 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_777
timestamp 1679581782
transform 1 0 146208 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_784
timestamp 1679581782
transform 1 0 146880 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_791
timestamp 1679581782
transform 1 0 147552 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_798
timestamp 1679581782
transform 1 0 148224 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_805
timestamp 1679581782
transform 1 0 148896 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_812
timestamp 1679581782
transform 1 0 149568 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_819
timestamp 1679581782
transform 1 0 150240 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_826
timestamp 1679581782
transform 1 0 150912 0 1 85428
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_833
timestamp 1679581782
transform 1 0 151584 0 1 85428
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_840
timestamp 1677579658
transform 1 0 152256 0 1 85428
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_0
timestamp 1679581782
transform 1 0 71616 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_7
timestamp 1679581782
transform 1 0 72288 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_14
timestamp 1679581782
transform 1 0 72960 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_21
timestamp 1679581782
transform 1 0 73632 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_28
timestamp 1679581782
transform 1 0 74304 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_35
timestamp 1679581782
transform 1 0 74976 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_42
timestamp 1679581782
transform 1 0 75648 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_49
timestamp 1679581782
transform 1 0 76320 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_56
timestamp 1679581782
transform 1 0 76992 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_63
timestamp 1679581782
transform 1 0 77664 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_70
timestamp 1679581782
transform 1 0 78336 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_77
timestamp 1679581782
transform 1 0 79008 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_84
timestamp 1679581782
transform 1 0 79680 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_91
timestamp 1679581782
transform 1 0 80352 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_98
timestamp 1679581782
transform 1 0 81024 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_105
timestamp 1679581782
transform 1 0 81696 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_112
timestamp 1679581782
transform 1 0 82368 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_119
timestamp 1679581782
transform 1 0 83040 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_126
timestamp 1679581782
transform 1 0 83712 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_133
timestamp 1679581782
transform 1 0 84384 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_140
timestamp 1679581782
transform 1 0 85056 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_147
timestamp 1679581782
transform 1 0 85728 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_154
timestamp 1679581782
transform 1 0 86400 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_161
timestamp 1679581782
transform 1 0 87072 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_168
timestamp 1679581782
transform 1 0 87744 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_175
timestamp 1679581782
transform 1 0 88416 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_182
timestamp 1679581782
transform 1 0 89088 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_189
timestamp 1679581782
transform 1 0 89760 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_196
timestamp 1679581782
transform 1 0 90432 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_203
timestamp 1679581782
transform 1 0 91104 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_210
timestamp 1679581782
transform 1 0 91776 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_217
timestamp 1679581782
transform 1 0 92448 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_224
timestamp 1679581782
transform 1 0 93120 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_231
timestamp 1679581782
transform 1 0 93792 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_238
timestamp 1679581782
transform 1 0 94464 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_245
timestamp 1679581782
transform 1 0 95136 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_252
timestamp 1679581782
transform 1 0 95808 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_259
timestamp 1679581782
transform 1 0 96480 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_266
timestamp 1679581782
transform 1 0 97152 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_273
timestamp 1679581782
transform 1 0 97824 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_280
timestamp 1679581782
transform 1 0 98496 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_287
timestamp 1679581782
transform 1 0 99168 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_294
timestamp 1679581782
transform 1 0 99840 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_301
timestamp 1679581782
transform 1 0 100512 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_308
timestamp 1679581782
transform 1 0 101184 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_315
timestamp 1679581782
transform 1 0 101856 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_322
timestamp 1679581782
transform 1 0 102528 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_329
timestamp 1679581782
transform 1 0 103200 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_336
timestamp 1679581782
transform 1 0 103872 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_343
timestamp 1679581782
transform 1 0 104544 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_350
timestamp 1679581782
transform 1 0 105216 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_357
timestamp 1679581782
transform 1 0 105888 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_364
timestamp 1679581782
transform 1 0 106560 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_371
timestamp 1679581782
transform 1 0 107232 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_378
timestamp 1679581782
transform 1 0 107904 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_385
timestamp 1679581782
transform 1 0 108576 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_392
timestamp 1679581782
transform 1 0 109248 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_399
timestamp 1679581782
transform 1 0 109920 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_406
timestamp 1679581782
transform 1 0 110592 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_413
timestamp 1679581782
transform 1 0 111264 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_420
timestamp 1679581782
transform 1 0 111936 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_427
timestamp 1679581782
transform 1 0 112608 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_434
timestamp 1679581782
transform 1 0 113280 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_441
timestamp 1679581782
transform 1 0 113952 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_448
timestamp 1679581782
transform 1 0 114624 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_455
timestamp 1679581782
transform 1 0 115296 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_462
timestamp 1679581782
transform 1 0 115968 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_469
timestamp 1679581782
transform 1 0 116640 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_476
timestamp 1679581782
transform 1 0 117312 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_483
timestamp 1679581782
transform 1 0 117984 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_490
timestamp 1679581782
transform 1 0 118656 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_497
timestamp 1679581782
transform 1 0 119328 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_504
timestamp 1679581782
transform 1 0 120000 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_511
timestamp 1679581782
transform 1 0 120672 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_518
timestamp 1679581782
transform 1 0 121344 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_525
timestamp 1679581782
transform 1 0 122016 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_532
timestamp 1679581782
transform 1 0 122688 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_539
timestamp 1679581782
transform 1 0 123360 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_546
timestamp 1679581782
transform 1 0 124032 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_553
timestamp 1679581782
transform 1 0 124704 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_560
timestamp 1679581782
transform 1 0 125376 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_567
timestamp 1679581782
transform 1 0 126048 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_574
timestamp 1679581782
transform 1 0 126720 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_581
timestamp 1679581782
transform 1 0 127392 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_588
timestamp 1679581782
transform 1 0 128064 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_595
timestamp 1679581782
transform 1 0 128736 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_602
timestamp 1679581782
transform 1 0 129408 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_609
timestamp 1679581782
transform 1 0 130080 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_616
timestamp 1679581782
transform 1 0 130752 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_623
timestamp 1679581782
transform 1 0 131424 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_630
timestamp 1679581782
transform 1 0 132096 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_637
timestamp 1679581782
transform 1 0 132768 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_644
timestamp 1679581782
transform 1 0 133440 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_651
timestamp 1679581782
transform 1 0 134112 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_658
timestamp 1679581782
transform 1 0 134784 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_665
timestamp 1679581782
transform 1 0 135456 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_672
timestamp 1679581782
transform 1 0 136128 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_679
timestamp 1679581782
transform 1 0 136800 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_686
timestamp 1679581782
transform 1 0 137472 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_693
timestamp 1679581782
transform 1 0 138144 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_700
timestamp 1679581782
transform 1 0 138816 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_707
timestamp 1679581782
transform 1 0 139488 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_714
timestamp 1679581782
transform 1 0 140160 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_721
timestamp 1679581782
transform 1 0 140832 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_728
timestamp 1679581782
transform 1 0 141504 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_735
timestamp 1679581782
transform 1 0 142176 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_742
timestamp 1679581782
transform 1 0 142848 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_749
timestamp 1679581782
transform 1 0 143520 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_756
timestamp 1679581782
transform 1 0 144192 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_763
timestamp 1679581782
transform 1 0 144864 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_770
timestamp 1679581782
transform 1 0 145536 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_777
timestamp 1679581782
transform 1 0 146208 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_784
timestamp 1679581782
transform 1 0 146880 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_791
timestamp 1679581782
transform 1 0 147552 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_798
timestamp 1679581782
transform 1 0 148224 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_805
timestamp 1679581782
transform 1 0 148896 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_812
timestamp 1679581782
transform 1 0 149568 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_819
timestamp 1679581782
transform 1 0 150240 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_826
timestamp 1679581782
transform 1 0 150912 0 -1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_833
timestamp 1679581782
transform 1 0 151584 0 -1 86940
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_840
timestamp 1677579658
transform 1 0 152256 0 -1 86940
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_0
timestamp 1679581782
transform 1 0 71616 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_7
timestamp 1679581782
transform 1 0 72288 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_14
timestamp 1679581782
transform 1 0 72960 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_21
timestamp 1679581782
transform 1 0 73632 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_28
timestamp 1679581782
transform 1 0 74304 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_35
timestamp 1679581782
transform 1 0 74976 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_42
timestamp 1679581782
transform 1 0 75648 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_49
timestamp 1679581782
transform 1 0 76320 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_56
timestamp 1679581782
transform 1 0 76992 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_63
timestamp 1679581782
transform 1 0 77664 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_70
timestamp 1679581782
transform 1 0 78336 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_77
timestamp 1679581782
transform 1 0 79008 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_84
timestamp 1679581782
transform 1 0 79680 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_91
timestamp 1679581782
transform 1 0 80352 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_98
timestamp 1679581782
transform 1 0 81024 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_105
timestamp 1679581782
transform 1 0 81696 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_112
timestamp 1679581782
transform 1 0 82368 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_119
timestamp 1679581782
transform 1 0 83040 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_126
timestamp 1679581782
transform 1 0 83712 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_133
timestamp 1679581782
transform 1 0 84384 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_140
timestamp 1679581782
transform 1 0 85056 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_147
timestamp 1679581782
transform 1 0 85728 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_154
timestamp 1679581782
transform 1 0 86400 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_161
timestamp 1679581782
transform 1 0 87072 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_168
timestamp 1679581782
transform 1 0 87744 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_175
timestamp 1679581782
transform 1 0 88416 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_182
timestamp 1679581782
transform 1 0 89088 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_189
timestamp 1679581782
transform 1 0 89760 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_196
timestamp 1679581782
transform 1 0 90432 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_203
timestamp 1679581782
transform 1 0 91104 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_210
timestamp 1679581782
transform 1 0 91776 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_217
timestamp 1679581782
transform 1 0 92448 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_224
timestamp 1679581782
transform 1 0 93120 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_231
timestamp 1679581782
transform 1 0 93792 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_238
timestamp 1679581782
transform 1 0 94464 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_245
timestamp 1679581782
transform 1 0 95136 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_252
timestamp 1679581782
transform 1 0 95808 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_259
timestamp 1679581782
transform 1 0 96480 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_266
timestamp 1679581782
transform 1 0 97152 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_273
timestamp 1679581782
transform 1 0 97824 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_280
timestamp 1679581782
transform 1 0 98496 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_287
timestamp 1679581782
transform 1 0 99168 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_294
timestamp 1679581782
transform 1 0 99840 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_301
timestamp 1679581782
transform 1 0 100512 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_308
timestamp 1679581782
transform 1 0 101184 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_315
timestamp 1679581782
transform 1 0 101856 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_322
timestamp 1679581782
transform 1 0 102528 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_329
timestamp 1679581782
transform 1 0 103200 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_336
timestamp 1679581782
transform 1 0 103872 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_343
timestamp 1679581782
transform 1 0 104544 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_350
timestamp 1679581782
transform 1 0 105216 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_357
timestamp 1679581782
transform 1 0 105888 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_364
timestamp 1679581782
transform 1 0 106560 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_371
timestamp 1679581782
transform 1 0 107232 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_378
timestamp 1679581782
transform 1 0 107904 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_385
timestamp 1679581782
transform 1 0 108576 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_392
timestamp 1679581782
transform 1 0 109248 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_399
timestamp 1679581782
transform 1 0 109920 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_406
timestamp 1679581782
transform 1 0 110592 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_413
timestamp 1679581782
transform 1 0 111264 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_420
timestamp 1679581782
transform 1 0 111936 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_427
timestamp 1679581782
transform 1 0 112608 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_434
timestamp 1679581782
transform 1 0 113280 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_441
timestamp 1679581782
transform 1 0 113952 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_448
timestamp 1679581782
transform 1 0 114624 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_455
timestamp 1679581782
transform 1 0 115296 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_462
timestamp 1679581782
transform 1 0 115968 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_469
timestamp 1679581782
transform 1 0 116640 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_476
timestamp 1679581782
transform 1 0 117312 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_483
timestamp 1679581782
transform 1 0 117984 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_490
timestamp 1679581782
transform 1 0 118656 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_497
timestamp 1679581782
transform 1 0 119328 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_504
timestamp 1679581782
transform 1 0 120000 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_511
timestamp 1679581782
transform 1 0 120672 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_518
timestamp 1679581782
transform 1 0 121344 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_525
timestamp 1679581782
transform 1 0 122016 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_532
timestamp 1679581782
transform 1 0 122688 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_539
timestamp 1679581782
transform 1 0 123360 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_546
timestamp 1679581782
transform 1 0 124032 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_553
timestamp 1679581782
transform 1 0 124704 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_560
timestamp 1679581782
transform 1 0 125376 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_567
timestamp 1679581782
transform 1 0 126048 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_574
timestamp 1679581782
transform 1 0 126720 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_581
timestamp 1679581782
transform 1 0 127392 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_588
timestamp 1679581782
transform 1 0 128064 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_595
timestamp 1679581782
transform 1 0 128736 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_602
timestamp 1679581782
transform 1 0 129408 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_609
timestamp 1679581782
transform 1 0 130080 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_616
timestamp 1679581782
transform 1 0 130752 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_623
timestamp 1679581782
transform 1 0 131424 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_630
timestamp 1679581782
transform 1 0 132096 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_637
timestamp 1679581782
transform 1 0 132768 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_644
timestamp 1679581782
transform 1 0 133440 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_651
timestamp 1679581782
transform 1 0 134112 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_658
timestamp 1679581782
transform 1 0 134784 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_665
timestamp 1679581782
transform 1 0 135456 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_672
timestamp 1679581782
transform 1 0 136128 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_679
timestamp 1679581782
transform 1 0 136800 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_686
timestamp 1679581782
transform 1 0 137472 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_693
timestamp 1679581782
transform 1 0 138144 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_700
timestamp 1679581782
transform 1 0 138816 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_707
timestamp 1679581782
transform 1 0 139488 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_714
timestamp 1679581782
transform 1 0 140160 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_721
timestamp 1679581782
transform 1 0 140832 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_728
timestamp 1679581782
transform 1 0 141504 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_735
timestamp 1679581782
transform 1 0 142176 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_742
timestamp 1679581782
transform 1 0 142848 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_749
timestamp 1679581782
transform 1 0 143520 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_756
timestamp 1679581782
transform 1 0 144192 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_763
timestamp 1679581782
transform 1 0 144864 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_770
timestamp 1679581782
transform 1 0 145536 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_777
timestamp 1679581782
transform 1 0 146208 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_784
timestamp 1679581782
transform 1 0 146880 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_791
timestamp 1679581782
transform 1 0 147552 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_798
timestamp 1679581782
transform 1 0 148224 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_805
timestamp 1679581782
transform 1 0 148896 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_812
timestamp 1679581782
transform 1 0 149568 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_819
timestamp 1679581782
transform 1 0 150240 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_826
timestamp 1679581782
transform 1 0 150912 0 1 86940
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_833
timestamp 1679581782
transform 1 0 151584 0 1 86940
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_840
timestamp 1677579658
transform 1 0 152256 0 1 86940
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_0
timestamp 1679581782
transform 1 0 71616 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_7
timestamp 1679581782
transform 1 0 72288 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_14
timestamp 1679581782
transform 1 0 72960 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_21
timestamp 1679581782
transform 1 0 73632 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_28
timestamp 1679581782
transform 1 0 74304 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_35
timestamp 1679581782
transform 1 0 74976 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_42
timestamp 1679581782
transform 1 0 75648 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_49
timestamp 1679581782
transform 1 0 76320 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_56
timestamp 1679581782
transform 1 0 76992 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_63
timestamp 1679581782
transform 1 0 77664 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_70
timestamp 1679581782
transform 1 0 78336 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_77
timestamp 1679581782
transform 1 0 79008 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_84
timestamp 1679581782
transform 1 0 79680 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_91
timestamp 1679581782
transform 1 0 80352 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_98
timestamp 1679581782
transform 1 0 81024 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_105
timestamp 1679581782
transform 1 0 81696 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_112
timestamp 1679581782
transform 1 0 82368 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_119
timestamp 1679581782
transform 1 0 83040 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_126
timestamp 1679581782
transform 1 0 83712 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_133
timestamp 1679581782
transform 1 0 84384 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_140
timestamp 1679581782
transform 1 0 85056 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_147
timestamp 1679581782
transform 1 0 85728 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_154
timestamp 1679581782
transform 1 0 86400 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_161
timestamp 1679581782
transform 1 0 87072 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_168
timestamp 1679581782
transform 1 0 87744 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_175
timestamp 1679581782
transform 1 0 88416 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_182
timestamp 1679581782
transform 1 0 89088 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_189
timestamp 1679581782
transform 1 0 89760 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_196
timestamp 1679581782
transform 1 0 90432 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_203
timestamp 1679581782
transform 1 0 91104 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_210
timestamp 1679581782
transform 1 0 91776 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_217
timestamp 1679581782
transform 1 0 92448 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_224
timestamp 1679581782
transform 1 0 93120 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_231
timestamp 1679581782
transform 1 0 93792 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_238
timestamp 1679581782
transform 1 0 94464 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_245
timestamp 1679581782
transform 1 0 95136 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_252
timestamp 1679581782
transform 1 0 95808 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_259
timestamp 1679581782
transform 1 0 96480 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_266
timestamp 1679581782
transform 1 0 97152 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_273
timestamp 1679581782
transform 1 0 97824 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_280
timestamp 1679581782
transform 1 0 98496 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_287
timestamp 1679581782
transform 1 0 99168 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_294
timestamp 1679581782
transform 1 0 99840 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_301
timestamp 1679581782
transform 1 0 100512 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_308
timestamp 1679581782
transform 1 0 101184 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_315
timestamp 1679581782
transform 1 0 101856 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_322
timestamp 1679581782
transform 1 0 102528 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_329
timestamp 1679581782
transform 1 0 103200 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_336
timestamp 1679581782
transform 1 0 103872 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_343
timestamp 1679581782
transform 1 0 104544 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_350
timestamp 1679581782
transform 1 0 105216 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_357
timestamp 1679581782
transform 1 0 105888 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_364
timestamp 1679581782
transform 1 0 106560 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_371
timestamp 1679581782
transform 1 0 107232 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_378
timestamp 1679581782
transform 1 0 107904 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_385
timestamp 1679581782
transform 1 0 108576 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_392
timestamp 1679581782
transform 1 0 109248 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_399
timestamp 1679581782
transform 1 0 109920 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_406
timestamp 1679581782
transform 1 0 110592 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_413
timestamp 1679581782
transform 1 0 111264 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_420
timestamp 1679581782
transform 1 0 111936 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_427
timestamp 1679581782
transform 1 0 112608 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_434
timestamp 1679581782
transform 1 0 113280 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_441
timestamp 1679581782
transform 1 0 113952 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_448
timestamp 1679581782
transform 1 0 114624 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_455
timestamp 1679581782
transform 1 0 115296 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_462
timestamp 1679581782
transform 1 0 115968 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_469
timestamp 1679581782
transform 1 0 116640 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_476
timestamp 1679581782
transform 1 0 117312 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_483
timestamp 1679581782
transform 1 0 117984 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_490
timestamp 1679581782
transform 1 0 118656 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_497
timestamp 1679581782
transform 1 0 119328 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_504
timestamp 1679581782
transform 1 0 120000 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_511
timestamp 1679581782
transform 1 0 120672 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_518
timestamp 1679581782
transform 1 0 121344 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_525
timestamp 1679581782
transform 1 0 122016 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_532
timestamp 1679581782
transform 1 0 122688 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_539
timestamp 1679581782
transform 1 0 123360 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_546
timestamp 1679581782
transform 1 0 124032 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_553
timestamp 1679581782
transform 1 0 124704 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_560
timestamp 1679581782
transform 1 0 125376 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_567
timestamp 1679581782
transform 1 0 126048 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_574
timestamp 1679581782
transform 1 0 126720 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_581
timestamp 1679581782
transform 1 0 127392 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_588
timestamp 1679581782
transform 1 0 128064 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_595
timestamp 1679581782
transform 1 0 128736 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_602
timestamp 1679581782
transform 1 0 129408 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_609
timestamp 1679581782
transform 1 0 130080 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_616
timestamp 1679581782
transform 1 0 130752 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_623
timestamp 1679581782
transform 1 0 131424 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_630
timestamp 1679581782
transform 1 0 132096 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_637
timestamp 1679581782
transform 1 0 132768 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_644
timestamp 1679581782
transform 1 0 133440 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_651
timestamp 1679581782
transform 1 0 134112 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_658
timestamp 1679581782
transform 1 0 134784 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_665
timestamp 1679581782
transform 1 0 135456 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_672
timestamp 1679581782
transform 1 0 136128 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_679
timestamp 1679581782
transform 1 0 136800 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_686
timestamp 1679581782
transform 1 0 137472 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_693
timestamp 1679581782
transform 1 0 138144 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_700
timestamp 1679581782
transform 1 0 138816 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_707
timestamp 1679581782
transform 1 0 139488 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_714
timestamp 1679581782
transform 1 0 140160 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_721
timestamp 1679581782
transform 1 0 140832 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_728
timestamp 1679581782
transform 1 0 141504 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_735
timestamp 1679581782
transform 1 0 142176 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_742
timestamp 1679581782
transform 1 0 142848 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_749
timestamp 1679581782
transform 1 0 143520 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_756
timestamp 1679581782
transform 1 0 144192 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_763
timestamp 1679581782
transform 1 0 144864 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_770
timestamp 1679581782
transform 1 0 145536 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_777
timestamp 1679581782
transform 1 0 146208 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_784
timestamp 1679581782
transform 1 0 146880 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_791
timestamp 1679581782
transform 1 0 147552 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_798
timestamp 1679581782
transform 1 0 148224 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_805
timestamp 1679581782
transform 1 0 148896 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_812
timestamp 1679581782
transform 1 0 149568 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_819
timestamp 1679581782
transform 1 0 150240 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_826
timestamp 1679581782
transform 1 0 150912 0 -1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_833
timestamp 1679581782
transform 1 0 151584 0 -1 88452
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_840
timestamp 1677579658
transform 1 0 152256 0 -1 88452
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_0
timestamp 1679581782
transform 1 0 71616 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_7
timestamp 1679581782
transform 1 0 72288 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_14
timestamp 1679581782
transform 1 0 72960 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_21
timestamp 1679581782
transform 1 0 73632 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_28
timestamp 1679581782
transform 1 0 74304 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_35
timestamp 1679581782
transform 1 0 74976 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_42
timestamp 1679581782
transform 1 0 75648 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_49
timestamp 1679581782
transform 1 0 76320 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_56
timestamp 1679581782
transform 1 0 76992 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_63
timestamp 1679581782
transform 1 0 77664 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_70
timestamp 1679581782
transform 1 0 78336 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_77
timestamp 1679581782
transform 1 0 79008 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_84
timestamp 1679581782
transform 1 0 79680 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_91
timestamp 1679581782
transform 1 0 80352 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_98
timestamp 1679581782
transform 1 0 81024 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_105
timestamp 1679581782
transform 1 0 81696 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_112
timestamp 1679581782
transform 1 0 82368 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_119
timestamp 1679581782
transform 1 0 83040 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_126
timestamp 1679581782
transform 1 0 83712 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_133
timestamp 1679581782
transform 1 0 84384 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_140
timestamp 1679581782
transform 1 0 85056 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_147
timestamp 1679581782
transform 1 0 85728 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_154
timestamp 1679581782
transform 1 0 86400 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_161
timestamp 1679581782
transform 1 0 87072 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_168
timestamp 1679581782
transform 1 0 87744 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_175
timestamp 1679581782
transform 1 0 88416 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_182
timestamp 1679581782
transform 1 0 89088 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_189
timestamp 1679581782
transform 1 0 89760 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_196
timestamp 1679581782
transform 1 0 90432 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_203
timestamp 1679581782
transform 1 0 91104 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_210
timestamp 1679581782
transform 1 0 91776 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_217
timestamp 1679581782
transform 1 0 92448 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_224
timestamp 1679581782
transform 1 0 93120 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_231
timestamp 1679581782
transform 1 0 93792 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_238
timestamp 1679581782
transform 1 0 94464 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_245
timestamp 1679581782
transform 1 0 95136 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_252
timestamp 1679581782
transform 1 0 95808 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_259
timestamp 1679581782
transform 1 0 96480 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_266
timestamp 1679581782
transform 1 0 97152 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_273
timestamp 1679581782
transform 1 0 97824 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_280
timestamp 1679581782
transform 1 0 98496 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_287
timestamp 1679581782
transform 1 0 99168 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_294
timestamp 1679581782
transform 1 0 99840 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_301
timestamp 1679581782
transform 1 0 100512 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_308
timestamp 1679581782
transform 1 0 101184 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_315
timestamp 1679581782
transform 1 0 101856 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_322
timestamp 1679581782
transform 1 0 102528 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_329
timestamp 1679581782
transform 1 0 103200 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_336
timestamp 1679581782
transform 1 0 103872 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_343
timestamp 1679581782
transform 1 0 104544 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_350
timestamp 1679581782
transform 1 0 105216 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_357
timestamp 1679581782
transform 1 0 105888 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_364
timestamp 1679581782
transform 1 0 106560 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_371
timestamp 1679581782
transform 1 0 107232 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_378
timestamp 1679581782
transform 1 0 107904 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_385
timestamp 1679581782
transform 1 0 108576 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_392
timestamp 1679581782
transform 1 0 109248 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_399
timestamp 1679581782
transform 1 0 109920 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_406
timestamp 1679581782
transform 1 0 110592 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_413
timestamp 1679581782
transform 1 0 111264 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_420
timestamp 1679581782
transform 1 0 111936 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_427
timestamp 1679581782
transform 1 0 112608 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_434
timestamp 1679581782
transform 1 0 113280 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_441
timestamp 1679581782
transform 1 0 113952 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_448
timestamp 1679581782
transform 1 0 114624 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_455
timestamp 1679581782
transform 1 0 115296 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_462
timestamp 1679581782
transform 1 0 115968 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_469
timestamp 1679581782
transform 1 0 116640 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_476
timestamp 1679581782
transform 1 0 117312 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_483
timestamp 1679581782
transform 1 0 117984 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_490
timestamp 1679581782
transform 1 0 118656 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_497
timestamp 1679581782
transform 1 0 119328 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_504
timestamp 1679581782
transform 1 0 120000 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_511
timestamp 1679581782
transform 1 0 120672 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_518
timestamp 1679581782
transform 1 0 121344 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_525
timestamp 1679581782
transform 1 0 122016 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_532
timestamp 1679581782
transform 1 0 122688 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_539
timestamp 1679581782
transform 1 0 123360 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_546
timestamp 1679581782
transform 1 0 124032 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_553
timestamp 1679581782
transform 1 0 124704 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_560
timestamp 1679581782
transform 1 0 125376 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_567
timestamp 1679581782
transform 1 0 126048 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_574
timestamp 1679581782
transform 1 0 126720 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_581
timestamp 1679581782
transform 1 0 127392 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_588
timestamp 1679581782
transform 1 0 128064 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_595
timestamp 1679581782
transform 1 0 128736 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_602
timestamp 1679581782
transform 1 0 129408 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_609
timestamp 1679581782
transform 1 0 130080 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_616
timestamp 1679581782
transform 1 0 130752 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_623
timestamp 1679581782
transform 1 0 131424 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_630
timestamp 1679581782
transform 1 0 132096 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_637
timestamp 1679581782
transform 1 0 132768 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_644
timestamp 1679581782
transform 1 0 133440 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_651
timestamp 1679581782
transform 1 0 134112 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_658
timestamp 1679581782
transform 1 0 134784 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_665
timestamp 1679581782
transform 1 0 135456 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_672
timestamp 1679581782
transform 1 0 136128 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_679
timestamp 1679581782
transform 1 0 136800 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_686
timestamp 1679581782
transform 1 0 137472 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_693
timestamp 1679581782
transform 1 0 138144 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_700
timestamp 1679581782
transform 1 0 138816 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_707
timestamp 1679581782
transform 1 0 139488 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_714
timestamp 1679581782
transform 1 0 140160 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_721
timestamp 1679581782
transform 1 0 140832 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_728
timestamp 1679581782
transform 1 0 141504 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_735
timestamp 1679581782
transform 1 0 142176 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_742
timestamp 1679581782
transform 1 0 142848 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_749
timestamp 1679581782
transform 1 0 143520 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_756
timestamp 1679581782
transform 1 0 144192 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_763
timestamp 1679581782
transform 1 0 144864 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_770
timestamp 1679581782
transform 1 0 145536 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_777
timestamp 1679581782
transform 1 0 146208 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_784
timestamp 1679581782
transform 1 0 146880 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_791
timestamp 1679581782
transform 1 0 147552 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_798
timestamp 1679581782
transform 1 0 148224 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_805
timestamp 1679581782
transform 1 0 148896 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_812
timestamp 1679581782
transform 1 0 149568 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_819
timestamp 1679581782
transform 1 0 150240 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_826
timestamp 1679581782
transform 1 0 150912 0 1 88452
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_833
timestamp 1679581782
transform 1 0 151584 0 1 88452
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_840
timestamp 1677579658
transform 1 0 152256 0 1 88452
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_0
timestamp 1679581782
transform 1 0 71616 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_7
timestamp 1679581782
transform 1 0 72288 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_14
timestamp 1679581782
transform 1 0 72960 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_21
timestamp 1679581782
transform 1 0 73632 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_28
timestamp 1679581782
transform 1 0 74304 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_35
timestamp 1679581782
transform 1 0 74976 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_42
timestamp 1679581782
transform 1 0 75648 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_49
timestamp 1679581782
transform 1 0 76320 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_56
timestamp 1679581782
transform 1 0 76992 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_63
timestamp 1679581782
transform 1 0 77664 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_70
timestamp 1679581782
transform 1 0 78336 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_77
timestamp 1679581782
transform 1 0 79008 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_84
timestamp 1679581782
transform 1 0 79680 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_91
timestamp 1679581782
transform 1 0 80352 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_98
timestamp 1679581782
transform 1 0 81024 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_105
timestamp 1679581782
transform 1 0 81696 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_112
timestamp 1679581782
transform 1 0 82368 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_119
timestamp 1679581782
transform 1 0 83040 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_126
timestamp 1679581782
transform 1 0 83712 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_133
timestamp 1679581782
transform 1 0 84384 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_140
timestamp 1679581782
transform 1 0 85056 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_147
timestamp 1679581782
transform 1 0 85728 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_154
timestamp 1679581782
transform 1 0 86400 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_161
timestamp 1679581782
transform 1 0 87072 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_168
timestamp 1679581782
transform 1 0 87744 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_175
timestamp 1679581782
transform 1 0 88416 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_182
timestamp 1679581782
transform 1 0 89088 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_189
timestamp 1679581782
transform 1 0 89760 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_196
timestamp 1679581782
transform 1 0 90432 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_203
timestamp 1679581782
transform 1 0 91104 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_210
timestamp 1679581782
transform 1 0 91776 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_217
timestamp 1679581782
transform 1 0 92448 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_224
timestamp 1679581782
transform 1 0 93120 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_231
timestamp 1679581782
transform 1 0 93792 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_238
timestamp 1679581782
transform 1 0 94464 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_245
timestamp 1679581782
transform 1 0 95136 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_252
timestamp 1679581782
transform 1 0 95808 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_259
timestamp 1679581782
transform 1 0 96480 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_266
timestamp 1679581782
transform 1 0 97152 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_273
timestamp 1679581782
transform 1 0 97824 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_280
timestamp 1679581782
transform 1 0 98496 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_287
timestamp 1679581782
transform 1 0 99168 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_294
timestamp 1679581782
transform 1 0 99840 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_301
timestamp 1679581782
transform 1 0 100512 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_308
timestamp 1679581782
transform 1 0 101184 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_315
timestamp 1679581782
transform 1 0 101856 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_322
timestamp 1679581782
transform 1 0 102528 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_329
timestamp 1679581782
transform 1 0 103200 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_336
timestamp 1679581782
transform 1 0 103872 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_343
timestamp 1679581782
transform 1 0 104544 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_350
timestamp 1679581782
transform 1 0 105216 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_357
timestamp 1679581782
transform 1 0 105888 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_364
timestamp 1679581782
transform 1 0 106560 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_371
timestamp 1679581782
transform 1 0 107232 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_378
timestamp 1679581782
transform 1 0 107904 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_385
timestamp 1679581782
transform 1 0 108576 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_392
timestamp 1679581782
transform 1 0 109248 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_399
timestamp 1679581782
transform 1 0 109920 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_406
timestamp 1679581782
transform 1 0 110592 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_413
timestamp 1679581782
transform 1 0 111264 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_420
timestamp 1679581782
transform 1 0 111936 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_427
timestamp 1679581782
transform 1 0 112608 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_434
timestamp 1679581782
transform 1 0 113280 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_441
timestamp 1679581782
transform 1 0 113952 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_448
timestamp 1679581782
transform 1 0 114624 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_455
timestamp 1679581782
transform 1 0 115296 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_462
timestamp 1679581782
transform 1 0 115968 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_469
timestamp 1679581782
transform 1 0 116640 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_476
timestamp 1679581782
transform 1 0 117312 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_483
timestamp 1679581782
transform 1 0 117984 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_490
timestamp 1679581782
transform 1 0 118656 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_497
timestamp 1679581782
transform 1 0 119328 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_504
timestamp 1679581782
transform 1 0 120000 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_511
timestamp 1679581782
transform 1 0 120672 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_518
timestamp 1679581782
transform 1 0 121344 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_525
timestamp 1679581782
transform 1 0 122016 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_532
timestamp 1679581782
transform 1 0 122688 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_539
timestamp 1679581782
transform 1 0 123360 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_546
timestamp 1679581782
transform 1 0 124032 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_553
timestamp 1679581782
transform 1 0 124704 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_560
timestamp 1679581782
transform 1 0 125376 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_567
timestamp 1679581782
transform 1 0 126048 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_574
timestamp 1679581782
transform 1 0 126720 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_581
timestamp 1679581782
transform 1 0 127392 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_588
timestamp 1679581782
transform 1 0 128064 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_595
timestamp 1679581782
transform 1 0 128736 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_602
timestamp 1679581782
transform 1 0 129408 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_609
timestamp 1679581782
transform 1 0 130080 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_616
timestamp 1679581782
transform 1 0 130752 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_623
timestamp 1679581782
transform 1 0 131424 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_630
timestamp 1679581782
transform 1 0 132096 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_637
timestamp 1679581782
transform 1 0 132768 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_644
timestamp 1679581782
transform 1 0 133440 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_651
timestamp 1679581782
transform 1 0 134112 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_658
timestamp 1679581782
transform 1 0 134784 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_665
timestamp 1679581782
transform 1 0 135456 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_672
timestamp 1679581782
transform 1 0 136128 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_679
timestamp 1679581782
transform 1 0 136800 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_686
timestamp 1679581782
transform 1 0 137472 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_693
timestamp 1679581782
transform 1 0 138144 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_700
timestamp 1679581782
transform 1 0 138816 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_707
timestamp 1679581782
transform 1 0 139488 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_714
timestamp 1679581782
transform 1 0 140160 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_721
timestamp 1679581782
transform 1 0 140832 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_728
timestamp 1679581782
transform 1 0 141504 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_735
timestamp 1679581782
transform 1 0 142176 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_742
timestamp 1679581782
transform 1 0 142848 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_749
timestamp 1679581782
transform 1 0 143520 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_756
timestamp 1679581782
transform 1 0 144192 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_763
timestamp 1679581782
transform 1 0 144864 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_770
timestamp 1679581782
transform 1 0 145536 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_777
timestamp 1679581782
transform 1 0 146208 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_784
timestamp 1679581782
transform 1 0 146880 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_791
timestamp 1679581782
transform 1 0 147552 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_798
timestamp 1679581782
transform 1 0 148224 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_805
timestamp 1679581782
transform 1 0 148896 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_812
timestamp 1679581782
transform 1 0 149568 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_819
timestamp 1679581782
transform 1 0 150240 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_826
timestamp 1679581782
transform 1 0 150912 0 -1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_833
timestamp 1679581782
transform 1 0 151584 0 -1 89964
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_840
timestamp 1677579658
transform 1 0 152256 0 -1 89964
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_0
timestamp 1679581782
transform 1 0 71616 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_7
timestamp 1679581782
transform 1 0 72288 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_14
timestamp 1679581782
transform 1 0 72960 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_21
timestamp 1679581782
transform 1 0 73632 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_28
timestamp 1679581782
transform 1 0 74304 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_35
timestamp 1679581782
transform 1 0 74976 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_42
timestamp 1679581782
transform 1 0 75648 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_49
timestamp 1679581782
transform 1 0 76320 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_56
timestamp 1679581782
transform 1 0 76992 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_63
timestamp 1679581782
transform 1 0 77664 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_70
timestamp 1679581782
transform 1 0 78336 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_77
timestamp 1679581782
transform 1 0 79008 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_84
timestamp 1679581782
transform 1 0 79680 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_91
timestamp 1679581782
transform 1 0 80352 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_98
timestamp 1679581782
transform 1 0 81024 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_105
timestamp 1679581782
transform 1 0 81696 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_112
timestamp 1679581782
transform 1 0 82368 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_119
timestamp 1679581782
transform 1 0 83040 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_126
timestamp 1679581782
transform 1 0 83712 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_133
timestamp 1679581782
transform 1 0 84384 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_140
timestamp 1679581782
transform 1 0 85056 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_147
timestamp 1679581782
transform 1 0 85728 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_154
timestamp 1679581782
transform 1 0 86400 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_161
timestamp 1679581782
transform 1 0 87072 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_168
timestamp 1679581782
transform 1 0 87744 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_175
timestamp 1679581782
transform 1 0 88416 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_182
timestamp 1679581782
transform 1 0 89088 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_189
timestamp 1679581782
transform 1 0 89760 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_196
timestamp 1679581782
transform 1 0 90432 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_203
timestamp 1679581782
transform 1 0 91104 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_210
timestamp 1679581782
transform 1 0 91776 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_217
timestamp 1679581782
transform 1 0 92448 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_224
timestamp 1679581782
transform 1 0 93120 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_231
timestamp 1679581782
transform 1 0 93792 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_238
timestamp 1679581782
transform 1 0 94464 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_245
timestamp 1679581782
transform 1 0 95136 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_252
timestamp 1679581782
transform 1 0 95808 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_259
timestamp 1679581782
transform 1 0 96480 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_266
timestamp 1679581782
transform 1 0 97152 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_273
timestamp 1679581782
transform 1 0 97824 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_280
timestamp 1679581782
transform 1 0 98496 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_287
timestamp 1679581782
transform 1 0 99168 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_294
timestamp 1679581782
transform 1 0 99840 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_301
timestamp 1679581782
transform 1 0 100512 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_308
timestamp 1679581782
transform 1 0 101184 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_315
timestamp 1679581782
transform 1 0 101856 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_322
timestamp 1679581782
transform 1 0 102528 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_329
timestamp 1679581782
transform 1 0 103200 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_336
timestamp 1679581782
transform 1 0 103872 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_343
timestamp 1679581782
transform 1 0 104544 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_350
timestamp 1679581782
transform 1 0 105216 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_357
timestamp 1679581782
transform 1 0 105888 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_364
timestamp 1679581782
transform 1 0 106560 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_371
timestamp 1679581782
transform 1 0 107232 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_378
timestamp 1679581782
transform 1 0 107904 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_385
timestamp 1679581782
transform 1 0 108576 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_392
timestamp 1679581782
transform 1 0 109248 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_399
timestamp 1679581782
transform 1 0 109920 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_406
timestamp 1679581782
transform 1 0 110592 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_413
timestamp 1679581782
transform 1 0 111264 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_420
timestamp 1679581782
transform 1 0 111936 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_427
timestamp 1679581782
transform 1 0 112608 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_434
timestamp 1679581782
transform 1 0 113280 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_441
timestamp 1679581782
transform 1 0 113952 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_448
timestamp 1679581782
transform 1 0 114624 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_455
timestamp 1679581782
transform 1 0 115296 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_462
timestamp 1679581782
transform 1 0 115968 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_469
timestamp 1679581782
transform 1 0 116640 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_476
timestamp 1679581782
transform 1 0 117312 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_483
timestamp 1679581782
transform 1 0 117984 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_490
timestamp 1679581782
transform 1 0 118656 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_497
timestamp 1679581782
transform 1 0 119328 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_504
timestamp 1679581782
transform 1 0 120000 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_511
timestamp 1679581782
transform 1 0 120672 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_518
timestamp 1679581782
transform 1 0 121344 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_525
timestamp 1679581782
transform 1 0 122016 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_532
timestamp 1679581782
transform 1 0 122688 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_539
timestamp 1679581782
transform 1 0 123360 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_546
timestamp 1679581782
transform 1 0 124032 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_553
timestamp 1679581782
transform 1 0 124704 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_560
timestamp 1679581782
transform 1 0 125376 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_567
timestamp 1679581782
transform 1 0 126048 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_574
timestamp 1679581782
transform 1 0 126720 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_581
timestamp 1679581782
transform 1 0 127392 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_588
timestamp 1679581782
transform 1 0 128064 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_595
timestamp 1679581782
transform 1 0 128736 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_602
timestamp 1679581782
transform 1 0 129408 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_609
timestamp 1679581782
transform 1 0 130080 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_616
timestamp 1679581782
transform 1 0 130752 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_623
timestamp 1679581782
transform 1 0 131424 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_630
timestamp 1679581782
transform 1 0 132096 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_637
timestamp 1679581782
transform 1 0 132768 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_644
timestamp 1679581782
transform 1 0 133440 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_651
timestamp 1679581782
transform 1 0 134112 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_658
timestamp 1679581782
transform 1 0 134784 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_665
timestamp 1679581782
transform 1 0 135456 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_672
timestamp 1679581782
transform 1 0 136128 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_679
timestamp 1679581782
transform 1 0 136800 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_686
timestamp 1679581782
transform 1 0 137472 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_693
timestamp 1679581782
transform 1 0 138144 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_700
timestamp 1679581782
transform 1 0 138816 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_707
timestamp 1679581782
transform 1 0 139488 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_714
timestamp 1679581782
transform 1 0 140160 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_721
timestamp 1679581782
transform 1 0 140832 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_728
timestamp 1679581782
transform 1 0 141504 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_735
timestamp 1679581782
transform 1 0 142176 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_742
timestamp 1679581782
transform 1 0 142848 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_749
timestamp 1679581782
transform 1 0 143520 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_756
timestamp 1679581782
transform 1 0 144192 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_763
timestamp 1679581782
transform 1 0 144864 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_770
timestamp 1679581782
transform 1 0 145536 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_777
timestamp 1679581782
transform 1 0 146208 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_784
timestamp 1679581782
transform 1 0 146880 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_791
timestamp 1679581782
transform 1 0 147552 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_798
timestamp 1679581782
transform 1 0 148224 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_805
timestamp 1679581782
transform 1 0 148896 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_812
timestamp 1679581782
transform 1 0 149568 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_819
timestamp 1679581782
transform 1 0 150240 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_826
timestamp 1679581782
transform 1 0 150912 0 1 89964
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_833
timestamp 1679581782
transform 1 0 151584 0 1 89964
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_840
timestamp 1677579658
transform 1 0 152256 0 1 89964
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_0
timestamp 1679581782
transform 1 0 71616 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_7
timestamp 1679581782
transform 1 0 72288 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_14
timestamp 1679581782
transform 1 0 72960 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_21
timestamp 1679581782
transform 1 0 73632 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_28
timestamp 1679581782
transform 1 0 74304 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_35
timestamp 1679581782
transform 1 0 74976 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_42
timestamp 1679581782
transform 1 0 75648 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_49
timestamp 1679581782
transform 1 0 76320 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_56
timestamp 1679581782
transform 1 0 76992 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_63
timestamp 1679581782
transform 1 0 77664 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_70
timestamp 1679581782
transform 1 0 78336 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_77
timestamp 1679581782
transform 1 0 79008 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_84
timestamp 1679581782
transform 1 0 79680 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_91
timestamp 1679581782
transform 1 0 80352 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_98
timestamp 1679581782
transform 1 0 81024 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_105
timestamp 1679581782
transform 1 0 81696 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_112
timestamp 1679581782
transform 1 0 82368 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_119
timestamp 1679581782
transform 1 0 83040 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_126
timestamp 1679581782
transform 1 0 83712 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_133
timestamp 1679581782
transform 1 0 84384 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_140
timestamp 1679581782
transform 1 0 85056 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_147
timestamp 1679581782
transform 1 0 85728 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_154
timestamp 1679581782
transform 1 0 86400 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_161
timestamp 1679581782
transform 1 0 87072 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_168
timestamp 1679581782
transform 1 0 87744 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_175
timestamp 1679581782
transform 1 0 88416 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_182
timestamp 1679581782
transform 1 0 89088 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_189
timestamp 1679581782
transform 1 0 89760 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_196
timestamp 1679581782
transform 1 0 90432 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_203
timestamp 1679581782
transform 1 0 91104 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_210
timestamp 1679581782
transform 1 0 91776 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_217
timestamp 1679581782
transform 1 0 92448 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_224
timestamp 1679581782
transform 1 0 93120 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_231
timestamp 1679581782
transform 1 0 93792 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_238
timestamp 1679581782
transform 1 0 94464 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_245
timestamp 1679581782
transform 1 0 95136 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_252
timestamp 1679581782
transform 1 0 95808 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_259
timestamp 1679581782
transform 1 0 96480 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_266
timestamp 1679581782
transform 1 0 97152 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_273
timestamp 1679581782
transform 1 0 97824 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_280
timestamp 1679581782
transform 1 0 98496 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_287
timestamp 1679581782
transform 1 0 99168 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_294
timestamp 1679581782
transform 1 0 99840 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_301
timestamp 1679581782
transform 1 0 100512 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_308
timestamp 1679581782
transform 1 0 101184 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_315
timestamp 1679581782
transform 1 0 101856 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_322
timestamp 1679581782
transform 1 0 102528 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_329
timestamp 1679581782
transform 1 0 103200 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_336
timestamp 1679581782
transform 1 0 103872 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_343
timestamp 1679581782
transform 1 0 104544 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_350
timestamp 1679581782
transform 1 0 105216 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_357
timestamp 1679581782
transform 1 0 105888 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_364
timestamp 1679581782
transform 1 0 106560 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_371
timestamp 1679581782
transform 1 0 107232 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_378
timestamp 1679581782
transform 1 0 107904 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_385
timestamp 1679581782
transform 1 0 108576 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_392
timestamp 1679581782
transform 1 0 109248 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_399
timestamp 1679581782
transform 1 0 109920 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_406
timestamp 1679581782
transform 1 0 110592 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_413
timestamp 1679581782
transform 1 0 111264 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_420
timestamp 1679581782
transform 1 0 111936 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_427
timestamp 1679581782
transform 1 0 112608 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_434
timestamp 1679581782
transform 1 0 113280 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_441
timestamp 1679581782
transform 1 0 113952 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_448
timestamp 1679581782
transform 1 0 114624 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_455
timestamp 1679581782
transform 1 0 115296 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_462
timestamp 1679581782
transform 1 0 115968 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_469
timestamp 1679581782
transform 1 0 116640 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_476
timestamp 1679581782
transform 1 0 117312 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_483
timestamp 1679581782
transform 1 0 117984 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_490
timestamp 1679581782
transform 1 0 118656 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_497
timestamp 1679581782
transform 1 0 119328 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_504
timestamp 1679581782
transform 1 0 120000 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_511
timestamp 1679581782
transform 1 0 120672 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_518
timestamp 1679581782
transform 1 0 121344 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_525
timestamp 1679581782
transform 1 0 122016 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_532
timestamp 1679581782
transform 1 0 122688 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_539
timestamp 1679581782
transform 1 0 123360 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_546
timestamp 1679581782
transform 1 0 124032 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_553
timestamp 1679581782
transform 1 0 124704 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_560
timestamp 1679581782
transform 1 0 125376 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_567
timestamp 1679581782
transform 1 0 126048 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_574
timestamp 1679581782
transform 1 0 126720 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_581
timestamp 1679581782
transform 1 0 127392 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_588
timestamp 1679581782
transform 1 0 128064 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_595
timestamp 1679581782
transform 1 0 128736 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_602
timestamp 1679581782
transform 1 0 129408 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_609
timestamp 1679581782
transform 1 0 130080 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_616
timestamp 1679581782
transform 1 0 130752 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_623
timestamp 1679581782
transform 1 0 131424 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_630
timestamp 1679581782
transform 1 0 132096 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_637
timestamp 1679581782
transform 1 0 132768 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_644
timestamp 1679581782
transform 1 0 133440 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_651
timestamp 1679581782
transform 1 0 134112 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_658
timestamp 1679581782
transform 1 0 134784 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_665
timestamp 1679581782
transform 1 0 135456 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_672
timestamp 1679581782
transform 1 0 136128 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_679
timestamp 1679581782
transform 1 0 136800 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_686
timestamp 1679581782
transform 1 0 137472 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_693
timestamp 1679581782
transform 1 0 138144 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_700
timestamp 1679581782
transform 1 0 138816 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_707
timestamp 1679581782
transform 1 0 139488 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_714
timestamp 1679581782
transform 1 0 140160 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_721
timestamp 1679581782
transform 1 0 140832 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_728
timestamp 1679581782
transform 1 0 141504 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_735
timestamp 1679581782
transform 1 0 142176 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_742
timestamp 1679581782
transform 1 0 142848 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_749
timestamp 1679581782
transform 1 0 143520 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_756
timestamp 1679581782
transform 1 0 144192 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_763
timestamp 1679581782
transform 1 0 144864 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_770
timestamp 1679581782
transform 1 0 145536 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_777
timestamp 1679581782
transform 1 0 146208 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_784
timestamp 1679581782
transform 1 0 146880 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_791
timestamp 1679581782
transform 1 0 147552 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_798
timestamp 1679581782
transform 1 0 148224 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_805
timestamp 1679581782
transform 1 0 148896 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_812
timestamp 1679581782
transform 1 0 149568 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_819
timestamp 1679581782
transform 1 0 150240 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_826
timestamp 1679581782
transform 1 0 150912 0 -1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_833
timestamp 1679581782
transform 1 0 151584 0 -1 91476
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_840
timestamp 1677579658
transform 1 0 152256 0 -1 91476
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_0
timestamp 1679581782
transform 1 0 71616 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_7
timestamp 1679581782
transform 1 0 72288 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_14
timestamp 1679581782
transform 1 0 72960 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_21
timestamp 1679581782
transform 1 0 73632 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_28
timestamp 1679581782
transform 1 0 74304 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_35
timestamp 1679581782
transform 1 0 74976 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_42
timestamp 1679581782
transform 1 0 75648 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_49
timestamp 1679581782
transform 1 0 76320 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_56
timestamp 1679581782
transform 1 0 76992 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_63
timestamp 1679581782
transform 1 0 77664 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_70
timestamp 1679581782
transform 1 0 78336 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_77
timestamp 1679581782
transform 1 0 79008 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_84
timestamp 1679581782
transform 1 0 79680 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_91
timestamp 1679581782
transform 1 0 80352 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_98
timestamp 1679581782
transform 1 0 81024 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_105
timestamp 1679581782
transform 1 0 81696 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_112
timestamp 1679581782
transform 1 0 82368 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_119
timestamp 1679581782
transform 1 0 83040 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_126
timestamp 1679581782
transform 1 0 83712 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_133
timestamp 1679581782
transform 1 0 84384 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_140
timestamp 1679581782
transform 1 0 85056 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_147
timestamp 1679581782
transform 1 0 85728 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_154
timestamp 1679581782
transform 1 0 86400 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_161
timestamp 1679581782
transform 1 0 87072 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_168
timestamp 1679581782
transform 1 0 87744 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_175
timestamp 1679581782
transform 1 0 88416 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_182
timestamp 1679581782
transform 1 0 89088 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_189
timestamp 1679581782
transform 1 0 89760 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_196
timestamp 1679581782
transform 1 0 90432 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_203
timestamp 1679581782
transform 1 0 91104 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_210
timestamp 1679581782
transform 1 0 91776 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_217
timestamp 1679581782
transform 1 0 92448 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_224
timestamp 1679581782
transform 1 0 93120 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_231
timestamp 1679581782
transform 1 0 93792 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_238
timestamp 1679581782
transform 1 0 94464 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_245
timestamp 1679581782
transform 1 0 95136 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_252
timestamp 1679581782
transform 1 0 95808 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_259
timestamp 1679581782
transform 1 0 96480 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_266
timestamp 1679581782
transform 1 0 97152 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_273
timestamp 1679581782
transform 1 0 97824 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_280
timestamp 1679581782
transform 1 0 98496 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_287
timestamp 1679581782
transform 1 0 99168 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_294
timestamp 1679581782
transform 1 0 99840 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_301
timestamp 1679581782
transform 1 0 100512 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_308
timestamp 1679581782
transform 1 0 101184 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_315
timestamp 1679581782
transform 1 0 101856 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_322
timestamp 1679581782
transform 1 0 102528 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_329
timestamp 1679581782
transform 1 0 103200 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_336
timestamp 1679581782
transform 1 0 103872 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_343
timestamp 1679581782
transform 1 0 104544 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_350
timestamp 1679581782
transform 1 0 105216 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_357
timestamp 1679581782
transform 1 0 105888 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_364
timestamp 1679581782
transform 1 0 106560 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_371
timestamp 1679581782
transform 1 0 107232 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_378
timestamp 1679581782
transform 1 0 107904 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_385
timestamp 1679581782
transform 1 0 108576 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_392
timestamp 1679581782
transform 1 0 109248 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_399
timestamp 1679581782
transform 1 0 109920 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_406
timestamp 1679581782
transform 1 0 110592 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_413
timestamp 1679581782
transform 1 0 111264 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_420
timestamp 1679581782
transform 1 0 111936 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_427
timestamp 1679581782
transform 1 0 112608 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_434
timestamp 1679581782
transform 1 0 113280 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_441
timestamp 1679581782
transform 1 0 113952 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_448
timestamp 1679581782
transform 1 0 114624 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_455
timestamp 1679581782
transform 1 0 115296 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_462
timestamp 1679581782
transform 1 0 115968 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_469
timestamp 1679581782
transform 1 0 116640 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_476
timestamp 1679581782
transform 1 0 117312 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_483
timestamp 1679581782
transform 1 0 117984 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_490
timestamp 1679581782
transform 1 0 118656 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_497
timestamp 1679581782
transform 1 0 119328 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_504
timestamp 1679581782
transform 1 0 120000 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_511
timestamp 1679581782
transform 1 0 120672 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_518
timestamp 1679581782
transform 1 0 121344 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_525
timestamp 1679581782
transform 1 0 122016 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_532
timestamp 1679581782
transform 1 0 122688 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_539
timestamp 1679581782
transform 1 0 123360 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_546
timestamp 1679581782
transform 1 0 124032 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_553
timestamp 1679581782
transform 1 0 124704 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_560
timestamp 1679581782
transform 1 0 125376 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_567
timestamp 1679581782
transform 1 0 126048 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_574
timestamp 1679581782
transform 1 0 126720 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_581
timestamp 1679581782
transform 1 0 127392 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_588
timestamp 1679581782
transform 1 0 128064 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_595
timestamp 1679581782
transform 1 0 128736 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_602
timestamp 1679581782
transform 1 0 129408 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_609
timestamp 1679581782
transform 1 0 130080 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_616
timestamp 1679581782
transform 1 0 130752 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_623
timestamp 1679581782
transform 1 0 131424 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_630
timestamp 1679581782
transform 1 0 132096 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_637
timestamp 1679581782
transform 1 0 132768 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_644
timestamp 1679581782
transform 1 0 133440 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_651
timestamp 1679581782
transform 1 0 134112 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_658
timestamp 1679581782
transform 1 0 134784 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_665
timestamp 1679581782
transform 1 0 135456 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_672
timestamp 1679581782
transform 1 0 136128 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_679
timestamp 1679581782
transform 1 0 136800 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_686
timestamp 1679581782
transform 1 0 137472 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_693
timestamp 1679581782
transform 1 0 138144 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_700
timestamp 1679581782
transform 1 0 138816 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_707
timestamp 1679581782
transform 1 0 139488 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_714
timestamp 1679581782
transform 1 0 140160 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_721
timestamp 1679581782
transform 1 0 140832 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_728
timestamp 1679581782
transform 1 0 141504 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_735
timestamp 1679581782
transform 1 0 142176 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_742
timestamp 1679581782
transform 1 0 142848 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_749
timestamp 1679581782
transform 1 0 143520 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_756
timestamp 1679581782
transform 1 0 144192 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_763
timestamp 1679581782
transform 1 0 144864 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_770
timestamp 1679581782
transform 1 0 145536 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_777
timestamp 1679581782
transform 1 0 146208 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_784
timestamp 1679581782
transform 1 0 146880 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_791
timestamp 1679581782
transform 1 0 147552 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_798
timestamp 1679581782
transform 1 0 148224 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_805
timestamp 1679581782
transform 1 0 148896 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_812
timestamp 1679581782
transform 1 0 149568 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_819
timestamp 1679581782
transform 1 0 150240 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_826
timestamp 1679581782
transform 1 0 150912 0 1 91476
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_833
timestamp 1679581782
transform 1 0 151584 0 1 91476
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_840
timestamp 1677579658
transform 1 0 152256 0 1 91476
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 71616 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679581782
transform 1 0 72288 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679581782
transform 1 0 72960 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679581782
transform 1 0 73632 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_28
timestamp 1679581782
transform 1 0 74304 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_35
timestamp 1679581782
transform 1 0 74976 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_42
timestamp 1679581782
transform 1 0 75648 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_49
timestamp 1679581782
transform 1 0 76320 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_56
timestamp 1679581782
transform 1 0 76992 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_63
timestamp 1679581782
transform 1 0 77664 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_70
timestamp 1679581782
transform 1 0 78336 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_77
timestamp 1679581782
transform 1 0 79008 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_84
timestamp 1679581782
transform 1 0 79680 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_91
timestamp 1679581782
transform 1 0 80352 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_98
timestamp 1679581782
transform 1 0 81024 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_105
timestamp 1679581782
transform 1 0 81696 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_112
timestamp 1679581782
transform 1 0 82368 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_119
timestamp 1679581782
transform 1 0 83040 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_126
timestamp 1679581782
transform 1 0 83712 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_133
timestamp 1679581782
transform 1 0 84384 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_140
timestamp 1679581782
transform 1 0 85056 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_147
timestamp 1679581782
transform 1 0 85728 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_154
timestamp 1679581782
transform 1 0 86400 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_161
timestamp 1679581782
transform 1 0 87072 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_168
timestamp 1679581782
transform 1 0 87744 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_175
timestamp 1679581782
transform 1 0 88416 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_182
timestamp 1679581782
transform 1 0 89088 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_189
timestamp 1679581782
transform 1 0 89760 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_196
timestamp 1679581782
transform 1 0 90432 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_203
timestamp 1679581782
transform 1 0 91104 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_210
timestamp 1679581782
transform 1 0 91776 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_217
timestamp 1679581782
transform 1 0 92448 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_224
timestamp 1679581782
transform 1 0 93120 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_231
timestamp 1679581782
transform 1 0 93792 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_238
timestamp 1679581782
transform 1 0 94464 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_245
timestamp 1679581782
transform 1 0 95136 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_252
timestamp 1679581782
transform 1 0 95808 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_259
timestamp 1679581782
transform 1 0 96480 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_266
timestamp 1679581782
transform 1 0 97152 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_273
timestamp 1679581782
transform 1 0 97824 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_280
timestamp 1679581782
transform 1 0 98496 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_287
timestamp 1679581782
transform 1 0 99168 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_294
timestamp 1679581782
transform 1 0 99840 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_301
timestamp 1679581782
transform 1 0 100512 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_308
timestamp 1679581782
transform 1 0 101184 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_315
timestamp 1679581782
transform 1 0 101856 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_322
timestamp 1679581782
transform 1 0 102528 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_329
timestamp 1679581782
transform 1 0 103200 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_336
timestamp 1679581782
transform 1 0 103872 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_343
timestamp 1679581782
transform 1 0 104544 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_350
timestamp 1679581782
transform 1 0 105216 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_357
timestamp 1679581782
transform 1 0 105888 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_364
timestamp 1679581782
transform 1 0 106560 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_371
timestamp 1679581782
transform 1 0 107232 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_378
timestamp 1679581782
transform 1 0 107904 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_385
timestamp 1679581782
transform 1 0 108576 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_392
timestamp 1679581782
transform 1 0 109248 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_399
timestamp 1679581782
transform 1 0 109920 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_406
timestamp 1679581782
transform 1 0 110592 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_413
timestamp 1679581782
transform 1 0 111264 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_420
timestamp 1679581782
transform 1 0 111936 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_427
timestamp 1679581782
transform 1 0 112608 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_434
timestamp 1679581782
transform 1 0 113280 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_441
timestamp 1679581782
transform 1 0 113952 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_448
timestamp 1679581782
transform 1 0 114624 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_455
timestamp 1679581782
transform 1 0 115296 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_462
timestamp 1679581782
transform 1 0 115968 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_469
timestamp 1679581782
transform 1 0 116640 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_476
timestamp 1679581782
transform 1 0 117312 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_483
timestamp 1679581782
transform 1 0 117984 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_490
timestamp 1679581782
transform 1 0 118656 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_497
timestamp 1679581782
transform 1 0 119328 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_504
timestamp 1679581782
transform 1 0 120000 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_511
timestamp 1679581782
transform 1 0 120672 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_518
timestamp 1679581782
transform 1 0 121344 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_525
timestamp 1679581782
transform 1 0 122016 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_532
timestamp 1679581782
transform 1 0 122688 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_539
timestamp 1679581782
transform 1 0 123360 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_546
timestamp 1679581782
transform 1 0 124032 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_553
timestamp 1679581782
transform 1 0 124704 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_560
timestamp 1679581782
transform 1 0 125376 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_567
timestamp 1679581782
transform 1 0 126048 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_574
timestamp 1679581782
transform 1 0 126720 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_581
timestamp 1679581782
transform 1 0 127392 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_588
timestamp 1679581782
transform 1 0 128064 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_595
timestamp 1679581782
transform 1 0 128736 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_602
timestamp 1679581782
transform 1 0 129408 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_609
timestamp 1679581782
transform 1 0 130080 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_616
timestamp 1679581782
transform 1 0 130752 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_623
timestamp 1679581782
transform 1 0 131424 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_630
timestamp 1679581782
transform 1 0 132096 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_637
timestamp 1679581782
transform 1 0 132768 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_644
timestamp 1679581782
transform 1 0 133440 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_651
timestamp 1679581782
transform 1 0 134112 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_658
timestamp 1679581782
transform 1 0 134784 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_665
timestamp 1679581782
transform 1 0 135456 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_672
timestamp 1679581782
transform 1 0 136128 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_679
timestamp 1679581782
transform 1 0 136800 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_686
timestamp 1679581782
transform 1 0 137472 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_693
timestamp 1679581782
transform 1 0 138144 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_700
timestamp 1679581782
transform 1 0 138816 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_707
timestamp 1679581782
transform 1 0 139488 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_714
timestamp 1679581782
transform 1 0 140160 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_721
timestamp 1679581782
transform 1 0 140832 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_728
timestamp 1679581782
transform 1 0 141504 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_735
timestamp 1679581782
transform 1 0 142176 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_742
timestamp 1679581782
transform 1 0 142848 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_749
timestamp 1679581782
transform 1 0 143520 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_756
timestamp 1679581782
transform 1 0 144192 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_763
timestamp 1679581782
transform 1 0 144864 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_770
timestamp 1679581782
transform 1 0 145536 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_777
timestamp 1679581782
transform 1 0 146208 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_784
timestamp 1679581782
transform 1 0 146880 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_791
timestamp 1679581782
transform 1 0 147552 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_798
timestamp 1679581782
transform 1 0 148224 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_805
timestamp 1679581782
transform 1 0 148896 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_812
timestamp 1679581782
transform 1 0 149568 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_819
timestamp 1679581782
transform 1 0 150240 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_826
timestamp 1679581782
transform 1 0 150912 0 -1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_833
timestamp 1679581782
transform 1 0 151584 0 -1 92988
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_840
timestamp 1677579658
transform 1 0 152256 0 -1 92988
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_0
timestamp 1679581782
transform 1 0 71616 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_7
timestamp 1679581782
transform 1 0 72288 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_14
timestamp 1679581782
transform 1 0 72960 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_21
timestamp 1679581782
transform 1 0 73632 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_28
timestamp 1679581782
transform 1 0 74304 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_35
timestamp 1679581782
transform 1 0 74976 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_42
timestamp 1679581782
transform 1 0 75648 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_49
timestamp 1679581782
transform 1 0 76320 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_56
timestamp 1679581782
transform 1 0 76992 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_63
timestamp 1679581782
transform 1 0 77664 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_70
timestamp 1679581782
transform 1 0 78336 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_77
timestamp 1679581782
transform 1 0 79008 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_84
timestamp 1679581782
transform 1 0 79680 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_91
timestamp 1679581782
transform 1 0 80352 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_98
timestamp 1679581782
transform 1 0 81024 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_105
timestamp 1679581782
transform 1 0 81696 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_112
timestamp 1679581782
transform 1 0 82368 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_119
timestamp 1679581782
transform 1 0 83040 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_126
timestamp 1679581782
transform 1 0 83712 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_133
timestamp 1679581782
transform 1 0 84384 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_140
timestamp 1679581782
transform 1 0 85056 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_147
timestamp 1679581782
transform 1 0 85728 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_154
timestamp 1679581782
transform 1 0 86400 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_161
timestamp 1679581782
transform 1 0 87072 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_168
timestamp 1679581782
transform 1 0 87744 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_175
timestamp 1679581782
transform 1 0 88416 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_182
timestamp 1679581782
transform 1 0 89088 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_189
timestamp 1679581782
transform 1 0 89760 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_196
timestamp 1679581782
transform 1 0 90432 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_203
timestamp 1679581782
transform 1 0 91104 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_210
timestamp 1679581782
transform 1 0 91776 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_217
timestamp 1679581782
transform 1 0 92448 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_224
timestamp 1679581782
transform 1 0 93120 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_231
timestamp 1679581782
transform 1 0 93792 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_238
timestamp 1679581782
transform 1 0 94464 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_245
timestamp 1679581782
transform 1 0 95136 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_252
timestamp 1679581782
transform 1 0 95808 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_259
timestamp 1679581782
transform 1 0 96480 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_266
timestamp 1679581782
transform 1 0 97152 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_273
timestamp 1679581782
transform 1 0 97824 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_280
timestamp 1679581782
transform 1 0 98496 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_287
timestamp 1679581782
transform 1 0 99168 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_294
timestamp 1679581782
transform 1 0 99840 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_301
timestamp 1679581782
transform 1 0 100512 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_308
timestamp 1679581782
transform 1 0 101184 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_315
timestamp 1679581782
transform 1 0 101856 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_322
timestamp 1679581782
transform 1 0 102528 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_329
timestamp 1679581782
transform 1 0 103200 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_336
timestamp 1679581782
transform 1 0 103872 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_343
timestamp 1679581782
transform 1 0 104544 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_350
timestamp 1679581782
transform 1 0 105216 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_357
timestamp 1679581782
transform 1 0 105888 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_364
timestamp 1679581782
transform 1 0 106560 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_371
timestamp 1679581782
transform 1 0 107232 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_378
timestamp 1679581782
transform 1 0 107904 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_385
timestamp 1679581782
transform 1 0 108576 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_392
timestamp 1679581782
transform 1 0 109248 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_399
timestamp 1679581782
transform 1 0 109920 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_406
timestamp 1679581782
transform 1 0 110592 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_413
timestamp 1679581782
transform 1 0 111264 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_420
timestamp 1679581782
transform 1 0 111936 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_427
timestamp 1679581782
transform 1 0 112608 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_434
timestamp 1679581782
transform 1 0 113280 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_441
timestamp 1679581782
transform 1 0 113952 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_448
timestamp 1679581782
transform 1 0 114624 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_455
timestamp 1679581782
transform 1 0 115296 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_462
timestamp 1679581782
transform 1 0 115968 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_469
timestamp 1679581782
transform 1 0 116640 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_476
timestamp 1679581782
transform 1 0 117312 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_483
timestamp 1679581782
transform 1 0 117984 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_490
timestamp 1679581782
transform 1 0 118656 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_497
timestamp 1679581782
transform 1 0 119328 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_504
timestamp 1679581782
transform 1 0 120000 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_511
timestamp 1679581782
transform 1 0 120672 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_518
timestamp 1679581782
transform 1 0 121344 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_525
timestamp 1679581782
transform 1 0 122016 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_532
timestamp 1679581782
transform 1 0 122688 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_539
timestamp 1679581782
transform 1 0 123360 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_546
timestamp 1679581782
transform 1 0 124032 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_553
timestamp 1679581782
transform 1 0 124704 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_560
timestamp 1679581782
transform 1 0 125376 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_567
timestamp 1679581782
transform 1 0 126048 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_574
timestamp 1679581782
transform 1 0 126720 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_581
timestamp 1679581782
transform 1 0 127392 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_588
timestamp 1679581782
transform 1 0 128064 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_595
timestamp 1679581782
transform 1 0 128736 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_602
timestamp 1679581782
transform 1 0 129408 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_609
timestamp 1679581782
transform 1 0 130080 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_616
timestamp 1679581782
transform 1 0 130752 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_623
timestamp 1679581782
transform 1 0 131424 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_630
timestamp 1679581782
transform 1 0 132096 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_637
timestamp 1679581782
transform 1 0 132768 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_644
timestamp 1679581782
transform 1 0 133440 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_651
timestamp 1679581782
transform 1 0 134112 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_658
timestamp 1679581782
transform 1 0 134784 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_665
timestamp 1679581782
transform 1 0 135456 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_672
timestamp 1679581782
transform 1 0 136128 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_679
timestamp 1679581782
transform 1 0 136800 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_686
timestamp 1679581782
transform 1 0 137472 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_693
timestamp 1679581782
transform 1 0 138144 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_700
timestamp 1679581782
transform 1 0 138816 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_707
timestamp 1679581782
transform 1 0 139488 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_714
timestamp 1679581782
transform 1 0 140160 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_721
timestamp 1679581782
transform 1 0 140832 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_728
timestamp 1679581782
transform 1 0 141504 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_735
timestamp 1679581782
transform 1 0 142176 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_742
timestamp 1679581782
transform 1 0 142848 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_749
timestamp 1679581782
transform 1 0 143520 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_756
timestamp 1679581782
transform 1 0 144192 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_763
timestamp 1679581782
transform 1 0 144864 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_770
timestamp 1679581782
transform 1 0 145536 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_777
timestamp 1679581782
transform 1 0 146208 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_784
timestamp 1679581782
transform 1 0 146880 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_791
timestamp 1679581782
transform 1 0 147552 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_798
timestamp 1679581782
transform 1 0 148224 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_805
timestamp 1679581782
transform 1 0 148896 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_812
timestamp 1679581782
transform 1 0 149568 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_819
timestamp 1679581782
transform 1 0 150240 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_826
timestamp 1679581782
transform 1 0 150912 0 1 92988
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_833
timestamp 1679581782
transform 1 0 151584 0 1 92988
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_840
timestamp 1677579658
transform 1 0 152256 0 1 92988
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_0
timestamp 1679581782
transform 1 0 71616 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_7
timestamp 1679581782
transform 1 0 72288 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_14
timestamp 1679581782
transform 1 0 72960 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_21
timestamp 1679581782
transform 1 0 73632 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_28
timestamp 1679581782
transform 1 0 74304 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_35
timestamp 1679581782
transform 1 0 74976 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_42
timestamp 1679581782
transform 1 0 75648 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_49
timestamp 1679581782
transform 1 0 76320 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_56
timestamp 1679581782
transform 1 0 76992 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_63
timestamp 1679581782
transform 1 0 77664 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_70
timestamp 1679581782
transform 1 0 78336 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_77
timestamp 1679581782
transform 1 0 79008 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_84
timestamp 1679581782
transform 1 0 79680 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_91
timestamp 1679581782
transform 1 0 80352 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_98
timestamp 1679581782
transform 1 0 81024 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_105
timestamp 1679581782
transform 1 0 81696 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_112
timestamp 1679581782
transform 1 0 82368 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_119
timestamp 1679581782
transform 1 0 83040 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_126
timestamp 1679581782
transform 1 0 83712 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_133
timestamp 1679581782
transform 1 0 84384 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_140
timestamp 1679581782
transform 1 0 85056 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_147
timestamp 1679581782
transform 1 0 85728 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_154
timestamp 1679581782
transform 1 0 86400 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_161
timestamp 1679581782
transform 1 0 87072 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_168
timestamp 1679581782
transform 1 0 87744 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_175
timestamp 1679581782
transform 1 0 88416 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_182
timestamp 1679581782
transform 1 0 89088 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_189
timestamp 1679581782
transform 1 0 89760 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_196
timestamp 1679581782
transform 1 0 90432 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_203
timestamp 1679581782
transform 1 0 91104 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_210
timestamp 1679581782
transform 1 0 91776 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_217
timestamp 1679581782
transform 1 0 92448 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_224
timestamp 1679581782
transform 1 0 93120 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_231
timestamp 1679581782
transform 1 0 93792 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_238
timestamp 1679581782
transform 1 0 94464 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_245
timestamp 1679581782
transform 1 0 95136 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_252
timestamp 1679581782
transform 1 0 95808 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_259
timestamp 1679581782
transform 1 0 96480 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_266
timestamp 1679581782
transform 1 0 97152 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_273
timestamp 1679581782
transform 1 0 97824 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_280
timestamp 1679581782
transform 1 0 98496 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_287
timestamp 1679581782
transform 1 0 99168 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_294
timestamp 1679581782
transform 1 0 99840 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_301
timestamp 1679581782
transform 1 0 100512 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_308
timestamp 1679581782
transform 1 0 101184 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_315
timestamp 1679581782
transform 1 0 101856 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_322
timestamp 1679581782
transform 1 0 102528 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_329
timestamp 1679581782
transform 1 0 103200 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_336
timestamp 1679581782
transform 1 0 103872 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_343
timestamp 1679581782
transform 1 0 104544 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_350
timestamp 1679581782
transform 1 0 105216 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_357
timestamp 1679581782
transform 1 0 105888 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_364
timestamp 1679581782
transform 1 0 106560 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_371
timestamp 1679581782
transform 1 0 107232 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_378
timestamp 1679581782
transform 1 0 107904 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_385
timestamp 1679581782
transform 1 0 108576 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_392
timestamp 1679581782
transform 1 0 109248 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_399
timestamp 1679581782
transform 1 0 109920 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_406
timestamp 1679581782
transform 1 0 110592 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_413
timestamp 1679581782
transform 1 0 111264 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_420
timestamp 1679581782
transform 1 0 111936 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_427
timestamp 1679581782
transform 1 0 112608 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_434
timestamp 1679581782
transform 1 0 113280 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_441
timestamp 1679581782
transform 1 0 113952 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_448
timestamp 1679581782
transform 1 0 114624 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_455
timestamp 1679581782
transform 1 0 115296 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_462
timestamp 1679581782
transform 1 0 115968 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_469
timestamp 1679581782
transform 1 0 116640 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_476
timestamp 1679581782
transform 1 0 117312 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_483
timestamp 1679581782
transform 1 0 117984 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_490
timestamp 1679581782
transform 1 0 118656 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_497
timestamp 1679581782
transform 1 0 119328 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_504
timestamp 1679581782
transform 1 0 120000 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_511
timestamp 1679581782
transform 1 0 120672 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_518
timestamp 1679581782
transform 1 0 121344 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_525
timestamp 1679581782
transform 1 0 122016 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_532
timestamp 1679581782
transform 1 0 122688 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_539
timestamp 1679581782
transform 1 0 123360 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_546
timestamp 1679581782
transform 1 0 124032 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_553
timestamp 1679581782
transform 1 0 124704 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_560
timestamp 1679581782
transform 1 0 125376 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_567
timestamp 1679581782
transform 1 0 126048 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_574
timestamp 1679581782
transform 1 0 126720 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_581
timestamp 1679581782
transform 1 0 127392 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_588
timestamp 1679581782
transform 1 0 128064 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_595
timestamp 1679581782
transform 1 0 128736 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_602
timestamp 1679581782
transform 1 0 129408 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_609
timestamp 1679581782
transform 1 0 130080 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_616
timestamp 1679581782
transform 1 0 130752 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_623
timestamp 1679581782
transform 1 0 131424 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_630
timestamp 1679581782
transform 1 0 132096 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_637
timestamp 1679581782
transform 1 0 132768 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_644
timestamp 1679581782
transform 1 0 133440 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_651
timestamp 1679581782
transform 1 0 134112 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_658
timestamp 1679581782
transform 1 0 134784 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_665
timestamp 1679581782
transform 1 0 135456 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_672
timestamp 1679581782
transform 1 0 136128 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_679
timestamp 1679581782
transform 1 0 136800 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_686
timestamp 1679581782
transform 1 0 137472 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_693
timestamp 1679581782
transform 1 0 138144 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_700
timestamp 1679581782
transform 1 0 138816 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_707
timestamp 1679581782
transform 1 0 139488 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_714
timestamp 1679581782
transform 1 0 140160 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_721
timestamp 1679581782
transform 1 0 140832 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_728
timestamp 1679581782
transform 1 0 141504 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_735
timestamp 1679581782
transform 1 0 142176 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_742
timestamp 1679581782
transform 1 0 142848 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_749
timestamp 1679581782
transform 1 0 143520 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_756
timestamp 1679581782
transform 1 0 144192 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_763
timestamp 1679581782
transform 1 0 144864 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_770
timestamp 1679581782
transform 1 0 145536 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_777
timestamp 1679581782
transform 1 0 146208 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_784
timestamp 1679581782
transform 1 0 146880 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_791
timestamp 1679581782
transform 1 0 147552 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_798
timestamp 1679581782
transform 1 0 148224 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_805
timestamp 1679581782
transform 1 0 148896 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_812
timestamp 1679581782
transform 1 0 149568 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_819
timestamp 1679581782
transform 1 0 150240 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_826
timestamp 1679581782
transform 1 0 150912 0 -1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_833
timestamp 1679581782
transform 1 0 151584 0 -1 94500
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_840
timestamp 1677579658
transform 1 0 152256 0 -1 94500
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_0
timestamp 1679581782
transform 1 0 71616 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_7
timestamp 1679581782
transform 1 0 72288 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_14
timestamp 1679581782
transform 1 0 72960 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_21
timestamp 1679581782
transform 1 0 73632 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_28
timestamp 1679581782
transform 1 0 74304 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_35
timestamp 1679581782
transform 1 0 74976 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_42
timestamp 1679581782
transform 1 0 75648 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_49
timestamp 1679581782
transform 1 0 76320 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_56
timestamp 1679581782
transform 1 0 76992 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_63
timestamp 1679581782
transform 1 0 77664 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_70
timestamp 1679581782
transform 1 0 78336 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_77
timestamp 1679581782
transform 1 0 79008 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_84
timestamp 1679581782
transform 1 0 79680 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_91
timestamp 1679581782
transform 1 0 80352 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_98
timestamp 1679581782
transform 1 0 81024 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_105
timestamp 1679581782
transform 1 0 81696 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_112
timestamp 1679581782
transform 1 0 82368 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_119
timestamp 1679581782
transform 1 0 83040 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_126
timestamp 1679581782
transform 1 0 83712 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_133
timestamp 1679581782
transform 1 0 84384 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_140
timestamp 1679581782
transform 1 0 85056 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_147
timestamp 1679581782
transform 1 0 85728 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_154
timestamp 1679581782
transform 1 0 86400 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_161
timestamp 1679581782
transform 1 0 87072 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_168
timestamp 1679581782
transform 1 0 87744 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_175
timestamp 1679581782
transform 1 0 88416 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_182
timestamp 1679581782
transform 1 0 89088 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_189
timestamp 1679581782
transform 1 0 89760 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_196
timestamp 1679581782
transform 1 0 90432 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_203
timestamp 1679581782
transform 1 0 91104 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_210
timestamp 1679581782
transform 1 0 91776 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_217
timestamp 1679581782
transform 1 0 92448 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_224
timestamp 1679581782
transform 1 0 93120 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_231
timestamp 1679581782
transform 1 0 93792 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_238
timestamp 1679581782
transform 1 0 94464 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_245
timestamp 1679581782
transform 1 0 95136 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_252
timestamp 1679581782
transform 1 0 95808 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_259
timestamp 1679581782
transform 1 0 96480 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_266
timestamp 1679581782
transform 1 0 97152 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_273
timestamp 1679581782
transform 1 0 97824 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_280
timestamp 1679581782
transform 1 0 98496 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_287
timestamp 1679581782
transform 1 0 99168 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_294
timestamp 1679581782
transform 1 0 99840 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_301
timestamp 1679581782
transform 1 0 100512 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_308
timestamp 1679581782
transform 1 0 101184 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_315
timestamp 1679581782
transform 1 0 101856 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_322
timestamp 1679581782
transform 1 0 102528 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_329
timestamp 1679581782
transform 1 0 103200 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_336
timestamp 1679581782
transform 1 0 103872 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_343
timestamp 1679581782
transform 1 0 104544 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_350
timestamp 1679581782
transform 1 0 105216 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_357
timestamp 1679581782
transform 1 0 105888 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_364
timestamp 1679581782
transform 1 0 106560 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_371
timestamp 1679581782
transform 1 0 107232 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_378
timestamp 1679581782
transform 1 0 107904 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_385
timestamp 1679581782
transform 1 0 108576 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_392
timestamp 1679581782
transform 1 0 109248 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_399
timestamp 1679581782
transform 1 0 109920 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_406
timestamp 1679581782
transform 1 0 110592 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_413
timestamp 1679581782
transform 1 0 111264 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_420
timestamp 1679581782
transform 1 0 111936 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_427
timestamp 1679581782
transform 1 0 112608 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_434
timestamp 1679581782
transform 1 0 113280 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_441
timestamp 1679581782
transform 1 0 113952 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_448
timestamp 1679581782
transform 1 0 114624 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_455
timestamp 1679581782
transform 1 0 115296 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_462
timestamp 1679581782
transform 1 0 115968 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_469
timestamp 1679581782
transform 1 0 116640 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_476
timestamp 1679581782
transform 1 0 117312 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_483
timestamp 1679581782
transform 1 0 117984 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_490
timestamp 1679581782
transform 1 0 118656 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_497
timestamp 1679581782
transform 1 0 119328 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_504
timestamp 1679581782
transform 1 0 120000 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_511
timestamp 1679581782
transform 1 0 120672 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_518
timestamp 1679581782
transform 1 0 121344 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_525
timestamp 1679581782
transform 1 0 122016 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_532
timestamp 1679581782
transform 1 0 122688 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_539
timestamp 1679581782
transform 1 0 123360 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_546
timestamp 1679581782
transform 1 0 124032 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_553
timestamp 1679581782
transform 1 0 124704 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_560
timestamp 1679581782
transform 1 0 125376 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_567
timestamp 1679581782
transform 1 0 126048 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_574
timestamp 1679581782
transform 1 0 126720 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_581
timestamp 1679581782
transform 1 0 127392 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_588
timestamp 1679581782
transform 1 0 128064 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_595
timestamp 1679581782
transform 1 0 128736 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_602
timestamp 1679581782
transform 1 0 129408 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_609
timestamp 1679581782
transform 1 0 130080 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_616
timestamp 1679581782
transform 1 0 130752 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_623
timestamp 1679581782
transform 1 0 131424 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_630
timestamp 1679581782
transform 1 0 132096 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_637
timestamp 1679581782
transform 1 0 132768 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_644
timestamp 1679581782
transform 1 0 133440 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_651
timestamp 1679581782
transform 1 0 134112 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_658
timestamp 1679581782
transform 1 0 134784 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_665
timestamp 1679581782
transform 1 0 135456 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_672
timestamp 1679581782
transform 1 0 136128 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_679
timestamp 1679581782
transform 1 0 136800 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_686
timestamp 1679581782
transform 1 0 137472 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_693
timestamp 1679581782
transform 1 0 138144 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_700
timestamp 1679581782
transform 1 0 138816 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_707
timestamp 1679581782
transform 1 0 139488 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_714
timestamp 1679581782
transform 1 0 140160 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_721
timestamp 1679581782
transform 1 0 140832 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_728
timestamp 1679581782
transform 1 0 141504 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_735
timestamp 1679581782
transform 1 0 142176 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_742
timestamp 1679581782
transform 1 0 142848 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_749
timestamp 1679581782
transform 1 0 143520 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_756
timestamp 1679581782
transform 1 0 144192 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_763
timestamp 1679581782
transform 1 0 144864 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_770
timestamp 1679581782
transform 1 0 145536 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_777
timestamp 1679581782
transform 1 0 146208 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_784
timestamp 1679581782
transform 1 0 146880 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_791
timestamp 1679581782
transform 1 0 147552 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_798
timestamp 1679581782
transform 1 0 148224 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_805
timestamp 1679581782
transform 1 0 148896 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_812
timestamp 1679581782
transform 1 0 149568 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_819
timestamp 1679581782
transform 1 0 150240 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_826
timestamp 1679581782
transform 1 0 150912 0 1 94500
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_833
timestamp 1679581782
transform 1 0 151584 0 1 94500
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_840
timestamp 1677579658
transform 1 0 152256 0 1 94500
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_0
timestamp 1679581782
transform 1 0 71616 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_7
timestamp 1679581782
transform 1 0 72288 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_14
timestamp 1679581782
transform 1 0 72960 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_21
timestamp 1679581782
transform 1 0 73632 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_28
timestamp 1679581782
transform 1 0 74304 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_35
timestamp 1679581782
transform 1 0 74976 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_42
timestamp 1679581782
transform 1 0 75648 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_49
timestamp 1679581782
transform 1 0 76320 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_56
timestamp 1679581782
transform 1 0 76992 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_63
timestamp 1679581782
transform 1 0 77664 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_70
timestamp 1679581782
transform 1 0 78336 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_77
timestamp 1679581782
transform 1 0 79008 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_84
timestamp 1679581782
transform 1 0 79680 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_91
timestamp 1679581782
transform 1 0 80352 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_98
timestamp 1679581782
transform 1 0 81024 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_105
timestamp 1679581782
transform 1 0 81696 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_112
timestamp 1679581782
transform 1 0 82368 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_119
timestamp 1679581782
transform 1 0 83040 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_126
timestamp 1679581782
transform 1 0 83712 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_133
timestamp 1679581782
transform 1 0 84384 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_140
timestamp 1679581782
transform 1 0 85056 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_147
timestamp 1679581782
transform 1 0 85728 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_154
timestamp 1679581782
transform 1 0 86400 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_161
timestamp 1679581782
transform 1 0 87072 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_168
timestamp 1679581782
transform 1 0 87744 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_175
timestamp 1679581782
transform 1 0 88416 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_182
timestamp 1679581782
transform 1 0 89088 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_189
timestamp 1679581782
transform 1 0 89760 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_196
timestamp 1679581782
transform 1 0 90432 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_203
timestamp 1679581782
transform 1 0 91104 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_210
timestamp 1679581782
transform 1 0 91776 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_217
timestamp 1679581782
transform 1 0 92448 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_224
timestamp 1679581782
transform 1 0 93120 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_231
timestamp 1679581782
transform 1 0 93792 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_238
timestamp 1679581782
transform 1 0 94464 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_245
timestamp 1679581782
transform 1 0 95136 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_252
timestamp 1679581782
transform 1 0 95808 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_259
timestamp 1679581782
transform 1 0 96480 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_266
timestamp 1679581782
transform 1 0 97152 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_273
timestamp 1679581782
transform 1 0 97824 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_280
timestamp 1679581782
transform 1 0 98496 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_287
timestamp 1679581782
transform 1 0 99168 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_294
timestamp 1679581782
transform 1 0 99840 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_301
timestamp 1679581782
transform 1 0 100512 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_308
timestamp 1679581782
transform 1 0 101184 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_315
timestamp 1679581782
transform 1 0 101856 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_322
timestamp 1679581782
transform 1 0 102528 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_329
timestamp 1679581782
transform 1 0 103200 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_336
timestamp 1679581782
transform 1 0 103872 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_343
timestamp 1679581782
transform 1 0 104544 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_350
timestamp 1679581782
transform 1 0 105216 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_357
timestamp 1679581782
transform 1 0 105888 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_364
timestamp 1679581782
transform 1 0 106560 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_371
timestamp 1679581782
transform 1 0 107232 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_378
timestamp 1679581782
transform 1 0 107904 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_385
timestamp 1679581782
transform 1 0 108576 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_392
timestamp 1679581782
transform 1 0 109248 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_399
timestamp 1679581782
transform 1 0 109920 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_406
timestamp 1679581782
transform 1 0 110592 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_413
timestamp 1679581782
transform 1 0 111264 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_420
timestamp 1679581782
transform 1 0 111936 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_427
timestamp 1679581782
transform 1 0 112608 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_434
timestamp 1679581782
transform 1 0 113280 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_441
timestamp 1679581782
transform 1 0 113952 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_448
timestamp 1679581782
transform 1 0 114624 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_455
timestamp 1679581782
transform 1 0 115296 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_462
timestamp 1679581782
transform 1 0 115968 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_469
timestamp 1679581782
transform 1 0 116640 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_476
timestamp 1679581782
transform 1 0 117312 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_483
timestamp 1679581782
transform 1 0 117984 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_490
timestamp 1679581782
transform 1 0 118656 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_497
timestamp 1679581782
transform 1 0 119328 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_504
timestamp 1679581782
transform 1 0 120000 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_511
timestamp 1679581782
transform 1 0 120672 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_518
timestamp 1679581782
transform 1 0 121344 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_525
timestamp 1679581782
transform 1 0 122016 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_532
timestamp 1679581782
transform 1 0 122688 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_539
timestamp 1679581782
transform 1 0 123360 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_546
timestamp 1679581782
transform 1 0 124032 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_553
timestamp 1679581782
transform 1 0 124704 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_560
timestamp 1679581782
transform 1 0 125376 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_567
timestamp 1679581782
transform 1 0 126048 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_574
timestamp 1679581782
transform 1 0 126720 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_581
timestamp 1679581782
transform 1 0 127392 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_588
timestamp 1679581782
transform 1 0 128064 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_595
timestamp 1679581782
transform 1 0 128736 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_602
timestamp 1679581782
transform 1 0 129408 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_609
timestamp 1679581782
transform 1 0 130080 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_616
timestamp 1679581782
transform 1 0 130752 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_623
timestamp 1679581782
transform 1 0 131424 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_630
timestamp 1679581782
transform 1 0 132096 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_637
timestamp 1679581782
transform 1 0 132768 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_644
timestamp 1679581782
transform 1 0 133440 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_651
timestamp 1679581782
transform 1 0 134112 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_658
timestamp 1679581782
transform 1 0 134784 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_665
timestamp 1679581782
transform 1 0 135456 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_672
timestamp 1679581782
transform 1 0 136128 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_679
timestamp 1679581782
transform 1 0 136800 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_686
timestamp 1679581782
transform 1 0 137472 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_693
timestamp 1679581782
transform 1 0 138144 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_700
timestamp 1679581782
transform 1 0 138816 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_707
timestamp 1679581782
transform 1 0 139488 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_714
timestamp 1679581782
transform 1 0 140160 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_721
timestamp 1679581782
transform 1 0 140832 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_728
timestamp 1679581782
transform 1 0 141504 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_735
timestamp 1679581782
transform 1 0 142176 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_742
timestamp 1679581782
transform 1 0 142848 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_749
timestamp 1679581782
transform 1 0 143520 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_756
timestamp 1679581782
transform 1 0 144192 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_763
timestamp 1679581782
transform 1 0 144864 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_770
timestamp 1679581782
transform 1 0 145536 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_777
timestamp 1679581782
transform 1 0 146208 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_784
timestamp 1679581782
transform 1 0 146880 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_791
timestamp 1679581782
transform 1 0 147552 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_798
timestamp 1679581782
transform 1 0 148224 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_805
timestamp 1679581782
transform 1 0 148896 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_812
timestamp 1679581782
transform 1 0 149568 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_819
timestamp 1679581782
transform 1 0 150240 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_826
timestamp 1679581782
transform 1 0 150912 0 -1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_833
timestamp 1679581782
transform 1 0 151584 0 -1 96012
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_840
timestamp 1677579658
transform 1 0 152256 0 -1 96012
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_0
timestamp 1679581782
transform 1 0 71616 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_7
timestamp 1679581782
transform 1 0 72288 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_14
timestamp 1679581782
transform 1 0 72960 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_21
timestamp 1679581782
transform 1 0 73632 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_28
timestamp 1679581782
transform 1 0 74304 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_35
timestamp 1679581782
transform 1 0 74976 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_42
timestamp 1679581782
transform 1 0 75648 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_49
timestamp 1679581782
transform 1 0 76320 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_56
timestamp 1679581782
transform 1 0 76992 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_63
timestamp 1679581782
transform 1 0 77664 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_70
timestamp 1679581782
transform 1 0 78336 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_77
timestamp 1679581782
transform 1 0 79008 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_84
timestamp 1679581782
transform 1 0 79680 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_91
timestamp 1679581782
transform 1 0 80352 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_98
timestamp 1679581782
transform 1 0 81024 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_105
timestamp 1679581782
transform 1 0 81696 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_112
timestamp 1679581782
transform 1 0 82368 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_119
timestamp 1679581782
transform 1 0 83040 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_126
timestamp 1679581782
transform 1 0 83712 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_133
timestamp 1679581782
transform 1 0 84384 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_140
timestamp 1679581782
transform 1 0 85056 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_147
timestamp 1679581782
transform 1 0 85728 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_154
timestamp 1679581782
transform 1 0 86400 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_161
timestamp 1679581782
transform 1 0 87072 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_168
timestamp 1679581782
transform 1 0 87744 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_175
timestamp 1679581782
transform 1 0 88416 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_182
timestamp 1679581782
transform 1 0 89088 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_189
timestamp 1679581782
transform 1 0 89760 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_196
timestamp 1679581782
transform 1 0 90432 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_203
timestamp 1679581782
transform 1 0 91104 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_210
timestamp 1679581782
transform 1 0 91776 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_217
timestamp 1679581782
transform 1 0 92448 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_224
timestamp 1679581782
transform 1 0 93120 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_231
timestamp 1679581782
transform 1 0 93792 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_238
timestamp 1679581782
transform 1 0 94464 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_245
timestamp 1679581782
transform 1 0 95136 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_252
timestamp 1679581782
transform 1 0 95808 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_259
timestamp 1679581782
transform 1 0 96480 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_266
timestamp 1679581782
transform 1 0 97152 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_273
timestamp 1679581782
transform 1 0 97824 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_280
timestamp 1679581782
transform 1 0 98496 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_287
timestamp 1679581782
transform 1 0 99168 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_294
timestamp 1679581782
transform 1 0 99840 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_301
timestamp 1679581782
transform 1 0 100512 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_308
timestamp 1679581782
transform 1 0 101184 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_315
timestamp 1679581782
transform 1 0 101856 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_322
timestamp 1679581782
transform 1 0 102528 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_329
timestamp 1679581782
transform 1 0 103200 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_336
timestamp 1679581782
transform 1 0 103872 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_343
timestamp 1679581782
transform 1 0 104544 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_350
timestamp 1679581782
transform 1 0 105216 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_357
timestamp 1679581782
transform 1 0 105888 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_364
timestamp 1679581782
transform 1 0 106560 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_371
timestamp 1679581782
transform 1 0 107232 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_378
timestamp 1679581782
transform 1 0 107904 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_385
timestamp 1679581782
transform 1 0 108576 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_392
timestamp 1679581782
transform 1 0 109248 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_399
timestamp 1679581782
transform 1 0 109920 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_406
timestamp 1679581782
transform 1 0 110592 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_413
timestamp 1679581782
transform 1 0 111264 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_420
timestamp 1679581782
transform 1 0 111936 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_427
timestamp 1679581782
transform 1 0 112608 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_434
timestamp 1679581782
transform 1 0 113280 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_441
timestamp 1679581782
transform 1 0 113952 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_448
timestamp 1679581782
transform 1 0 114624 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_455
timestamp 1679581782
transform 1 0 115296 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_462
timestamp 1679581782
transform 1 0 115968 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_469
timestamp 1679581782
transform 1 0 116640 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_476
timestamp 1679581782
transform 1 0 117312 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_483
timestamp 1679581782
transform 1 0 117984 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_490
timestamp 1679581782
transform 1 0 118656 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_497
timestamp 1679581782
transform 1 0 119328 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_504
timestamp 1679581782
transform 1 0 120000 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_511
timestamp 1679581782
transform 1 0 120672 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_518
timestamp 1679581782
transform 1 0 121344 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_525
timestamp 1679581782
transform 1 0 122016 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_532
timestamp 1679581782
transform 1 0 122688 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_539
timestamp 1679581782
transform 1 0 123360 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_546
timestamp 1679581782
transform 1 0 124032 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_553
timestamp 1679581782
transform 1 0 124704 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_560
timestamp 1679581782
transform 1 0 125376 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_567
timestamp 1679581782
transform 1 0 126048 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_574
timestamp 1679581782
transform 1 0 126720 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_581
timestamp 1679581782
transform 1 0 127392 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_588
timestamp 1679581782
transform 1 0 128064 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_595
timestamp 1679581782
transform 1 0 128736 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_602
timestamp 1679581782
transform 1 0 129408 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_609
timestamp 1679581782
transform 1 0 130080 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_616
timestamp 1679581782
transform 1 0 130752 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_623
timestamp 1679581782
transform 1 0 131424 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_630
timestamp 1679581782
transform 1 0 132096 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_637
timestamp 1679581782
transform 1 0 132768 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_644
timestamp 1679581782
transform 1 0 133440 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_651
timestamp 1679581782
transform 1 0 134112 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_658
timestamp 1679581782
transform 1 0 134784 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_665
timestamp 1679581782
transform 1 0 135456 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_672
timestamp 1679581782
transform 1 0 136128 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_679
timestamp 1679581782
transform 1 0 136800 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_686
timestamp 1679581782
transform 1 0 137472 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_693
timestamp 1679581782
transform 1 0 138144 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_700
timestamp 1679581782
transform 1 0 138816 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_707
timestamp 1679581782
transform 1 0 139488 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_714
timestamp 1679581782
transform 1 0 140160 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_721
timestamp 1679581782
transform 1 0 140832 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_728
timestamp 1679581782
transform 1 0 141504 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_735
timestamp 1679581782
transform 1 0 142176 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_742
timestamp 1679581782
transform 1 0 142848 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_749
timestamp 1679581782
transform 1 0 143520 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_756
timestamp 1679581782
transform 1 0 144192 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_763
timestamp 1679581782
transform 1 0 144864 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_770
timestamp 1679581782
transform 1 0 145536 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_777
timestamp 1679581782
transform 1 0 146208 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_784
timestamp 1679581782
transform 1 0 146880 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_791
timestamp 1679581782
transform 1 0 147552 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_798
timestamp 1679581782
transform 1 0 148224 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_805
timestamp 1679581782
transform 1 0 148896 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_812
timestamp 1679581782
transform 1 0 149568 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_819
timestamp 1679581782
transform 1 0 150240 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_826
timestamp 1679581782
transform 1 0 150912 0 1 96012
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_833
timestamp 1679581782
transform 1 0 151584 0 1 96012
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_840
timestamp 1677579658
transform 1 0 152256 0 1 96012
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679581782
transform 1 0 71616 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1679581782
transform 1 0 72288 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1679581782
transform 1 0 72960 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_21
timestamp 1679581782
transform 1 0 73632 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_28
timestamp 1679581782
transform 1 0 74304 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_35
timestamp 1679581782
transform 1 0 74976 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_42
timestamp 1679581782
transform 1 0 75648 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_49
timestamp 1679581782
transform 1 0 76320 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_56
timestamp 1679581782
transform 1 0 76992 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_63
timestamp 1679581782
transform 1 0 77664 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_70
timestamp 1679581782
transform 1 0 78336 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_77
timestamp 1679581782
transform 1 0 79008 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_84
timestamp 1679581782
transform 1 0 79680 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_91
timestamp 1679581782
transform 1 0 80352 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_98
timestamp 1679581782
transform 1 0 81024 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_105
timestamp 1679581782
transform 1 0 81696 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_112
timestamp 1679581782
transform 1 0 82368 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_119
timestamp 1679581782
transform 1 0 83040 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_126
timestamp 1679581782
transform 1 0 83712 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_133
timestamp 1679581782
transform 1 0 84384 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_140
timestamp 1679581782
transform 1 0 85056 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_147
timestamp 1679581782
transform 1 0 85728 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_154
timestamp 1679581782
transform 1 0 86400 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_161
timestamp 1679581782
transform 1 0 87072 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_168
timestamp 1679581782
transform 1 0 87744 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_175
timestamp 1679581782
transform 1 0 88416 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_182
timestamp 1679581782
transform 1 0 89088 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_189
timestamp 1679581782
transform 1 0 89760 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_196
timestamp 1679581782
transform 1 0 90432 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_203
timestamp 1679581782
transform 1 0 91104 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_210
timestamp 1679581782
transform 1 0 91776 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_217
timestamp 1679581782
transform 1 0 92448 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_224
timestamp 1679581782
transform 1 0 93120 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_231
timestamp 1679581782
transform 1 0 93792 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_238
timestamp 1679581782
transform 1 0 94464 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_245
timestamp 1679581782
transform 1 0 95136 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_252
timestamp 1679581782
transform 1 0 95808 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_259
timestamp 1679581782
transform 1 0 96480 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_266
timestamp 1679581782
transform 1 0 97152 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_273
timestamp 1679581782
transform 1 0 97824 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_280
timestamp 1679581782
transform 1 0 98496 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_287
timestamp 1679581782
transform 1 0 99168 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_294
timestamp 1679581782
transform 1 0 99840 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_301
timestamp 1679581782
transform 1 0 100512 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_308
timestamp 1679581782
transform 1 0 101184 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_315
timestamp 1679581782
transform 1 0 101856 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_322
timestamp 1679581782
transform 1 0 102528 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_329
timestamp 1679581782
transform 1 0 103200 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_336
timestamp 1679581782
transform 1 0 103872 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_343
timestamp 1679581782
transform 1 0 104544 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_350
timestamp 1679581782
transform 1 0 105216 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_357
timestamp 1679581782
transform 1 0 105888 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_364
timestamp 1679581782
transform 1 0 106560 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_371
timestamp 1679581782
transform 1 0 107232 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_378
timestamp 1679581782
transform 1 0 107904 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_385
timestamp 1679581782
transform 1 0 108576 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_392
timestamp 1679581782
transform 1 0 109248 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_399
timestamp 1679581782
transform 1 0 109920 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_406
timestamp 1679581782
transform 1 0 110592 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_413
timestamp 1679581782
transform 1 0 111264 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_420
timestamp 1679581782
transform 1 0 111936 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_427
timestamp 1679581782
transform 1 0 112608 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_434
timestamp 1679581782
transform 1 0 113280 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_441
timestamp 1679581782
transform 1 0 113952 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_448
timestamp 1679581782
transform 1 0 114624 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_455
timestamp 1679581782
transform 1 0 115296 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_462
timestamp 1679581782
transform 1 0 115968 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_469
timestamp 1679581782
transform 1 0 116640 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_476
timestamp 1679581782
transform 1 0 117312 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_483
timestamp 1679581782
transform 1 0 117984 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_490
timestamp 1679581782
transform 1 0 118656 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_497
timestamp 1679581782
transform 1 0 119328 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_504
timestamp 1679581782
transform 1 0 120000 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_511
timestamp 1679581782
transform 1 0 120672 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_518
timestamp 1679581782
transform 1 0 121344 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_525
timestamp 1679581782
transform 1 0 122016 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_532
timestamp 1679581782
transform 1 0 122688 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_539
timestamp 1679581782
transform 1 0 123360 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_546
timestamp 1679581782
transform 1 0 124032 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_553
timestamp 1679581782
transform 1 0 124704 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_560
timestamp 1679581782
transform 1 0 125376 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_567
timestamp 1679581782
transform 1 0 126048 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_574
timestamp 1679581782
transform 1 0 126720 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_581
timestamp 1679581782
transform 1 0 127392 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_588
timestamp 1679581782
transform 1 0 128064 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_595
timestamp 1679581782
transform 1 0 128736 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_602
timestamp 1679581782
transform 1 0 129408 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_609
timestamp 1679581782
transform 1 0 130080 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_616
timestamp 1679581782
transform 1 0 130752 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_623
timestamp 1679581782
transform 1 0 131424 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_630
timestamp 1679581782
transform 1 0 132096 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_637
timestamp 1679581782
transform 1 0 132768 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_644
timestamp 1679581782
transform 1 0 133440 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_651
timestamp 1679581782
transform 1 0 134112 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_658
timestamp 1679581782
transform 1 0 134784 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_665
timestamp 1679581782
transform 1 0 135456 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_672
timestamp 1679581782
transform 1 0 136128 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_679
timestamp 1679581782
transform 1 0 136800 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_686
timestamp 1679581782
transform 1 0 137472 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_693
timestamp 1679581782
transform 1 0 138144 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_700
timestamp 1679581782
transform 1 0 138816 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_707
timestamp 1679581782
transform 1 0 139488 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_714
timestamp 1679581782
transform 1 0 140160 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_721
timestamp 1679581782
transform 1 0 140832 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_728
timestamp 1679581782
transform 1 0 141504 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_735
timestamp 1679581782
transform 1 0 142176 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_742
timestamp 1679581782
transform 1 0 142848 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_749
timestamp 1679581782
transform 1 0 143520 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_756
timestamp 1679581782
transform 1 0 144192 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_763
timestamp 1679581782
transform 1 0 144864 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_770
timestamp 1679581782
transform 1 0 145536 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_777
timestamp 1679581782
transform 1 0 146208 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_784
timestamp 1679581782
transform 1 0 146880 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_791
timestamp 1679581782
transform 1 0 147552 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_798
timestamp 1679581782
transform 1 0 148224 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_805
timestamp 1679581782
transform 1 0 148896 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_812
timestamp 1679581782
transform 1 0 149568 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_819
timestamp 1679581782
transform 1 0 150240 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_826
timestamp 1679581782
transform 1 0 150912 0 -1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_833
timestamp 1679581782
transform 1 0 151584 0 -1 97524
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_840
timestamp 1677579658
transform 1 0 152256 0 -1 97524
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 71616 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679581782
transform 1 0 72288 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679581782
transform 1 0 72960 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679581782
transform 1 0 73632 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679581782
transform 1 0 74304 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_35
timestamp 1679581782
transform 1 0 74976 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_42
timestamp 1679581782
transform 1 0 75648 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679581782
transform 1 0 76320 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_56
timestamp 1679581782
transform 1 0 76992 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_63
timestamp 1679581782
transform 1 0 77664 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_70
timestamp 1679581782
transform 1 0 78336 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_77
timestamp 1679581782
transform 1 0 79008 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_84
timestamp 1679581782
transform 1 0 79680 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_91
timestamp 1679581782
transform 1 0 80352 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_98
timestamp 1679581782
transform 1 0 81024 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_105
timestamp 1679581782
transform 1 0 81696 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_112
timestamp 1679581782
transform 1 0 82368 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_119
timestamp 1679581782
transform 1 0 83040 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_126
timestamp 1679581782
transform 1 0 83712 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_133
timestamp 1679581782
transform 1 0 84384 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_140
timestamp 1679581782
transform 1 0 85056 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_147
timestamp 1679581782
transform 1 0 85728 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_154
timestamp 1679581782
transform 1 0 86400 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_161
timestamp 1679581782
transform 1 0 87072 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_168
timestamp 1679581782
transform 1 0 87744 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_175
timestamp 1679581782
transform 1 0 88416 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_182
timestamp 1679581782
transform 1 0 89088 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_189
timestamp 1679581782
transform 1 0 89760 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_196
timestamp 1679581782
transform 1 0 90432 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_203
timestamp 1679581782
transform 1 0 91104 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_210
timestamp 1679581782
transform 1 0 91776 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_217
timestamp 1679581782
transform 1 0 92448 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_224
timestamp 1679581782
transform 1 0 93120 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_231
timestamp 1679581782
transform 1 0 93792 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_238
timestamp 1679581782
transform 1 0 94464 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_245
timestamp 1679581782
transform 1 0 95136 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_252
timestamp 1679581782
transform 1 0 95808 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_259
timestamp 1679581782
transform 1 0 96480 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_266
timestamp 1679581782
transform 1 0 97152 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_273
timestamp 1679581782
transform 1 0 97824 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_280
timestamp 1679581782
transform 1 0 98496 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_287
timestamp 1679581782
transform 1 0 99168 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_294
timestamp 1679581782
transform 1 0 99840 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_301
timestamp 1679581782
transform 1 0 100512 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_308
timestamp 1679581782
transform 1 0 101184 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_315
timestamp 1679581782
transform 1 0 101856 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_322
timestamp 1679581782
transform 1 0 102528 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_329
timestamp 1679581782
transform 1 0 103200 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_336
timestamp 1679581782
transform 1 0 103872 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_343
timestamp 1679581782
transform 1 0 104544 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_350
timestamp 1679581782
transform 1 0 105216 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_357
timestamp 1679581782
transform 1 0 105888 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_364
timestamp 1679581782
transform 1 0 106560 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_371
timestamp 1679581782
transform 1 0 107232 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_378
timestamp 1679581782
transform 1 0 107904 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_385
timestamp 1679581782
transform 1 0 108576 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_392
timestamp 1679581782
transform 1 0 109248 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_399
timestamp 1679581782
transform 1 0 109920 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_406
timestamp 1679581782
transform 1 0 110592 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_413
timestamp 1679581782
transform 1 0 111264 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_420
timestamp 1679581782
transform 1 0 111936 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_427
timestamp 1679581782
transform 1 0 112608 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_434
timestamp 1679581782
transform 1 0 113280 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_441
timestamp 1679581782
transform 1 0 113952 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_448
timestamp 1679581782
transform 1 0 114624 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_455
timestamp 1679581782
transform 1 0 115296 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_462
timestamp 1679581782
transform 1 0 115968 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_469
timestamp 1679581782
transform 1 0 116640 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_476
timestamp 1679581782
transform 1 0 117312 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_483
timestamp 1679581782
transform 1 0 117984 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_490
timestamp 1679581782
transform 1 0 118656 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_497
timestamp 1679581782
transform 1 0 119328 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_504
timestamp 1679581782
transform 1 0 120000 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_511
timestamp 1679581782
transform 1 0 120672 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_518
timestamp 1679581782
transform 1 0 121344 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_525
timestamp 1679581782
transform 1 0 122016 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_532
timestamp 1679581782
transform 1 0 122688 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_539
timestamp 1679581782
transform 1 0 123360 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_546
timestamp 1679581782
transform 1 0 124032 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_553
timestamp 1679581782
transform 1 0 124704 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_560
timestamp 1679581782
transform 1 0 125376 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_567
timestamp 1679581782
transform 1 0 126048 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_574
timestamp 1679581782
transform 1 0 126720 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_581
timestamp 1679581782
transform 1 0 127392 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_588
timestamp 1679581782
transform 1 0 128064 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_595
timestamp 1679581782
transform 1 0 128736 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_602
timestamp 1679581782
transform 1 0 129408 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_609
timestamp 1679581782
transform 1 0 130080 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_616
timestamp 1679581782
transform 1 0 130752 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_623
timestamp 1679581782
transform 1 0 131424 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_630
timestamp 1679581782
transform 1 0 132096 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_637
timestamp 1679581782
transform 1 0 132768 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_644
timestamp 1679581782
transform 1 0 133440 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_651
timestamp 1679581782
transform 1 0 134112 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_658
timestamp 1679581782
transform 1 0 134784 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_665
timestamp 1679581782
transform 1 0 135456 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_672
timestamp 1679581782
transform 1 0 136128 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_679
timestamp 1679581782
transform 1 0 136800 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_686
timestamp 1679581782
transform 1 0 137472 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_693
timestamp 1679581782
transform 1 0 138144 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_700
timestamp 1679581782
transform 1 0 138816 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_707
timestamp 1679581782
transform 1 0 139488 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_714
timestamp 1679581782
transform 1 0 140160 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_721
timestamp 1679581782
transform 1 0 140832 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_728
timestamp 1679581782
transform 1 0 141504 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_735
timestamp 1679581782
transform 1 0 142176 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_742
timestamp 1679581782
transform 1 0 142848 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_749
timestamp 1679581782
transform 1 0 143520 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_756
timestamp 1679581782
transform 1 0 144192 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_763
timestamp 1679581782
transform 1 0 144864 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_770
timestamp 1679581782
transform 1 0 145536 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_777
timestamp 1679581782
transform 1 0 146208 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_784
timestamp 1679581782
transform 1 0 146880 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_791
timestamp 1679581782
transform 1 0 147552 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_798
timestamp 1679581782
transform 1 0 148224 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_805
timestamp 1679581782
transform 1 0 148896 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_812
timestamp 1679581782
transform 1 0 149568 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_819
timestamp 1679581782
transform 1 0 150240 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_826
timestamp 1679581782
transform 1 0 150912 0 1 97524
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_833
timestamp 1679581782
transform 1 0 151584 0 1 97524
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_840
timestamp 1677579658
transform 1 0 152256 0 1 97524
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 71616 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679581782
transform 1 0 72288 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679581782
transform 1 0 72960 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679581782
transform 1 0 73632 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_28
timestamp 1679581782
transform 1 0 74304 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_35
timestamp 1679581782
transform 1 0 74976 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_42
timestamp 1679581782
transform 1 0 75648 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_49
timestamp 1679581782
transform 1 0 76320 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_56
timestamp 1679581782
transform 1 0 76992 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_63
timestamp 1679581782
transform 1 0 77664 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_70
timestamp 1679581782
transform 1 0 78336 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_77
timestamp 1679581782
transform 1 0 79008 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_84
timestamp 1679581782
transform 1 0 79680 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_91
timestamp 1679581782
transform 1 0 80352 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_98
timestamp 1679581782
transform 1 0 81024 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_105
timestamp 1679581782
transform 1 0 81696 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_112
timestamp 1679581782
transform 1 0 82368 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_119
timestamp 1679581782
transform 1 0 83040 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_126
timestamp 1679581782
transform 1 0 83712 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_133
timestamp 1679581782
transform 1 0 84384 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_140
timestamp 1679581782
transform 1 0 85056 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_147
timestamp 1679581782
transform 1 0 85728 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_154
timestamp 1679581782
transform 1 0 86400 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_161
timestamp 1679581782
transform 1 0 87072 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_168
timestamp 1679581782
transform 1 0 87744 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_175
timestamp 1679581782
transform 1 0 88416 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_182
timestamp 1679581782
transform 1 0 89088 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_189
timestamp 1679581782
transform 1 0 89760 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_196
timestamp 1679581782
transform 1 0 90432 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_203
timestamp 1679581782
transform 1 0 91104 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_210
timestamp 1679581782
transform 1 0 91776 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_217
timestamp 1679581782
transform 1 0 92448 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_224
timestamp 1679581782
transform 1 0 93120 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_231
timestamp 1679581782
transform 1 0 93792 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_238
timestamp 1679581782
transform 1 0 94464 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_245
timestamp 1679581782
transform 1 0 95136 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_252
timestamp 1679581782
transform 1 0 95808 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_259
timestamp 1679581782
transform 1 0 96480 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_266
timestamp 1679581782
transform 1 0 97152 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_273
timestamp 1679581782
transform 1 0 97824 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_280
timestamp 1679581782
transform 1 0 98496 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_287
timestamp 1679581782
transform 1 0 99168 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_294
timestamp 1679581782
transform 1 0 99840 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_301
timestamp 1679581782
transform 1 0 100512 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_308
timestamp 1679581782
transform 1 0 101184 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_315
timestamp 1679581782
transform 1 0 101856 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_322
timestamp 1679581782
transform 1 0 102528 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_329
timestamp 1679581782
transform 1 0 103200 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_336
timestamp 1679581782
transform 1 0 103872 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_343
timestamp 1679581782
transform 1 0 104544 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_350
timestamp 1679581782
transform 1 0 105216 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_357
timestamp 1679581782
transform 1 0 105888 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_364
timestamp 1679581782
transform 1 0 106560 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_371
timestamp 1679581782
transform 1 0 107232 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_378
timestamp 1679581782
transform 1 0 107904 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_385
timestamp 1679581782
transform 1 0 108576 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_392
timestamp 1679581782
transform 1 0 109248 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_399
timestamp 1679581782
transform 1 0 109920 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_406
timestamp 1679581782
transform 1 0 110592 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_413
timestamp 1679581782
transform 1 0 111264 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_420
timestamp 1679581782
transform 1 0 111936 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_427
timestamp 1679581782
transform 1 0 112608 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_434
timestamp 1679581782
transform 1 0 113280 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_441
timestamp 1679581782
transform 1 0 113952 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_448
timestamp 1679581782
transform 1 0 114624 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_455
timestamp 1679581782
transform 1 0 115296 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_462
timestamp 1679581782
transform 1 0 115968 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_469
timestamp 1679581782
transform 1 0 116640 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_476
timestamp 1679581782
transform 1 0 117312 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_483
timestamp 1679581782
transform 1 0 117984 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_490
timestamp 1679581782
transform 1 0 118656 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_497
timestamp 1679581782
transform 1 0 119328 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_504
timestamp 1679581782
transform 1 0 120000 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_511
timestamp 1679581782
transform 1 0 120672 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_518
timestamp 1679581782
transform 1 0 121344 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_525
timestamp 1679581782
transform 1 0 122016 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_532
timestamp 1679581782
transform 1 0 122688 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_539
timestamp 1679581782
transform 1 0 123360 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_546
timestamp 1679581782
transform 1 0 124032 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_553
timestamp 1679581782
transform 1 0 124704 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_560
timestamp 1679581782
transform 1 0 125376 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_567
timestamp 1679581782
transform 1 0 126048 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_574
timestamp 1679581782
transform 1 0 126720 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_581
timestamp 1679581782
transform 1 0 127392 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_588
timestamp 1679581782
transform 1 0 128064 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_595
timestamp 1679581782
transform 1 0 128736 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_602
timestamp 1679581782
transform 1 0 129408 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_609
timestamp 1679581782
transform 1 0 130080 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_616
timestamp 1679581782
transform 1 0 130752 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_623
timestamp 1679581782
transform 1 0 131424 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_630
timestamp 1679581782
transform 1 0 132096 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_637
timestamp 1679581782
transform 1 0 132768 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_644
timestamp 1679581782
transform 1 0 133440 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_651
timestamp 1679581782
transform 1 0 134112 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_658
timestamp 1679581782
transform 1 0 134784 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_665
timestamp 1679581782
transform 1 0 135456 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_672
timestamp 1679581782
transform 1 0 136128 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_679
timestamp 1679581782
transform 1 0 136800 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_686
timestamp 1679581782
transform 1 0 137472 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_693
timestamp 1679581782
transform 1 0 138144 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_700
timestamp 1679581782
transform 1 0 138816 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_707
timestamp 1679581782
transform 1 0 139488 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_714
timestamp 1679581782
transform 1 0 140160 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_721
timestamp 1679581782
transform 1 0 140832 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_728
timestamp 1679581782
transform 1 0 141504 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_735
timestamp 1679581782
transform 1 0 142176 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_742
timestamp 1679581782
transform 1 0 142848 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_749
timestamp 1679581782
transform 1 0 143520 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_756
timestamp 1679581782
transform 1 0 144192 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_763
timestamp 1679581782
transform 1 0 144864 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_770
timestamp 1679581782
transform 1 0 145536 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_777
timestamp 1679581782
transform 1 0 146208 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_784
timestamp 1679581782
transform 1 0 146880 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_791
timestamp 1679581782
transform 1 0 147552 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_798
timestamp 1679581782
transform 1 0 148224 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_805
timestamp 1679581782
transform 1 0 148896 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_812
timestamp 1679581782
transform 1 0 149568 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_819
timestamp 1679581782
transform 1 0 150240 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_826
timestamp 1679581782
transform 1 0 150912 0 -1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_833
timestamp 1679581782
transform 1 0 151584 0 -1 99036
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_840
timestamp 1677579658
transform 1 0 152256 0 -1 99036
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 71616 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679581782
transform 1 0 72288 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679581782
transform 1 0 72960 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679581782
transform 1 0 73632 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679581782
transform 1 0 74304 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679581782
transform 1 0 74976 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679581782
transform 1 0 75648 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679581782
transform 1 0 76320 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_56
timestamp 1679581782
transform 1 0 76992 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_63
timestamp 1679581782
transform 1 0 77664 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_70
timestamp 1679581782
transform 1 0 78336 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_77
timestamp 1679581782
transform 1 0 79008 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_84
timestamp 1679581782
transform 1 0 79680 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_91
timestamp 1679581782
transform 1 0 80352 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_98
timestamp 1679581782
transform 1 0 81024 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_105
timestamp 1679581782
transform 1 0 81696 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_112
timestamp 1679581782
transform 1 0 82368 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_119
timestamp 1679581782
transform 1 0 83040 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679581782
transform 1 0 83712 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_133
timestamp 1679581782
transform 1 0 84384 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_140
timestamp 1679581782
transform 1 0 85056 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_147
timestamp 1679581782
transform 1 0 85728 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_154
timestamp 1679581782
transform 1 0 86400 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_161
timestamp 1679581782
transform 1 0 87072 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_168
timestamp 1679581782
transform 1 0 87744 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_175
timestamp 1679581782
transform 1 0 88416 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_182
timestamp 1679581782
transform 1 0 89088 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_189
timestamp 1679581782
transform 1 0 89760 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_196
timestamp 1679581782
transform 1 0 90432 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_203
timestamp 1679581782
transform 1 0 91104 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_210
timestamp 1679581782
transform 1 0 91776 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_217
timestamp 1679581782
transform 1 0 92448 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_224
timestamp 1679581782
transform 1 0 93120 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_231
timestamp 1679581782
transform 1 0 93792 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_238
timestamp 1679581782
transform 1 0 94464 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_245
timestamp 1679581782
transform 1 0 95136 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_252
timestamp 1679581782
transform 1 0 95808 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_259
timestamp 1679581782
transform 1 0 96480 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_266
timestamp 1679581782
transform 1 0 97152 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_273
timestamp 1679581782
transform 1 0 97824 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_280
timestamp 1679581782
transform 1 0 98496 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_287
timestamp 1679581782
transform 1 0 99168 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_294
timestamp 1679581782
transform 1 0 99840 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_301
timestamp 1679581782
transform 1 0 100512 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_308
timestamp 1679581782
transform 1 0 101184 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_315
timestamp 1679581782
transform 1 0 101856 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_322
timestamp 1679581782
transform 1 0 102528 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_329
timestamp 1679581782
transform 1 0 103200 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_336
timestamp 1679581782
transform 1 0 103872 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_343
timestamp 1679581782
transform 1 0 104544 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_350
timestamp 1679581782
transform 1 0 105216 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_357
timestamp 1679581782
transform 1 0 105888 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_364
timestamp 1679581782
transform 1 0 106560 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_371
timestamp 1679581782
transform 1 0 107232 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_378
timestamp 1679581782
transform 1 0 107904 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_385
timestamp 1679581782
transform 1 0 108576 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_392
timestamp 1679581782
transform 1 0 109248 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_399
timestamp 1679581782
transform 1 0 109920 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_406
timestamp 1679581782
transform 1 0 110592 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_413
timestamp 1679581782
transform 1 0 111264 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_420
timestamp 1679581782
transform 1 0 111936 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_427
timestamp 1679581782
transform 1 0 112608 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_434
timestamp 1679581782
transform 1 0 113280 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_441
timestamp 1679581782
transform 1 0 113952 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_448
timestamp 1679581782
transform 1 0 114624 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_455
timestamp 1679581782
transform 1 0 115296 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_462
timestamp 1679581782
transform 1 0 115968 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_469
timestamp 1679581782
transform 1 0 116640 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_476
timestamp 1679581782
transform 1 0 117312 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_483
timestamp 1679581782
transform 1 0 117984 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_490
timestamp 1679581782
transform 1 0 118656 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_497
timestamp 1679581782
transform 1 0 119328 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_504
timestamp 1679581782
transform 1 0 120000 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_511
timestamp 1679581782
transform 1 0 120672 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_518
timestamp 1679581782
transform 1 0 121344 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_525
timestamp 1679581782
transform 1 0 122016 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_532
timestamp 1679581782
transform 1 0 122688 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_539
timestamp 1679581782
transform 1 0 123360 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_546
timestamp 1679581782
transform 1 0 124032 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_553
timestamp 1679581782
transform 1 0 124704 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_560
timestamp 1679581782
transform 1 0 125376 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_567
timestamp 1679581782
transform 1 0 126048 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_574
timestamp 1679581782
transform 1 0 126720 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_581
timestamp 1679581782
transform 1 0 127392 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_588
timestamp 1679581782
transform 1 0 128064 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_595
timestamp 1679581782
transform 1 0 128736 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_602
timestamp 1679581782
transform 1 0 129408 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_609
timestamp 1679581782
transform 1 0 130080 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_616
timestamp 1679581782
transform 1 0 130752 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_623
timestamp 1679581782
transform 1 0 131424 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_630
timestamp 1679581782
transform 1 0 132096 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_637
timestamp 1679581782
transform 1 0 132768 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_644
timestamp 1679581782
transform 1 0 133440 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_651
timestamp 1679581782
transform 1 0 134112 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_658
timestamp 1679581782
transform 1 0 134784 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_665
timestamp 1679581782
transform 1 0 135456 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_672
timestamp 1679581782
transform 1 0 136128 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_679
timestamp 1679581782
transform 1 0 136800 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_686
timestamp 1679581782
transform 1 0 137472 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_693
timestamp 1679581782
transform 1 0 138144 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_700
timestamp 1679581782
transform 1 0 138816 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_707
timestamp 1679581782
transform 1 0 139488 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_714
timestamp 1679581782
transform 1 0 140160 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_721
timestamp 1679581782
transform 1 0 140832 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_728
timestamp 1679581782
transform 1 0 141504 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_735
timestamp 1679581782
transform 1 0 142176 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_742
timestamp 1679581782
transform 1 0 142848 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_749
timestamp 1679581782
transform 1 0 143520 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_756
timestamp 1679581782
transform 1 0 144192 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_763
timestamp 1679581782
transform 1 0 144864 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_770
timestamp 1679581782
transform 1 0 145536 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_777
timestamp 1679581782
transform 1 0 146208 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_784
timestamp 1679581782
transform 1 0 146880 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_791
timestamp 1679581782
transform 1 0 147552 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_798
timestamp 1679581782
transform 1 0 148224 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_805
timestamp 1679581782
transform 1 0 148896 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_812
timestamp 1679581782
transform 1 0 149568 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_819
timestamp 1679581782
transform 1 0 150240 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_826
timestamp 1679581782
transform 1 0 150912 0 1 99036
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_833
timestamp 1679581782
transform 1 0 151584 0 1 99036
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_840
timestamp 1677579658
transform 1 0 152256 0 1 99036
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679581782
transform 1 0 71616 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679581782
transform 1 0 72288 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679581782
transform 1 0 72960 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679581782
transform 1 0 73632 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679581782
transform 1 0 74304 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679581782
transform 1 0 74976 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679581782
transform 1 0 75648 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679581782
transform 1 0 76320 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679581782
transform 1 0 76992 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679581782
transform 1 0 77664 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_70
timestamp 1679581782
transform 1 0 78336 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_77
timestamp 1679581782
transform 1 0 79008 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_84
timestamp 1679581782
transform 1 0 79680 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_91
timestamp 1679581782
transform 1 0 80352 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679581782
transform 1 0 81024 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679581782
transform 1 0 81696 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679581782
transform 1 0 82368 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679581782
transform 1 0 83040 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679581782
transform 1 0 83712 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679581782
transform 1 0 84384 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679581782
transform 1 0 85056 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_147
timestamp 1679581782
transform 1 0 85728 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_154
timestamp 1679581782
transform 1 0 86400 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_161
timestamp 1679581782
transform 1 0 87072 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_168
timestamp 1679581782
transform 1 0 87744 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_175
timestamp 1679581782
transform 1 0 88416 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_182
timestamp 1679581782
transform 1 0 89088 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_189
timestamp 1679581782
transform 1 0 89760 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_196
timestamp 1679581782
transform 1 0 90432 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_203
timestamp 1679581782
transform 1 0 91104 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_210
timestamp 1679581782
transform 1 0 91776 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_217
timestamp 1679581782
transform 1 0 92448 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_224
timestamp 1679581782
transform 1 0 93120 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_231
timestamp 1679581782
transform 1 0 93792 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_238
timestamp 1679581782
transform 1 0 94464 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_245
timestamp 1679581782
transform 1 0 95136 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_252
timestamp 1679581782
transform 1 0 95808 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_259
timestamp 1679581782
transform 1 0 96480 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_266
timestamp 1679581782
transform 1 0 97152 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_273
timestamp 1679581782
transform 1 0 97824 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_280
timestamp 1679581782
transform 1 0 98496 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_287
timestamp 1679581782
transform 1 0 99168 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_294
timestamp 1679581782
transform 1 0 99840 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_301
timestamp 1679581782
transform 1 0 100512 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_308
timestamp 1679581782
transform 1 0 101184 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_315
timestamp 1679581782
transform 1 0 101856 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_322
timestamp 1679581782
transform 1 0 102528 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_329
timestamp 1679581782
transform 1 0 103200 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_336
timestamp 1679581782
transform 1 0 103872 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_343
timestamp 1679581782
transform 1 0 104544 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_350
timestamp 1679581782
transform 1 0 105216 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_357
timestamp 1679581782
transform 1 0 105888 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_364
timestamp 1679581782
transform 1 0 106560 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_371
timestamp 1679581782
transform 1 0 107232 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_378
timestamp 1679581782
transform 1 0 107904 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_385
timestamp 1679581782
transform 1 0 108576 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_392
timestamp 1679581782
transform 1 0 109248 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_399
timestamp 1679581782
transform 1 0 109920 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_406
timestamp 1679581782
transform 1 0 110592 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_413
timestamp 1679581782
transform 1 0 111264 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_420
timestamp 1679581782
transform 1 0 111936 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_427
timestamp 1679581782
transform 1 0 112608 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_434
timestamp 1679581782
transform 1 0 113280 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_441
timestamp 1679581782
transform 1 0 113952 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_448
timestamp 1679581782
transform 1 0 114624 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_455
timestamp 1679581782
transform 1 0 115296 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_462
timestamp 1679581782
transform 1 0 115968 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_469
timestamp 1679581782
transform 1 0 116640 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_476
timestamp 1679581782
transform 1 0 117312 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_483
timestamp 1679581782
transform 1 0 117984 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_490
timestamp 1679581782
transform 1 0 118656 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_497
timestamp 1679581782
transform 1 0 119328 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_504
timestamp 1679581782
transform 1 0 120000 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_511
timestamp 1679581782
transform 1 0 120672 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_518
timestamp 1679581782
transform 1 0 121344 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_525
timestamp 1679581782
transform 1 0 122016 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_532
timestamp 1679581782
transform 1 0 122688 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_539
timestamp 1679581782
transform 1 0 123360 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_546
timestamp 1679581782
transform 1 0 124032 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_553
timestamp 1679581782
transform 1 0 124704 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_560
timestamp 1679581782
transform 1 0 125376 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_567
timestamp 1679581782
transform 1 0 126048 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_574
timestamp 1679581782
transform 1 0 126720 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_581
timestamp 1679581782
transform 1 0 127392 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_588
timestamp 1679581782
transform 1 0 128064 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_595
timestamp 1679581782
transform 1 0 128736 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_602
timestamp 1679581782
transform 1 0 129408 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_609
timestamp 1679581782
transform 1 0 130080 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_616
timestamp 1679581782
transform 1 0 130752 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_623
timestamp 1679581782
transform 1 0 131424 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_630
timestamp 1679581782
transform 1 0 132096 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_637
timestamp 1679581782
transform 1 0 132768 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_644
timestamp 1679581782
transform 1 0 133440 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_651
timestamp 1679581782
transform 1 0 134112 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_658
timestamp 1679581782
transform 1 0 134784 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_665
timestamp 1679581782
transform 1 0 135456 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_672
timestamp 1679581782
transform 1 0 136128 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_679
timestamp 1679581782
transform 1 0 136800 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_686
timestamp 1679581782
transform 1 0 137472 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_693
timestamp 1679581782
transform 1 0 138144 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_700
timestamp 1679581782
transform 1 0 138816 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_707
timestamp 1679581782
transform 1 0 139488 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_714
timestamp 1679581782
transform 1 0 140160 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_721
timestamp 1679581782
transform 1 0 140832 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_728
timestamp 1679581782
transform 1 0 141504 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_735
timestamp 1679581782
transform 1 0 142176 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_742
timestamp 1679581782
transform 1 0 142848 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_749
timestamp 1679581782
transform 1 0 143520 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_756
timestamp 1679581782
transform 1 0 144192 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_763
timestamp 1679581782
transform 1 0 144864 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_770
timestamp 1679581782
transform 1 0 145536 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_777
timestamp 1679581782
transform 1 0 146208 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_784
timestamp 1679581782
transform 1 0 146880 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_791
timestamp 1679581782
transform 1 0 147552 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_798
timestamp 1679581782
transform 1 0 148224 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_805
timestamp 1679581782
transform 1 0 148896 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_812
timestamp 1679581782
transform 1 0 149568 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_819
timestamp 1679581782
transform 1 0 150240 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_826
timestamp 1679581782
transform 1 0 150912 0 -1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_833
timestamp 1679581782
transform 1 0 151584 0 -1 100548
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_840
timestamp 1677579658
transform 1 0 152256 0 -1 100548
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 71616 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679581782
transform 1 0 72288 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679581782
transform 1 0 72960 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679581782
transform 1 0 73632 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679581782
transform 1 0 74304 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679581782
transform 1 0 74976 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679581782
transform 1 0 75648 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679581782
transform 1 0 76320 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_56
timestamp 1679581782
transform 1 0 76992 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_63
timestamp 1679581782
transform 1 0 77664 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_70
timestamp 1679581782
transform 1 0 78336 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_77
timestamp 1679581782
transform 1 0 79008 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_84
timestamp 1679581782
transform 1 0 79680 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_91
timestamp 1679581782
transform 1 0 80352 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_98
timestamp 1679581782
transform 1 0 81024 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_105
timestamp 1679581782
transform 1 0 81696 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_112
timestamp 1679581782
transform 1 0 82368 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_119
timestamp 1679581782
transform 1 0 83040 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_126
timestamp 1679581782
transform 1 0 83712 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_133
timestamp 1679581782
transform 1 0 84384 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_140
timestamp 1679581782
transform 1 0 85056 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_147
timestamp 1679581782
transform 1 0 85728 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_154
timestamp 1679581782
transform 1 0 86400 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_161
timestamp 1679581782
transform 1 0 87072 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_168
timestamp 1679581782
transform 1 0 87744 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_175
timestamp 1679581782
transform 1 0 88416 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_182
timestamp 1679581782
transform 1 0 89088 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_189
timestamp 1679581782
transform 1 0 89760 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_196
timestamp 1679581782
transform 1 0 90432 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_203
timestamp 1679581782
transform 1 0 91104 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_210
timestamp 1679581782
transform 1 0 91776 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_217
timestamp 1679581782
transform 1 0 92448 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_224
timestamp 1679581782
transform 1 0 93120 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_231
timestamp 1679581782
transform 1 0 93792 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_238
timestamp 1679581782
transform 1 0 94464 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_245
timestamp 1679581782
transform 1 0 95136 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_252
timestamp 1679581782
transform 1 0 95808 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_259
timestamp 1679581782
transform 1 0 96480 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_266
timestamp 1679581782
transform 1 0 97152 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_273
timestamp 1679581782
transform 1 0 97824 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_280
timestamp 1679581782
transform 1 0 98496 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_287
timestamp 1679581782
transform 1 0 99168 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_294
timestamp 1679581782
transform 1 0 99840 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_301
timestamp 1679581782
transform 1 0 100512 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_308
timestamp 1679581782
transform 1 0 101184 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_315
timestamp 1679581782
transform 1 0 101856 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_322
timestamp 1679581782
transform 1 0 102528 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_329
timestamp 1679581782
transform 1 0 103200 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_336
timestamp 1679581782
transform 1 0 103872 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_343
timestamp 1679581782
transform 1 0 104544 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_350
timestamp 1679581782
transform 1 0 105216 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_357
timestamp 1679581782
transform 1 0 105888 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_364
timestamp 1679581782
transform 1 0 106560 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_371
timestamp 1679581782
transform 1 0 107232 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_378
timestamp 1679581782
transform 1 0 107904 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_385
timestamp 1679581782
transform 1 0 108576 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_392
timestamp 1679581782
transform 1 0 109248 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_399
timestamp 1679581782
transform 1 0 109920 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_406
timestamp 1679581782
transform 1 0 110592 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_413
timestamp 1679581782
transform 1 0 111264 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_420
timestamp 1679581782
transform 1 0 111936 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_427
timestamp 1679581782
transform 1 0 112608 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_434
timestamp 1679581782
transform 1 0 113280 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_441
timestamp 1679581782
transform 1 0 113952 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_448
timestamp 1679581782
transform 1 0 114624 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_455
timestamp 1679581782
transform 1 0 115296 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_462
timestamp 1679581782
transform 1 0 115968 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_469
timestamp 1679581782
transform 1 0 116640 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_476
timestamp 1679581782
transform 1 0 117312 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_483
timestamp 1679581782
transform 1 0 117984 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_490
timestamp 1679581782
transform 1 0 118656 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_497
timestamp 1679581782
transform 1 0 119328 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_504
timestamp 1679581782
transform 1 0 120000 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_511
timestamp 1679581782
transform 1 0 120672 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_518
timestamp 1679581782
transform 1 0 121344 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_525
timestamp 1679581782
transform 1 0 122016 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_532
timestamp 1679581782
transform 1 0 122688 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_539
timestamp 1679581782
transform 1 0 123360 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_546
timestamp 1679581782
transform 1 0 124032 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_553
timestamp 1679581782
transform 1 0 124704 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_560
timestamp 1679581782
transform 1 0 125376 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_567
timestamp 1679581782
transform 1 0 126048 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_574
timestamp 1679581782
transform 1 0 126720 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_581
timestamp 1679581782
transform 1 0 127392 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_588
timestamp 1679581782
transform 1 0 128064 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_595
timestamp 1679581782
transform 1 0 128736 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_602
timestamp 1679581782
transform 1 0 129408 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_609
timestamp 1679581782
transform 1 0 130080 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_616
timestamp 1679581782
transform 1 0 130752 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_623
timestamp 1679581782
transform 1 0 131424 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_630
timestamp 1679581782
transform 1 0 132096 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_637
timestamp 1679581782
transform 1 0 132768 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_644
timestamp 1679581782
transform 1 0 133440 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_651
timestamp 1679581782
transform 1 0 134112 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_658
timestamp 1679581782
transform 1 0 134784 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_665
timestamp 1679581782
transform 1 0 135456 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_672
timestamp 1679581782
transform 1 0 136128 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_679
timestamp 1679581782
transform 1 0 136800 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_686
timestamp 1679581782
transform 1 0 137472 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_693
timestamp 1679581782
transform 1 0 138144 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_700
timestamp 1679581782
transform 1 0 138816 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_707
timestamp 1679581782
transform 1 0 139488 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_714
timestamp 1679581782
transform 1 0 140160 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_721
timestamp 1679581782
transform 1 0 140832 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_728
timestamp 1679581782
transform 1 0 141504 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_735
timestamp 1679581782
transform 1 0 142176 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_742
timestamp 1679581782
transform 1 0 142848 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_749
timestamp 1679581782
transform 1 0 143520 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_756
timestamp 1679581782
transform 1 0 144192 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_763
timestamp 1679581782
transform 1 0 144864 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_770
timestamp 1679581782
transform 1 0 145536 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_777
timestamp 1679581782
transform 1 0 146208 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_784
timestamp 1679581782
transform 1 0 146880 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_791
timestamp 1679581782
transform 1 0 147552 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_798
timestamp 1679581782
transform 1 0 148224 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_805
timestamp 1679581782
transform 1 0 148896 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_812
timestamp 1679581782
transform 1 0 149568 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_819
timestamp 1679581782
transform 1 0 150240 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_826
timestamp 1679581782
transform 1 0 150912 0 1 100548
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_833
timestamp 1679581782
transform 1 0 151584 0 1 100548
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_840
timestamp 1677579658
transform 1 0 152256 0 1 100548
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679581782
transform 1 0 71616 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679581782
transform 1 0 72288 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679581782
transform 1 0 72960 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679581782
transform 1 0 73632 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_28
timestamp 1679581782
transform 1 0 74304 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_35
timestamp 1679581782
transform 1 0 74976 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_42
timestamp 1679581782
transform 1 0 75648 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_49
timestamp 1679581782
transform 1 0 76320 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_56
timestamp 1679581782
transform 1 0 76992 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_63
timestamp 1679581782
transform 1 0 77664 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_70
timestamp 1679581782
transform 1 0 78336 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_77
timestamp 1679581782
transform 1 0 79008 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_84
timestamp 1679581782
transform 1 0 79680 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_91
timestamp 1679581782
transform 1 0 80352 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_98
timestamp 1679581782
transform 1 0 81024 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_105
timestamp 1679581782
transform 1 0 81696 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_112
timestamp 1679581782
transform 1 0 82368 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_119
timestamp 1679581782
transform 1 0 83040 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_126
timestamp 1679581782
transform 1 0 83712 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_133
timestamp 1679581782
transform 1 0 84384 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_140
timestamp 1679581782
transform 1 0 85056 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_147
timestamp 1679581782
transform 1 0 85728 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_154
timestamp 1679581782
transform 1 0 86400 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_161
timestamp 1679581782
transform 1 0 87072 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_168
timestamp 1679581782
transform 1 0 87744 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_175
timestamp 1679581782
transform 1 0 88416 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_182
timestamp 1679581782
transform 1 0 89088 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_189
timestamp 1679581782
transform 1 0 89760 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_196
timestamp 1679581782
transform 1 0 90432 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_203
timestamp 1679581782
transform 1 0 91104 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_210
timestamp 1679581782
transform 1 0 91776 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_217
timestamp 1679581782
transform 1 0 92448 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_224
timestamp 1679581782
transform 1 0 93120 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_231
timestamp 1679581782
transform 1 0 93792 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_238
timestamp 1679581782
transform 1 0 94464 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_245
timestamp 1679581782
transform 1 0 95136 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_252
timestamp 1679581782
transform 1 0 95808 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_259
timestamp 1679581782
transform 1 0 96480 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_266
timestamp 1679581782
transform 1 0 97152 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_273
timestamp 1679581782
transform 1 0 97824 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_280
timestamp 1679581782
transform 1 0 98496 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_287
timestamp 1679581782
transform 1 0 99168 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_294
timestamp 1679581782
transform 1 0 99840 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_301
timestamp 1679581782
transform 1 0 100512 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_308
timestamp 1679581782
transform 1 0 101184 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_315
timestamp 1679581782
transform 1 0 101856 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_322
timestamp 1679581782
transform 1 0 102528 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_329
timestamp 1679581782
transform 1 0 103200 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_336
timestamp 1679581782
transform 1 0 103872 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_343
timestamp 1679581782
transform 1 0 104544 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_350
timestamp 1679581782
transform 1 0 105216 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_357
timestamp 1679581782
transform 1 0 105888 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_364
timestamp 1679581782
transform 1 0 106560 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_371
timestamp 1679581782
transform 1 0 107232 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_378
timestamp 1679581782
transform 1 0 107904 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_385
timestamp 1679581782
transform 1 0 108576 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_392
timestamp 1679581782
transform 1 0 109248 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_399
timestamp 1679581782
transform 1 0 109920 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_406
timestamp 1679581782
transform 1 0 110592 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_413
timestamp 1679581782
transform 1 0 111264 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_420
timestamp 1679581782
transform 1 0 111936 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_427
timestamp 1679581782
transform 1 0 112608 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_434
timestamp 1679581782
transform 1 0 113280 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_441
timestamp 1679581782
transform 1 0 113952 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_448
timestamp 1679581782
transform 1 0 114624 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_455
timestamp 1679581782
transform 1 0 115296 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_462
timestamp 1679581782
transform 1 0 115968 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_469
timestamp 1679581782
transform 1 0 116640 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_476
timestamp 1679581782
transform 1 0 117312 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_483
timestamp 1679581782
transform 1 0 117984 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_490
timestamp 1679581782
transform 1 0 118656 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_497
timestamp 1679581782
transform 1 0 119328 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_504
timestamp 1679581782
transform 1 0 120000 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_511
timestamp 1679581782
transform 1 0 120672 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_518
timestamp 1679581782
transform 1 0 121344 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_525
timestamp 1679581782
transform 1 0 122016 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_532
timestamp 1679581782
transform 1 0 122688 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_539
timestamp 1679581782
transform 1 0 123360 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_546
timestamp 1679581782
transform 1 0 124032 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_553
timestamp 1679581782
transform 1 0 124704 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_560
timestamp 1679581782
transform 1 0 125376 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_567
timestamp 1679581782
transform 1 0 126048 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_574
timestamp 1679581782
transform 1 0 126720 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_581
timestamp 1679581782
transform 1 0 127392 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_588
timestamp 1679581782
transform 1 0 128064 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_595
timestamp 1679581782
transform 1 0 128736 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_602
timestamp 1679581782
transform 1 0 129408 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_609
timestamp 1679581782
transform 1 0 130080 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_616
timestamp 1679581782
transform 1 0 130752 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_623
timestamp 1679581782
transform 1 0 131424 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_630
timestamp 1679581782
transform 1 0 132096 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_637
timestamp 1679581782
transform 1 0 132768 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_644
timestamp 1679581782
transform 1 0 133440 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_651
timestamp 1679581782
transform 1 0 134112 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_658
timestamp 1679581782
transform 1 0 134784 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_665
timestamp 1679581782
transform 1 0 135456 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_672
timestamp 1679581782
transform 1 0 136128 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_679
timestamp 1679581782
transform 1 0 136800 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_686
timestamp 1679581782
transform 1 0 137472 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_693
timestamp 1679581782
transform 1 0 138144 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_700
timestamp 1679581782
transform 1 0 138816 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_707
timestamp 1679581782
transform 1 0 139488 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_714
timestamp 1679581782
transform 1 0 140160 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_721
timestamp 1679581782
transform 1 0 140832 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_728
timestamp 1679581782
transform 1 0 141504 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_735
timestamp 1679581782
transform 1 0 142176 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_742
timestamp 1679581782
transform 1 0 142848 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_749
timestamp 1679581782
transform 1 0 143520 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_756
timestamp 1679581782
transform 1 0 144192 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_763
timestamp 1679581782
transform 1 0 144864 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_770
timestamp 1679581782
transform 1 0 145536 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_777
timestamp 1679581782
transform 1 0 146208 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_784
timestamp 1679581782
transform 1 0 146880 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_791
timestamp 1679581782
transform 1 0 147552 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_798
timestamp 1679581782
transform 1 0 148224 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_805
timestamp 1679581782
transform 1 0 148896 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_812
timestamp 1679581782
transform 1 0 149568 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_819
timestamp 1679581782
transform 1 0 150240 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_826
timestamp 1679581782
transform 1 0 150912 0 -1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_833
timestamp 1679581782
transform 1 0 151584 0 -1 102060
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_840
timestamp 1677579658
transform 1 0 152256 0 -1 102060
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679581782
transform 1 0 71616 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679581782
transform 1 0 72288 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679581782
transform 1 0 72960 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679581782
transform 1 0 73632 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_28
timestamp 1679581782
transform 1 0 74304 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_35
timestamp 1679581782
transform 1 0 74976 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_42
timestamp 1679581782
transform 1 0 75648 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_49
timestamp 1679581782
transform 1 0 76320 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_56
timestamp 1679581782
transform 1 0 76992 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_63
timestamp 1679581782
transform 1 0 77664 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_70
timestamp 1679581782
transform 1 0 78336 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_77
timestamp 1679581782
transform 1 0 79008 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_84
timestamp 1679581782
transform 1 0 79680 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_91
timestamp 1679581782
transform 1 0 80352 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_98
timestamp 1679581782
transform 1 0 81024 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_105
timestamp 1679581782
transform 1 0 81696 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_112
timestamp 1679581782
transform 1 0 82368 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_119
timestamp 1679581782
transform 1 0 83040 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_126
timestamp 1679581782
transform 1 0 83712 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_133
timestamp 1679581782
transform 1 0 84384 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_140
timestamp 1679581782
transform 1 0 85056 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_147
timestamp 1679581782
transform 1 0 85728 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_154
timestamp 1679581782
transform 1 0 86400 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_161
timestamp 1679581782
transform 1 0 87072 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_168
timestamp 1679581782
transform 1 0 87744 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_175
timestamp 1679581782
transform 1 0 88416 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_182
timestamp 1679581782
transform 1 0 89088 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_189
timestamp 1679581782
transform 1 0 89760 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_196
timestamp 1679581782
transform 1 0 90432 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_203
timestamp 1679581782
transform 1 0 91104 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_210
timestamp 1679581782
transform 1 0 91776 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_217
timestamp 1679581782
transform 1 0 92448 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_224
timestamp 1679581782
transform 1 0 93120 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_231
timestamp 1679581782
transform 1 0 93792 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_238
timestamp 1679581782
transform 1 0 94464 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_245
timestamp 1679581782
transform 1 0 95136 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_252
timestamp 1679581782
transform 1 0 95808 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_259
timestamp 1679581782
transform 1 0 96480 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_266
timestamp 1679581782
transform 1 0 97152 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_273
timestamp 1679581782
transform 1 0 97824 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_280
timestamp 1679581782
transform 1 0 98496 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_287
timestamp 1679581782
transform 1 0 99168 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_294
timestamp 1679581782
transform 1 0 99840 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_301
timestamp 1679581782
transform 1 0 100512 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_308
timestamp 1679581782
transform 1 0 101184 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_315
timestamp 1679581782
transform 1 0 101856 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_322
timestamp 1679581782
transform 1 0 102528 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_329
timestamp 1679581782
transform 1 0 103200 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_336
timestamp 1679581782
transform 1 0 103872 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_343
timestamp 1679581782
transform 1 0 104544 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_350
timestamp 1679581782
transform 1 0 105216 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_357
timestamp 1679581782
transform 1 0 105888 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_364
timestamp 1679581782
transform 1 0 106560 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_371
timestamp 1679581782
transform 1 0 107232 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_378
timestamp 1679581782
transform 1 0 107904 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_385
timestamp 1679581782
transform 1 0 108576 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_392
timestamp 1679581782
transform 1 0 109248 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_399
timestamp 1679581782
transform 1 0 109920 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_406
timestamp 1679581782
transform 1 0 110592 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_413
timestamp 1679581782
transform 1 0 111264 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_420
timestamp 1679581782
transform 1 0 111936 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_427
timestamp 1679581782
transform 1 0 112608 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_434
timestamp 1679581782
transform 1 0 113280 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_441
timestamp 1679581782
transform 1 0 113952 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_448
timestamp 1679581782
transform 1 0 114624 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_455
timestamp 1679581782
transform 1 0 115296 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_462
timestamp 1679581782
transform 1 0 115968 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_469
timestamp 1679581782
transform 1 0 116640 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_476
timestamp 1679581782
transform 1 0 117312 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_483
timestamp 1679581782
transform 1 0 117984 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_490
timestamp 1679581782
transform 1 0 118656 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_497
timestamp 1679581782
transform 1 0 119328 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_504
timestamp 1679581782
transform 1 0 120000 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_511
timestamp 1679581782
transform 1 0 120672 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_518
timestamp 1679581782
transform 1 0 121344 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_525
timestamp 1679581782
transform 1 0 122016 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_532
timestamp 1679581782
transform 1 0 122688 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_539
timestamp 1679581782
transform 1 0 123360 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_546
timestamp 1679581782
transform 1 0 124032 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_553
timestamp 1679581782
transform 1 0 124704 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_560
timestamp 1679581782
transform 1 0 125376 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_567
timestamp 1679581782
transform 1 0 126048 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_574
timestamp 1679581782
transform 1 0 126720 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_581
timestamp 1679581782
transform 1 0 127392 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_588
timestamp 1679581782
transform 1 0 128064 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_595
timestamp 1679581782
transform 1 0 128736 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_602
timestamp 1679581782
transform 1 0 129408 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_609
timestamp 1679581782
transform 1 0 130080 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_616
timestamp 1679581782
transform 1 0 130752 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_623
timestamp 1679581782
transform 1 0 131424 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_630
timestamp 1679581782
transform 1 0 132096 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_637
timestamp 1679581782
transform 1 0 132768 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_644
timestamp 1679581782
transform 1 0 133440 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_651
timestamp 1679581782
transform 1 0 134112 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_658
timestamp 1679581782
transform 1 0 134784 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_665
timestamp 1679581782
transform 1 0 135456 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_672
timestamp 1679581782
transform 1 0 136128 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_679
timestamp 1679581782
transform 1 0 136800 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_686
timestamp 1679581782
transform 1 0 137472 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_693
timestamp 1679581782
transform 1 0 138144 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_700
timestamp 1679581782
transform 1 0 138816 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_707
timestamp 1679581782
transform 1 0 139488 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_714
timestamp 1679581782
transform 1 0 140160 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_721
timestamp 1679581782
transform 1 0 140832 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_728
timestamp 1679581782
transform 1 0 141504 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_735
timestamp 1679581782
transform 1 0 142176 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_742
timestamp 1679581782
transform 1 0 142848 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_749
timestamp 1679581782
transform 1 0 143520 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_756
timestamp 1679581782
transform 1 0 144192 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_763
timestamp 1679581782
transform 1 0 144864 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_770
timestamp 1679581782
transform 1 0 145536 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_777
timestamp 1679581782
transform 1 0 146208 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_784
timestamp 1679581782
transform 1 0 146880 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_791
timestamp 1679581782
transform 1 0 147552 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_798
timestamp 1679581782
transform 1 0 148224 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_805
timestamp 1679581782
transform 1 0 148896 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_812
timestamp 1679581782
transform 1 0 149568 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_819
timestamp 1679581782
transform 1 0 150240 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_826
timestamp 1679581782
transform 1 0 150912 0 1 102060
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_833
timestamp 1679581782
transform 1 0 151584 0 1 102060
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_840
timestamp 1677579658
transform 1 0 152256 0 1 102060
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 71616 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679581782
transform 1 0 72288 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679581782
transform 1 0 72960 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679581782
transform 1 0 73632 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679581782
transform 1 0 74304 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679581782
transform 1 0 74976 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679581782
transform 1 0 75648 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679581782
transform 1 0 76320 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679581782
transform 1 0 76992 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_63
timestamp 1679581782
transform 1 0 77664 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_70
timestamp 1679581782
transform 1 0 78336 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_77
timestamp 1679581782
transform 1 0 79008 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_84
timestamp 1679581782
transform 1 0 79680 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_91
timestamp 1679581782
transform 1 0 80352 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_98
timestamp 1679581782
transform 1 0 81024 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_105
timestamp 1679581782
transform 1 0 81696 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_112
timestamp 1679581782
transform 1 0 82368 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_119
timestamp 1679581782
transform 1 0 83040 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_126
timestamp 1679581782
transform 1 0 83712 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_133
timestamp 1679581782
transform 1 0 84384 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_140
timestamp 1679581782
transform 1 0 85056 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_147
timestamp 1679581782
transform 1 0 85728 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_154
timestamp 1679581782
transform 1 0 86400 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679581782
transform 1 0 87072 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_168
timestamp 1679581782
transform 1 0 87744 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_175
timestamp 1679581782
transform 1 0 88416 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_182
timestamp 1679581782
transform 1 0 89088 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_189
timestamp 1679581782
transform 1 0 89760 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_196
timestamp 1679581782
transform 1 0 90432 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_203
timestamp 1679581782
transform 1 0 91104 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_210
timestamp 1679581782
transform 1 0 91776 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_217
timestamp 1679581782
transform 1 0 92448 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_224
timestamp 1679581782
transform 1 0 93120 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_231
timestamp 1679581782
transform 1 0 93792 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_238
timestamp 1679581782
transform 1 0 94464 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_245
timestamp 1679581782
transform 1 0 95136 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_252
timestamp 1679581782
transform 1 0 95808 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_259
timestamp 1679581782
transform 1 0 96480 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_266
timestamp 1679581782
transform 1 0 97152 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_273
timestamp 1679581782
transform 1 0 97824 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_280
timestamp 1679581782
transform 1 0 98496 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_287
timestamp 1679581782
transform 1 0 99168 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_294
timestamp 1679581782
transform 1 0 99840 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_301
timestamp 1679581782
transform 1 0 100512 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_308
timestamp 1679581782
transform 1 0 101184 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_315
timestamp 1679581782
transform 1 0 101856 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_322
timestamp 1679581782
transform 1 0 102528 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_329
timestamp 1679581782
transform 1 0 103200 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_336
timestamp 1679581782
transform 1 0 103872 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_343
timestamp 1679581782
transform 1 0 104544 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_350
timestamp 1679581782
transform 1 0 105216 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_357
timestamp 1679581782
transform 1 0 105888 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_364
timestamp 1679581782
transform 1 0 106560 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_371
timestamp 1679581782
transform 1 0 107232 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_378
timestamp 1679581782
transform 1 0 107904 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_385
timestamp 1679581782
transform 1 0 108576 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_392
timestamp 1679581782
transform 1 0 109248 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_399
timestamp 1679581782
transform 1 0 109920 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_406
timestamp 1679581782
transform 1 0 110592 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_413
timestamp 1679581782
transform 1 0 111264 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_420
timestamp 1679581782
transform 1 0 111936 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_427
timestamp 1679581782
transform 1 0 112608 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_434
timestamp 1679581782
transform 1 0 113280 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_441
timestamp 1679581782
transform 1 0 113952 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_448
timestamp 1679581782
transform 1 0 114624 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_455
timestamp 1679581782
transform 1 0 115296 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_462
timestamp 1679581782
transform 1 0 115968 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_469
timestamp 1679581782
transform 1 0 116640 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_476
timestamp 1679581782
transform 1 0 117312 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_483
timestamp 1679581782
transform 1 0 117984 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_490
timestamp 1679581782
transform 1 0 118656 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_497
timestamp 1679581782
transform 1 0 119328 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_504
timestamp 1679581782
transform 1 0 120000 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_511
timestamp 1679581782
transform 1 0 120672 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_518
timestamp 1679581782
transform 1 0 121344 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_525
timestamp 1679581782
transform 1 0 122016 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_532
timestamp 1679581782
transform 1 0 122688 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_539
timestamp 1679581782
transform 1 0 123360 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_546
timestamp 1679581782
transform 1 0 124032 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_553
timestamp 1679581782
transform 1 0 124704 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_560
timestamp 1679581782
transform 1 0 125376 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_567
timestamp 1679581782
transform 1 0 126048 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_574
timestamp 1679581782
transform 1 0 126720 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_581
timestamp 1679581782
transform 1 0 127392 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_588
timestamp 1679581782
transform 1 0 128064 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_595
timestamp 1679581782
transform 1 0 128736 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_602
timestamp 1679581782
transform 1 0 129408 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_609
timestamp 1679581782
transform 1 0 130080 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_616
timestamp 1679581782
transform 1 0 130752 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_623
timestamp 1679581782
transform 1 0 131424 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_630
timestamp 1679581782
transform 1 0 132096 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_637
timestamp 1679581782
transform 1 0 132768 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_644
timestamp 1679581782
transform 1 0 133440 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_651
timestamp 1679581782
transform 1 0 134112 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_658
timestamp 1679581782
transform 1 0 134784 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_665
timestamp 1679581782
transform 1 0 135456 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_672
timestamp 1679581782
transform 1 0 136128 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_679
timestamp 1679581782
transform 1 0 136800 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_686
timestamp 1679581782
transform 1 0 137472 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_693
timestamp 1679581782
transform 1 0 138144 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_700
timestamp 1679581782
transform 1 0 138816 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_707
timestamp 1679581782
transform 1 0 139488 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_714
timestamp 1679581782
transform 1 0 140160 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_721
timestamp 1679581782
transform 1 0 140832 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_728
timestamp 1679581782
transform 1 0 141504 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_735
timestamp 1679581782
transform 1 0 142176 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_742
timestamp 1679581782
transform 1 0 142848 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_749
timestamp 1679581782
transform 1 0 143520 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_756
timestamp 1679581782
transform 1 0 144192 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_763
timestamp 1679581782
transform 1 0 144864 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_770
timestamp 1679581782
transform 1 0 145536 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_777
timestamp 1679581782
transform 1 0 146208 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_784
timestamp 1679581782
transform 1 0 146880 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_791
timestamp 1679581782
transform 1 0 147552 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_798
timestamp 1679581782
transform 1 0 148224 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_805
timestamp 1679581782
transform 1 0 148896 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_812
timestamp 1679581782
transform 1 0 149568 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_819
timestamp 1679581782
transform 1 0 150240 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_826
timestamp 1679581782
transform 1 0 150912 0 -1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_833
timestamp 1679581782
transform 1 0 151584 0 -1 103572
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_840
timestamp 1677579658
transform 1 0 152256 0 -1 103572
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679581782
transform 1 0 71616 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679581782
transform 1 0 72288 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679581782
transform 1 0 72960 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679581782
transform 1 0 73632 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679581782
transform 1 0 74304 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679581782
transform 1 0 74976 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679581782
transform 1 0 75648 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_49
timestamp 1679581782
transform 1 0 76320 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_56
timestamp 1679581782
transform 1 0 76992 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_63
timestamp 1679581782
transform 1 0 77664 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_70
timestamp 1679581782
transform 1 0 78336 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_77
timestamp 1679581782
transform 1 0 79008 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_84
timestamp 1679581782
transform 1 0 79680 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_91
timestamp 1679581782
transform 1 0 80352 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_98
timestamp 1679581782
transform 1 0 81024 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_105
timestamp 1679581782
transform 1 0 81696 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_112
timestamp 1679581782
transform 1 0 82368 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_119
timestamp 1679581782
transform 1 0 83040 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_126
timestamp 1679581782
transform 1 0 83712 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_133
timestamp 1679581782
transform 1 0 84384 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_140
timestamp 1679581782
transform 1 0 85056 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_147
timestamp 1679581782
transform 1 0 85728 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_154
timestamp 1679581782
transform 1 0 86400 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_161
timestamp 1679581782
transform 1 0 87072 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_168
timestamp 1679581782
transform 1 0 87744 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_175
timestamp 1679581782
transform 1 0 88416 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_182
timestamp 1679581782
transform 1 0 89088 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_189
timestamp 1679581782
transform 1 0 89760 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_196
timestamp 1679581782
transform 1 0 90432 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_203
timestamp 1679581782
transform 1 0 91104 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_210
timestamp 1679581782
transform 1 0 91776 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_217
timestamp 1679581782
transform 1 0 92448 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_224
timestamp 1679581782
transform 1 0 93120 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_231
timestamp 1679581782
transform 1 0 93792 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_238
timestamp 1679581782
transform 1 0 94464 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_245
timestamp 1679581782
transform 1 0 95136 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_252
timestamp 1679581782
transform 1 0 95808 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_259
timestamp 1679581782
transform 1 0 96480 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_266
timestamp 1679581782
transform 1 0 97152 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_273
timestamp 1679581782
transform 1 0 97824 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_280
timestamp 1679581782
transform 1 0 98496 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_287
timestamp 1679581782
transform 1 0 99168 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_294
timestamp 1679581782
transform 1 0 99840 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_301
timestamp 1679581782
transform 1 0 100512 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_308
timestamp 1679581782
transform 1 0 101184 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_315
timestamp 1679581782
transform 1 0 101856 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_322
timestamp 1679581782
transform 1 0 102528 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_329
timestamp 1679581782
transform 1 0 103200 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_336
timestamp 1679581782
transform 1 0 103872 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_343
timestamp 1679581782
transform 1 0 104544 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_350
timestamp 1679581782
transform 1 0 105216 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_357
timestamp 1679581782
transform 1 0 105888 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_364
timestamp 1679581782
transform 1 0 106560 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_371
timestamp 1679581782
transform 1 0 107232 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_378
timestamp 1679581782
transform 1 0 107904 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_385
timestamp 1679581782
transform 1 0 108576 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_392
timestamp 1679581782
transform 1 0 109248 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_399
timestamp 1679581782
transform 1 0 109920 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_406
timestamp 1679581782
transform 1 0 110592 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_413
timestamp 1679581782
transform 1 0 111264 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_420
timestamp 1679581782
transform 1 0 111936 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_427
timestamp 1679581782
transform 1 0 112608 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_434
timestamp 1679581782
transform 1 0 113280 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_441
timestamp 1679581782
transform 1 0 113952 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_448
timestamp 1679581782
transform 1 0 114624 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_455
timestamp 1679581782
transform 1 0 115296 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_462
timestamp 1679581782
transform 1 0 115968 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_469
timestamp 1679581782
transform 1 0 116640 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_476
timestamp 1679581782
transform 1 0 117312 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_483
timestamp 1679581782
transform 1 0 117984 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_490
timestamp 1679581782
transform 1 0 118656 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_497
timestamp 1679581782
transform 1 0 119328 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_504
timestamp 1679581782
transform 1 0 120000 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_511
timestamp 1679581782
transform 1 0 120672 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_518
timestamp 1679581782
transform 1 0 121344 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_525
timestamp 1679581782
transform 1 0 122016 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_532
timestamp 1679581782
transform 1 0 122688 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_539
timestamp 1679581782
transform 1 0 123360 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_546
timestamp 1679581782
transform 1 0 124032 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_553
timestamp 1679581782
transform 1 0 124704 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_560
timestamp 1679581782
transform 1 0 125376 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_567
timestamp 1679581782
transform 1 0 126048 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_574
timestamp 1679581782
transform 1 0 126720 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_581
timestamp 1679581782
transform 1 0 127392 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_588
timestamp 1679581782
transform 1 0 128064 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_595
timestamp 1679581782
transform 1 0 128736 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_602
timestamp 1679581782
transform 1 0 129408 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_609
timestamp 1679581782
transform 1 0 130080 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_616
timestamp 1679581782
transform 1 0 130752 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_623
timestamp 1679581782
transform 1 0 131424 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_630
timestamp 1679581782
transform 1 0 132096 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_637
timestamp 1679581782
transform 1 0 132768 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_644
timestamp 1679581782
transform 1 0 133440 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_651
timestamp 1679581782
transform 1 0 134112 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_658
timestamp 1679581782
transform 1 0 134784 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_665
timestamp 1679581782
transform 1 0 135456 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_672
timestamp 1679581782
transform 1 0 136128 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_679
timestamp 1679581782
transform 1 0 136800 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_686
timestamp 1679581782
transform 1 0 137472 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_693
timestamp 1679581782
transform 1 0 138144 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_700
timestamp 1679581782
transform 1 0 138816 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_707
timestamp 1679581782
transform 1 0 139488 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_714
timestamp 1679581782
transform 1 0 140160 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_721
timestamp 1679581782
transform 1 0 140832 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_728
timestamp 1679581782
transform 1 0 141504 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_735
timestamp 1679581782
transform 1 0 142176 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_742
timestamp 1679581782
transform 1 0 142848 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_749
timestamp 1679581782
transform 1 0 143520 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_756
timestamp 1679581782
transform 1 0 144192 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_763
timestamp 1679581782
transform 1 0 144864 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_770
timestamp 1679581782
transform 1 0 145536 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_777
timestamp 1679581782
transform 1 0 146208 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_784
timestamp 1679581782
transform 1 0 146880 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_791
timestamp 1679581782
transform 1 0 147552 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_798
timestamp 1679581782
transform 1 0 148224 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_805
timestamp 1679581782
transform 1 0 148896 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_812
timestamp 1679581782
transform 1 0 149568 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_819
timestamp 1679581782
transform 1 0 150240 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_826
timestamp 1679581782
transform 1 0 150912 0 1 103572
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_833
timestamp 1679581782
transform 1 0 151584 0 1 103572
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_840
timestamp 1677579658
transform 1 0 152256 0 1 103572
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 71616 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679581782
transform 1 0 72288 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679581782
transform 1 0 72960 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679581782
transform 1 0 73632 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679581782
transform 1 0 74304 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679581782
transform 1 0 74976 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679581782
transform 1 0 75648 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679581782
transform 1 0 76320 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679581782
transform 1 0 76992 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679581782
transform 1 0 77664 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679581782
transform 1 0 78336 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679581782
transform 1 0 79008 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679581782
transform 1 0 79680 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679581782
transform 1 0 80352 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679581782
transform 1 0 81024 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679581782
transform 1 0 81696 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_112
timestamp 1679581782
transform 1 0 82368 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_119
timestamp 1679581782
transform 1 0 83040 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_126
timestamp 1679581782
transform 1 0 83712 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_133
timestamp 1679581782
transform 1 0 84384 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_140
timestamp 1679581782
transform 1 0 85056 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_147
timestamp 1679581782
transform 1 0 85728 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_154
timestamp 1679581782
transform 1 0 86400 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_161
timestamp 1679581782
transform 1 0 87072 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_168
timestamp 1679581782
transform 1 0 87744 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_175
timestamp 1679581782
transform 1 0 88416 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_182
timestamp 1679581782
transform 1 0 89088 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_189
timestamp 1679581782
transform 1 0 89760 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_196
timestamp 1679581782
transform 1 0 90432 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_203
timestamp 1679581782
transform 1 0 91104 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_210
timestamp 1679581782
transform 1 0 91776 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_217
timestamp 1679581782
transform 1 0 92448 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_224
timestamp 1679581782
transform 1 0 93120 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_231
timestamp 1679581782
transform 1 0 93792 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_238
timestamp 1679581782
transform 1 0 94464 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_245
timestamp 1679581782
transform 1 0 95136 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_252
timestamp 1679581782
transform 1 0 95808 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_259
timestamp 1679581782
transform 1 0 96480 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_266
timestamp 1679581782
transform 1 0 97152 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_273
timestamp 1679581782
transform 1 0 97824 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_280
timestamp 1679581782
transform 1 0 98496 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_287
timestamp 1679581782
transform 1 0 99168 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_294
timestamp 1679581782
transform 1 0 99840 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_301
timestamp 1679581782
transform 1 0 100512 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_308
timestamp 1679581782
transform 1 0 101184 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_315
timestamp 1679581782
transform 1 0 101856 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_322
timestamp 1679581782
transform 1 0 102528 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_329
timestamp 1679581782
transform 1 0 103200 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_336
timestamp 1679581782
transform 1 0 103872 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_343
timestamp 1679581782
transform 1 0 104544 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_350
timestamp 1679581782
transform 1 0 105216 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_357
timestamp 1679581782
transform 1 0 105888 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_364
timestamp 1679581782
transform 1 0 106560 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_371
timestamp 1679581782
transform 1 0 107232 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_378
timestamp 1679581782
transform 1 0 107904 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_385
timestamp 1679581782
transform 1 0 108576 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_392
timestamp 1679581782
transform 1 0 109248 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_399
timestamp 1679581782
transform 1 0 109920 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_406
timestamp 1679581782
transform 1 0 110592 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_413
timestamp 1679581782
transform 1 0 111264 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_420
timestamp 1679581782
transform 1 0 111936 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_427
timestamp 1679581782
transform 1 0 112608 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_434
timestamp 1679581782
transform 1 0 113280 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_441
timestamp 1679581782
transform 1 0 113952 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_448
timestamp 1679581782
transform 1 0 114624 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_455
timestamp 1679581782
transform 1 0 115296 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_462
timestamp 1679581782
transform 1 0 115968 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_469
timestamp 1679581782
transform 1 0 116640 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_476
timestamp 1679581782
transform 1 0 117312 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_483
timestamp 1679581782
transform 1 0 117984 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_490
timestamp 1679581782
transform 1 0 118656 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_497
timestamp 1679581782
transform 1 0 119328 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_504
timestamp 1679581782
transform 1 0 120000 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_511
timestamp 1679581782
transform 1 0 120672 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_518
timestamp 1679581782
transform 1 0 121344 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_525
timestamp 1679581782
transform 1 0 122016 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_532
timestamp 1679581782
transform 1 0 122688 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_539
timestamp 1679581782
transform 1 0 123360 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_546
timestamp 1679581782
transform 1 0 124032 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_553
timestamp 1679581782
transform 1 0 124704 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_560
timestamp 1679581782
transform 1 0 125376 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_567
timestamp 1679581782
transform 1 0 126048 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_574
timestamp 1679581782
transform 1 0 126720 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_581
timestamp 1679581782
transform 1 0 127392 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_588
timestamp 1679581782
transform 1 0 128064 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_595
timestamp 1679581782
transform 1 0 128736 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_602
timestamp 1679581782
transform 1 0 129408 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_609
timestamp 1679581782
transform 1 0 130080 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_616
timestamp 1679581782
transform 1 0 130752 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_623
timestamp 1679581782
transform 1 0 131424 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_630
timestamp 1679581782
transform 1 0 132096 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_637
timestamp 1679581782
transform 1 0 132768 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_644
timestamp 1679581782
transform 1 0 133440 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_651
timestamp 1679581782
transform 1 0 134112 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_658
timestamp 1679581782
transform 1 0 134784 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_665
timestamp 1679581782
transform 1 0 135456 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_672
timestamp 1679581782
transform 1 0 136128 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_679
timestamp 1679581782
transform 1 0 136800 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_686
timestamp 1679581782
transform 1 0 137472 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_693
timestamp 1679581782
transform 1 0 138144 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_700
timestamp 1679581782
transform 1 0 138816 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_707
timestamp 1679581782
transform 1 0 139488 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_714
timestamp 1679581782
transform 1 0 140160 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_721
timestamp 1679581782
transform 1 0 140832 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_728
timestamp 1679581782
transform 1 0 141504 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_735
timestamp 1679581782
transform 1 0 142176 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_742
timestamp 1679581782
transform 1 0 142848 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_749
timestamp 1679581782
transform 1 0 143520 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_756
timestamp 1679581782
transform 1 0 144192 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_763
timestamp 1679581782
transform 1 0 144864 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_770
timestamp 1679581782
transform 1 0 145536 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_777
timestamp 1679581782
transform 1 0 146208 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_784
timestamp 1679581782
transform 1 0 146880 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_791
timestamp 1679581782
transform 1 0 147552 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_798
timestamp 1679581782
transform 1 0 148224 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_805
timestamp 1679581782
transform 1 0 148896 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_812
timestamp 1679581782
transform 1 0 149568 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_819
timestamp 1679581782
transform 1 0 150240 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_826
timestamp 1679581782
transform 1 0 150912 0 -1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_833
timestamp 1679581782
transform 1 0 151584 0 -1 105084
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_840
timestamp 1677579658
transform 1 0 152256 0 -1 105084
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679581782
transform 1 0 71616 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679581782
transform 1 0 72288 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679581782
transform 1 0 72960 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679581782
transform 1 0 73632 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679581782
transform 1 0 74304 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679581782
transform 1 0 74976 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679581782
transform 1 0 75648 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679581782
transform 1 0 76320 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679581782
transform 1 0 76992 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_63
timestamp 1679581782
transform 1 0 77664 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_70
timestamp 1679581782
transform 1 0 78336 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_77
timestamp 1679581782
transform 1 0 79008 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_84
timestamp 1679581782
transform 1 0 79680 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_91
timestamp 1679581782
transform 1 0 80352 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_98
timestamp 1679581782
transform 1 0 81024 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_105
timestamp 1679581782
transform 1 0 81696 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_112
timestamp 1679581782
transform 1 0 82368 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_119
timestamp 1679581782
transform 1 0 83040 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_126
timestamp 1679581782
transform 1 0 83712 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_133
timestamp 1679581782
transform 1 0 84384 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_140
timestamp 1679581782
transform 1 0 85056 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_147
timestamp 1679581782
transform 1 0 85728 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_154
timestamp 1679581782
transform 1 0 86400 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_161
timestamp 1679581782
transform 1 0 87072 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_168
timestamp 1679581782
transform 1 0 87744 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_175
timestamp 1679581782
transform 1 0 88416 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_182
timestamp 1679581782
transform 1 0 89088 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_189
timestamp 1679581782
transform 1 0 89760 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_196
timestamp 1679581782
transform 1 0 90432 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_203
timestamp 1679581782
transform 1 0 91104 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_210
timestamp 1679581782
transform 1 0 91776 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_217
timestamp 1679581782
transform 1 0 92448 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_224
timestamp 1679581782
transform 1 0 93120 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_231
timestamp 1679581782
transform 1 0 93792 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_238
timestamp 1679581782
transform 1 0 94464 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_245
timestamp 1679581782
transform 1 0 95136 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_252
timestamp 1679581782
transform 1 0 95808 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_259
timestamp 1679581782
transform 1 0 96480 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_266
timestamp 1679581782
transform 1 0 97152 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_273
timestamp 1679581782
transform 1 0 97824 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_280
timestamp 1679581782
transform 1 0 98496 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_287
timestamp 1679581782
transform 1 0 99168 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_294
timestamp 1679581782
transform 1 0 99840 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_301
timestamp 1679581782
transform 1 0 100512 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_308
timestamp 1679581782
transform 1 0 101184 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_315
timestamp 1679581782
transform 1 0 101856 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_322
timestamp 1679581782
transform 1 0 102528 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_329
timestamp 1679581782
transform 1 0 103200 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_336
timestamp 1679581782
transform 1 0 103872 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_343
timestamp 1679581782
transform 1 0 104544 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_350
timestamp 1679581782
transform 1 0 105216 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_357
timestamp 1679581782
transform 1 0 105888 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_364
timestamp 1679581782
transform 1 0 106560 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_371
timestamp 1679581782
transform 1 0 107232 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_378
timestamp 1679581782
transform 1 0 107904 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_385
timestamp 1679581782
transform 1 0 108576 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_392
timestamp 1679581782
transform 1 0 109248 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_399
timestamp 1679581782
transform 1 0 109920 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_406
timestamp 1679581782
transform 1 0 110592 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_413
timestamp 1679581782
transform 1 0 111264 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_420
timestamp 1679581782
transform 1 0 111936 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_427
timestamp 1679581782
transform 1 0 112608 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_434
timestamp 1679581782
transform 1 0 113280 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_441
timestamp 1679581782
transform 1 0 113952 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_448
timestamp 1679581782
transform 1 0 114624 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_455
timestamp 1679581782
transform 1 0 115296 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_462
timestamp 1679581782
transform 1 0 115968 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_469
timestamp 1679581782
transform 1 0 116640 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_476
timestamp 1679581782
transform 1 0 117312 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_483
timestamp 1679581782
transform 1 0 117984 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_490
timestamp 1679581782
transform 1 0 118656 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_497
timestamp 1679581782
transform 1 0 119328 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_504
timestamp 1679581782
transform 1 0 120000 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_511
timestamp 1679581782
transform 1 0 120672 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_518
timestamp 1679581782
transform 1 0 121344 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_525
timestamp 1679581782
transform 1 0 122016 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_532
timestamp 1679581782
transform 1 0 122688 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_539
timestamp 1679581782
transform 1 0 123360 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_546
timestamp 1679581782
transform 1 0 124032 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_553
timestamp 1679581782
transform 1 0 124704 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_560
timestamp 1679581782
transform 1 0 125376 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_567
timestamp 1679581782
transform 1 0 126048 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_574
timestamp 1679581782
transform 1 0 126720 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_581
timestamp 1679581782
transform 1 0 127392 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_588
timestamp 1679581782
transform 1 0 128064 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_595
timestamp 1679581782
transform 1 0 128736 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_602
timestamp 1679581782
transform 1 0 129408 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_609
timestamp 1679581782
transform 1 0 130080 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_616
timestamp 1679581782
transform 1 0 130752 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_623
timestamp 1679581782
transform 1 0 131424 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_630
timestamp 1679581782
transform 1 0 132096 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_637
timestamp 1679581782
transform 1 0 132768 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_644
timestamp 1679581782
transform 1 0 133440 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_651
timestamp 1679581782
transform 1 0 134112 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_658
timestamp 1679581782
transform 1 0 134784 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_665
timestamp 1679581782
transform 1 0 135456 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_672
timestamp 1679581782
transform 1 0 136128 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_679
timestamp 1679581782
transform 1 0 136800 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_686
timestamp 1679581782
transform 1 0 137472 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_693
timestamp 1679581782
transform 1 0 138144 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_700
timestamp 1679581782
transform 1 0 138816 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_707
timestamp 1679581782
transform 1 0 139488 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_714
timestamp 1679581782
transform 1 0 140160 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_721
timestamp 1679581782
transform 1 0 140832 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_728
timestamp 1679581782
transform 1 0 141504 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_735
timestamp 1679581782
transform 1 0 142176 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_742
timestamp 1679581782
transform 1 0 142848 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_749
timestamp 1679581782
transform 1 0 143520 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_756
timestamp 1679581782
transform 1 0 144192 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_763
timestamp 1679581782
transform 1 0 144864 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_770
timestamp 1679581782
transform 1 0 145536 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_777
timestamp 1679581782
transform 1 0 146208 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_784
timestamp 1679581782
transform 1 0 146880 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_791
timestamp 1679581782
transform 1 0 147552 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_798
timestamp 1679581782
transform 1 0 148224 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_805
timestamp 1679581782
transform 1 0 148896 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_812
timestamp 1679581782
transform 1 0 149568 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_819
timestamp 1679581782
transform 1 0 150240 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_826
timestamp 1679581782
transform 1 0 150912 0 1 105084
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_833
timestamp 1679581782
transform 1 0 151584 0 1 105084
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_840
timestamp 1677579658
transform 1 0 152256 0 1 105084
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 71616 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679581782
transform 1 0 72288 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679581782
transform 1 0 72960 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679581782
transform 1 0 73632 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 74304 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 74976 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679581782
transform 1 0 75648 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679581782
transform 1 0 76320 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679581782
transform 1 0 76992 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679581782
transform 1 0 77664 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679581782
transform 1 0 78336 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679581782
transform 1 0 79008 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679581782
transform 1 0 79680 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679581782
transform 1 0 80352 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679581782
transform 1 0 81024 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679581782
transform 1 0 81696 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679581782
transform 1 0 82368 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_119
timestamp 1679581782
transform 1 0 83040 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_126
timestamp 1679581782
transform 1 0 83712 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_133
timestamp 1679581782
transform 1 0 84384 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_140
timestamp 1679581782
transform 1 0 85056 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_147
timestamp 1679581782
transform 1 0 85728 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_154
timestamp 1679581782
transform 1 0 86400 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_161
timestamp 1679581782
transform 1 0 87072 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_168
timestamp 1679581782
transform 1 0 87744 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_175
timestamp 1679581782
transform 1 0 88416 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_182
timestamp 1679581782
transform 1 0 89088 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_189
timestamp 1679581782
transform 1 0 89760 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_196
timestamp 1679581782
transform 1 0 90432 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_203
timestamp 1679581782
transform 1 0 91104 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_210
timestamp 1679581782
transform 1 0 91776 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_217
timestamp 1679581782
transform 1 0 92448 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_224
timestamp 1679581782
transform 1 0 93120 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_231
timestamp 1679581782
transform 1 0 93792 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_238
timestamp 1679581782
transform 1 0 94464 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_245
timestamp 1679581782
transform 1 0 95136 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_252
timestamp 1679581782
transform 1 0 95808 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_259
timestamp 1679581782
transform 1 0 96480 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_266
timestamp 1679581782
transform 1 0 97152 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_273
timestamp 1679581782
transform 1 0 97824 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_280
timestamp 1679581782
transform 1 0 98496 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_287
timestamp 1679581782
transform 1 0 99168 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_294
timestamp 1679581782
transform 1 0 99840 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_301
timestamp 1679581782
transform 1 0 100512 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_308
timestamp 1679581782
transform 1 0 101184 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_315
timestamp 1679581782
transform 1 0 101856 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_322
timestamp 1679581782
transform 1 0 102528 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_329
timestamp 1679581782
transform 1 0 103200 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_336
timestamp 1679581782
transform 1 0 103872 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_343
timestamp 1679581782
transform 1 0 104544 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_350
timestamp 1679581782
transform 1 0 105216 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_357
timestamp 1679581782
transform 1 0 105888 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_364
timestamp 1679581782
transform 1 0 106560 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_371
timestamp 1679581782
transform 1 0 107232 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_378
timestamp 1679581782
transform 1 0 107904 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_385
timestamp 1679581782
transform 1 0 108576 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_392
timestamp 1679581782
transform 1 0 109248 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_399
timestamp 1679581782
transform 1 0 109920 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_406
timestamp 1679581782
transform 1 0 110592 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_413
timestamp 1679581782
transform 1 0 111264 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_420
timestamp 1679581782
transform 1 0 111936 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_427
timestamp 1679581782
transform 1 0 112608 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_434
timestamp 1679581782
transform 1 0 113280 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_441
timestamp 1679581782
transform 1 0 113952 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_448
timestamp 1679581782
transform 1 0 114624 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_455
timestamp 1679581782
transform 1 0 115296 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_462
timestamp 1679581782
transform 1 0 115968 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_469
timestamp 1679581782
transform 1 0 116640 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_476
timestamp 1679581782
transform 1 0 117312 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_483
timestamp 1679581782
transform 1 0 117984 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_490
timestamp 1679581782
transform 1 0 118656 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_497
timestamp 1679581782
transform 1 0 119328 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_504
timestamp 1679581782
transform 1 0 120000 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_511
timestamp 1679581782
transform 1 0 120672 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_518
timestamp 1679581782
transform 1 0 121344 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_525
timestamp 1679581782
transform 1 0 122016 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_532
timestamp 1679581782
transform 1 0 122688 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_539
timestamp 1679581782
transform 1 0 123360 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_546
timestamp 1679581782
transform 1 0 124032 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_553
timestamp 1679581782
transform 1 0 124704 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_560
timestamp 1679581782
transform 1 0 125376 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_567
timestamp 1679581782
transform 1 0 126048 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_574
timestamp 1679581782
transform 1 0 126720 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_581
timestamp 1679581782
transform 1 0 127392 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_588
timestamp 1679581782
transform 1 0 128064 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_595
timestamp 1679581782
transform 1 0 128736 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_602
timestamp 1679581782
transform 1 0 129408 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_609
timestamp 1679581782
transform 1 0 130080 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_616
timestamp 1679581782
transform 1 0 130752 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_623
timestamp 1679581782
transform 1 0 131424 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_630
timestamp 1679581782
transform 1 0 132096 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_637
timestamp 1679581782
transform 1 0 132768 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_644
timestamp 1679581782
transform 1 0 133440 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_651
timestamp 1679581782
transform 1 0 134112 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_658
timestamp 1679581782
transform 1 0 134784 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_665
timestamp 1679581782
transform 1 0 135456 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_672
timestamp 1679581782
transform 1 0 136128 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_679
timestamp 1679581782
transform 1 0 136800 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_686
timestamp 1679581782
transform 1 0 137472 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_693
timestamp 1679581782
transform 1 0 138144 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_700
timestamp 1679581782
transform 1 0 138816 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_707
timestamp 1679581782
transform 1 0 139488 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_714
timestamp 1679581782
transform 1 0 140160 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_721
timestamp 1679581782
transform 1 0 140832 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_728
timestamp 1679581782
transform 1 0 141504 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_735
timestamp 1679581782
transform 1 0 142176 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_742
timestamp 1679581782
transform 1 0 142848 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_749
timestamp 1679581782
transform 1 0 143520 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_756
timestamp 1679581782
transform 1 0 144192 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_763
timestamp 1679581782
transform 1 0 144864 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_770
timestamp 1679581782
transform 1 0 145536 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_777
timestamp 1679581782
transform 1 0 146208 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_784
timestamp 1679581782
transform 1 0 146880 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_791
timestamp 1679581782
transform 1 0 147552 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_798
timestamp 1679581782
transform 1 0 148224 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_805
timestamp 1679581782
transform 1 0 148896 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_812
timestamp 1679581782
transform 1 0 149568 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_819
timestamp 1679581782
transform 1 0 150240 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_826
timestamp 1679581782
transform 1 0 150912 0 -1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_833
timestamp 1679581782
transform 1 0 151584 0 -1 106596
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_840
timestamp 1677579658
transform 1 0 152256 0 -1 106596
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679581782
transform 1 0 71616 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679581782
transform 1 0 72288 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679581782
transform 1 0 72960 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679581782
transform 1 0 73632 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679581782
transform 1 0 74304 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679581782
transform 1 0 74976 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679581782
transform 1 0 75648 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679581782
transform 1 0 76320 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679581782
transform 1 0 76992 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679581782
transform 1 0 77664 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679581782
transform 1 0 78336 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679581782
transform 1 0 79008 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679581782
transform 1 0 79680 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679581782
transform 1 0 80352 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679581782
transform 1 0 81024 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679581782
transform 1 0 81696 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679581782
transform 1 0 82368 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679581782
transform 1 0 83040 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679581782
transform 1 0 83712 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679581782
transform 1 0 84384 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679581782
transform 1 0 85056 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679581782
transform 1 0 85728 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679581782
transform 1 0 86400 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679581782
transform 1 0 87072 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679581782
transform 1 0 87744 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679581782
transform 1 0 88416 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_182
timestamp 1679581782
transform 1 0 89088 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_189
timestamp 1679581782
transform 1 0 89760 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_196
timestamp 1679581782
transform 1 0 90432 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679581782
transform 1 0 91104 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_210
timestamp 1679581782
transform 1 0 91776 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_217
timestamp 1679581782
transform 1 0 92448 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679581782
transform 1 0 93120 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679581782
transform 1 0 93792 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679581782
transform 1 0 94464 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679581782
transform 1 0 95136 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679581782
transform 1 0 95808 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679581782
transform 1 0 96480 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_266
timestamp 1679581782
transform 1 0 97152 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_273
timestamp 1679581782
transform 1 0 97824 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_280
timestamp 1679581782
transform 1 0 98496 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679581782
transform 1 0 99168 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679581782
transform 1 0 99840 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679581782
transform 1 0 100512 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679581782
transform 1 0 101184 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_315
timestamp 1679581782
transform 1 0 101856 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_322
timestamp 1679581782
transform 1 0 102528 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_329
timestamp 1679581782
transform 1 0 103200 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_336
timestamp 1679581782
transform 1 0 103872 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_343
timestamp 1679581782
transform 1 0 104544 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_350
timestamp 1679581782
transform 1 0 105216 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_357
timestamp 1679581782
transform 1 0 105888 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_364
timestamp 1679581782
transform 1 0 106560 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_371
timestamp 1679581782
transform 1 0 107232 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_378
timestamp 1679581782
transform 1 0 107904 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_385
timestamp 1679581782
transform 1 0 108576 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_392
timestamp 1679581782
transform 1 0 109248 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_399
timestamp 1679581782
transform 1 0 109920 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_406
timestamp 1679581782
transform 1 0 110592 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_413
timestamp 1679581782
transform 1 0 111264 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_420
timestamp 1679581782
transform 1 0 111936 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679581782
transform 1 0 112608 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679581782
transform 1 0 113280 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679581782
transform 1 0 113952 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679581782
transform 1 0 114624 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679581782
transform 1 0 115296 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679581782
transform 1 0 115968 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679581782
transform 1 0 116640 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679581782
transform 1 0 117312 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679581782
transform 1 0 117984 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679581782
transform 1 0 118656 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_497
timestamp 1679581782
transform 1 0 119328 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_504
timestamp 1679581782
transform 1 0 120000 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_511
timestamp 1679581782
transform 1 0 120672 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_518
timestamp 1679581782
transform 1 0 121344 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_525
timestamp 1679581782
transform 1 0 122016 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_532
timestamp 1679581782
transform 1 0 122688 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_539
timestamp 1679581782
transform 1 0 123360 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_546
timestamp 1679581782
transform 1 0 124032 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_553
timestamp 1679581782
transform 1 0 124704 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_560
timestamp 1679581782
transform 1 0 125376 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_567
timestamp 1679581782
transform 1 0 126048 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_574
timestamp 1679581782
transform 1 0 126720 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_581
timestamp 1679581782
transform 1 0 127392 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_588
timestamp 1679581782
transform 1 0 128064 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_595
timestamp 1679581782
transform 1 0 128736 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_602
timestamp 1679581782
transform 1 0 129408 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_609
timestamp 1679581782
transform 1 0 130080 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_616
timestamp 1679581782
transform 1 0 130752 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_623
timestamp 1679581782
transform 1 0 131424 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_630
timestamp 1679581782
transform 1 0 132096 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_637
timestamp 1679581782
transform 1 0 132768 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_644
timestamp 1679581782
transform 1 0 133440 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_651
timestamp 1679581782
transform 1 0 134112 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_658
timestamp 1679581782
transform 1 0 134784 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_665
timestamp 1679581782
transform 1 0 135456 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_672
timestamp 1679581782
transform 1 0 136128 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_679
timestamp 1679581782
transform 1 0 136800 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_686
timestamp 1679581782
transform 1 0 137472 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_693
timestamp 1679581782
transform 1 0 138144 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_700
timestamp 1679581782
transform 1 0 138816 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_707
timestamp 1679581782
transform 1 0 139488 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_714
timestamp 1679581782
transform 1 0 140160 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_721
timestamp 1679581782
transform 1 0 140832 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_728
timestamp 1679581782
transform 1 0 141504 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_735
timestamp 1679581782
transform 1 0 142176 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_742
timestamp 1679581782
transform 1 0 142848 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_749
timestamp 1679581782
transform 1 0 143520 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_756
timestamp 1679581782
transform 1 0 144192 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_763
timestamp 1679581782
transform 1 0 144864 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_770
timestamp 1679581782
transform 1 0 145536 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_777
timestamp 1679581782
transform 1 0 146208 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_784
timestamp 1679581782
transform 1 0 146880 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_791
timestamp 1679581782
transform 1 0 147552 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_798
timestamp 1679581782
transform 1 0 148224 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_805
timestamp 1679581782
transform 1 0 148896 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_812
timestamp 1679581782
transform 1 0 149568 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_819
timestamp 1679581782
transform 1 0 150240 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_826
timestamp 1679581782
transform 1 0 150912 0 1 106596
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_833
timestamp 1679581782
transform 1 0 151584 0 1 106596
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_840
timestamp 1677579658
transform 1 0 152256 0 1 106596
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679581782
transform 1 0 71616 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679581782
transform 1 0 72288 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679581782
transform 1 0 72960 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679581782
transform 1 0 73632 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679581782
transform 1 0 74304 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679581782
transform 1 0 74976 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679581782
transform 1 0 75648 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679581782
transform 1 0 76320 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679581782
transform 1 0 76992 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679581782
transform 1 0 77664 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679581782
transform 1 0 78336 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679581782
transform 1 0 79008 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679581782
transform 1 0 79680 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679581782
transform 1 0 80352 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679581782
transform 1 0 81024 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679581782
transform 1 0 81696 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679581782
transform 1 0 82368 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679581782
transform 1 0 83040 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679581782
transform 1 0 83712 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679581782
transform 1 0 84384 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 85056 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679581782
transform 1 0 85728 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679581782
transform 1 0 86400 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679581782
transform 1 0 87072 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679581782
transform 1 0 87744 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679581782
transform 1 0 88416 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679581782
transform 1 0 89088 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679581782
transform 1 0 89760 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679581782
transform 1 0 90432 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679581782
transform 1 0 91104 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679581782
transform 1 0 91776 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679581782
transform 1 0 92448 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679581782
transform 1 0 93120 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679581782
transform 1 0 93792 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679581782
transform 1 0 94464 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679581782
transform 1 0 95136 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679581782
transform 1 0 95808 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679581782
transform 1 0 96480 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679581782
transform 1 0 97152 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679581782
transform 1 0 97824 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679581782
transform 1 0 98496 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679581782
transform 1 0 99168 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679581782
transform 1 0 99840 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679581782
transform 1 0 100512 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679581782
transform 1 0 101184 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679581782
transform 1 0 101856 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679581782
transform 1 0 102528 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679581782
transform 1 0 103200 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679581782
transform 1 0 103872 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679581782
transform 1 0 104544 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679581782
transform 1 0 105216 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679581782
transform 1 0 105888 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679581782
transform 1 0 106560 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679581782
transform 1 0 107232 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679581782
transform 1 0 107904 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679581782
transform 1 0 108576 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679581782
transform 1 0 109248 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679581782
transform 1 0 109920 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679581782
transform 1 0 110592 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679581782
transform 1 0 111264 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679581782
transform 1 0 111936 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679581782
transform 1 0 112608 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679581782
transform 1 0 113280 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679581782
transform 1 0 113952 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679581782
transform 1 0 114624 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679581782
transform 1 0 115296 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679581782
transform 1 0 115968 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679581782
transform 1 0 116640 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679581782
transform 1 0 117312 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679581782
transform 1 0 117984 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679581782
transform 1 0 118656 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679581782
transform 1 0 119328 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679581782
transform 1 0 120000 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679581782
transform 1 0 120672 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679581782
transform 1 0 121344 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679581782
transform 1 0 122016 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679581782
transform 1 0 122688 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679581782
transform 1 0 123360 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679581782
transform 1 0 124032 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679581782
transform 1 0 124704 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679581782
transform 1 0 125376 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679581782
transform 1 0 126048 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679581782
transform 1 0 126720 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679581782
transform 1 0 127392 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679581782
transform 1 0 128064 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679581782
transform 1 0 128736 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679581782
transform 1 0 129408 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679581782
transform 1 0 130080 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679581782
transform 1 0 130752 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679581782
transform 1 0 131424 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679581782
transform 1 0 132096 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679581782
transform 1 0 132768 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679581782
transform 1 0 133440 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679581782
transform 1 0 134112 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679581782
transform 1 0 134784 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679581782
transform 1 0 135456 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679581782
transform 1 0 136128 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679581782
transform 1 0 136800 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679581782
transform 1 0 137472 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679581782
transform 1 0 138144 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679581782
transform 1 0 138816 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679581782
transform 1 0 139488 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679581782
transform 1 0 140160 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679581782
transform 1 0 140832 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679581782
transform 1 0 141504 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679581782
transform 1 0 142176 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679581782
transform 1 0 142848 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679581782
transform 1 0 143520 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_756
timestamp 1679581782
transform 1 0 144192 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_763
timestamp 1679581782
transform 1 0 144864 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_770
timestamp 1679581782
transform 1 0 145536 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_777
timestamp 1679581782
transform 1 0 146208 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_784
timestamp 1679581782
transform 1 0 146880 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_791
timestamp 1679581782
transform 1 0 147552 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_798
timestamp 1679581782
transform 1 0 148224 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_805
timestamp 1679581782
transform 1 0 148896 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_812
timestamp 1679581782
transform 1 0 149568 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_819
timestamp 1679581782
transform 1 0 150240 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_826
timestamp 1679581782
transform 1 0 150912 0 -1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_833
timestamp 1679581782
transform 1 0 151584 0 -1 108108
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_840
timestamp 1677579658
transform 1 0 152256 0 -1 108108
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679581782
transform 1 0 71616 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679581782
transform 1 0 72288 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679581782
transform 1 0 72960 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679581782
transform 1 0 73632 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679581782
transform 1 0 74304 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679581782
transform 1 0 74976 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679581782
transform 1 0 75648 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679581782
transform 1 0 76320 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679581782
transform 1 0 76992 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679581782
transform 1 0 77664 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679581782
transform 1 0 78336 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679581782
transform 1 0 79008 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679581782
transform 1 0 79680 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679581782
transform 1 0 80352 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679581782
transform 1 0 81024 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679581782
transform 1 0 81696 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679581782
transform 1 0 82368 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679581782
transform 1 0 83040 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679581782
transform 1 0 83712 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679581782
transform 1 0 84384 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679581782
transform 1 0 85056 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679581782
transform 1 0 85728 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679581782
transform 1 0 86400 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679581782
transform 1 0 87072 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679581782
transform 1 0 87744 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679581782
transform 1 0 88416 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679581782
transform 1 0 89088 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679581782
transform 1 0 89760 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679581782
transform 1 0 90432 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679581782
transform 1 0 91104 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679581782
transform 1 0 91776 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679581782
transform 1 0 92448 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679581782
transform 1 0 93120 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679581782
transform 1 0 93792 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679581782
transform 1 0 94464 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679581782
transform 1 0 95136 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679581782
transform 1 0 95808 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679581782
transform 1 0 96480 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679581782
transform 1 0 97152 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679581782
transform 1 0 97824 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679581782
transform 1 0 98496 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679581782
transform 1 0 99168 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679581782
transform 1 0 99840 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679581782
transform 1 0 100512 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679581782
transform 1 0 101184 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679581782
transform 1 0 101856 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679581782
transform 1 0 102528 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679581782
transform 1 0 103200 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679581782
transform 1 0 103872 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679581782
transform 1 0 104544 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679581782
transform 1 0 105216 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679581782
transform 1 0 105888 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679581782
transform 1 0 106560 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679581782
transform 1 0 107232 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679581782
transform 1 0 107904 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679581782
transform 1 0 108576 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679581782
transform 1 0 109248 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679581782
transform 1 0 109920 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679581782
transform 1 0 110592 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679581782
transform 1 0 111264 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679581782
transform 1 0 111936 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679581782
transform 1 0 112608 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679581782
transform 1 0 113280 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679581782
transform 1 0 113952 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679581782
transform 1 0 114624 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679581782
transform 1 0 115296 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679581782
transform 1 0 115968 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679581782
transform 1 0 116640 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679581782
transform 1 0 117312 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679581782
transform 1 0 117984 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679581782
transform 1 0 118656 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679581782
transform 1 0 119328 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679581782
transform 1 0 120000 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679581782
transform 1 0 120672 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679581782
transform 1 0 121344 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679581782
transform 1 0 122016 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679581782
transform 1 0 122688 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679581782
transform 1 0 123360 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679581782
transform 1 0 124032 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679581782
transform 1 0 124704 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679581782
transform 1 0 125376 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_567
timestamp 1679581782
transform 1 0 126048 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_574
timestamp 1679581782
transform 1 0 126720 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_581
timestamp 1679581782
transform 1 0 127392 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_588
timestamp 1679581782
transform 1 0 128064 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_595
timestamp 1679581782
transform 1 0 128736 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_602
timestamp 1679581782
transform 1 0 129408 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_609
timestamp 1679581782
transform 1 0 130080 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_616
timestamp 1679581782
transform 1 0 130752 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_623
timestamp 1679581782
transform 1 0 131424 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_630
timestamp 1679581782
transform 1 0 132096 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_637
timestamp 1679581782
transform 1 0 132768 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_644
timestamp 1679581782
transform 1 0 133440 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_651
timestamp 1679581782
transform 1 0 134112 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_658
timestamp 1679581782
transform 1 0 134784 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_665
timestamp 1679581782
transform 1 0 135456 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_672
timestamp 1679581782
transform 1 0 136128 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_679
timestamp 1679581782
transform 1 0 136800 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_686
timestamp 1679581782
transform 1 0 137472 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_693
timestamp 1679581782
transform 1 0 138144 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_700
timestamp 1679581782
transform 1 0 138816 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_707
timestamp 1679581782
transform 1 0 139488 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_714
timestamp 1679581782
transform 1 0 140160 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_721
timestamp 1679581782
transform 1 0 140832 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_728
timestamp 1679581782
transform 1 0 141504 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_735
timestamp 1679581782
transform 1 0 142176 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_742
timestamp 1679581782
transform 1 0 142848 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_749
timestamp 1679581782
transform 1 0 143520 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_756
timestamp 1679581782
transform 1 0 144192 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_763
timestamp 1679581782
transform 1 0 144864 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_770
timestamp 1679581782
transform 1 0 145536 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_777
timestamp 1679581782
transform 1 0 146208 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_784
timestamp 1679581782
transform 1 0 146880 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_791
timestamp 1679581782
transform 1 0 147552 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_798
timestamp 1679581782
transform 1 0 148224 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_805
timestamp 1679581782
transform 1 0 148896 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_812
timestamp 1679581782
transform 1 0 149568 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_819
timestamp 1679581782
transform 1 0 150240 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_826
timestamp 1679581782
transform 1 0 150912 0 1 108108
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_833
timestamp 1679581782
transform 1 0 151584 0 1 108108
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_840
timestamp 1677579658
transform 1 0 152256 0 1 108108
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_0
timestamp 1679581782
transform 1 0 71616 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_7
timestamp 1679581782
transform 1 0 72288 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_14
timestamp 1679581782
transform 1 0 72960 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679581782
transform 1 0 73632 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_28
timestamp 1679581782
transform 1 0 74304 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_35
timestamp 1679581782
transform 1 0 74976 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_42
timestamp 1679581782
transform 1 0 75648 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_49
timestamp 1679581782
transform 1 0 76320 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_56
timestamp 1679581782
transform 1 0 76992 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_63
timestamp 1679581782
transform 1 0 77664 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_70
timestamp 1679581782
transform 1 0 78336 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_77
timestamp 1679581782
transform 1 0 79008 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_84
timestamp 1679581782
transform 1 0 79680 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_91
timestamp 1679581782
transform 1 0 80352 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_98
timestamp 1679581782
transform 1 0 81024 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_105
timestamp 1679581782
transform 1 0 81696 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_112
timestamp 1679581782
transform 1 0 82368 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_119
timestamp 1679581782
transform 1 0 83040 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_126
timestamp 1679581782
transform 1 0 83712 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_133
timestamp 1679581782
transform 1 0 84384 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_140
timestamp 1679581782
transform 1 0 85056 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_147
timestamp 1679581782
transform 1 0 85728 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_154
timestamp 1679581782
transform 1 0 86400 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_161
timestamp 1679581782
transform 1 0 87072 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_168
timestamp 1679581782
transform 1 0 87744 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_175
timestamp 1679581782
transform 1 0 88416 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_182
timestamp 1679581782
transform 1 0 89088 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_189
timestamp 1679581782
transform 1 0 89760 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_196
timestamp 1679581782
transform 1 0 90432 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_203
timestamp 1679581782
transform 1 0 91104 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_210
timestamp 1679581782
transform 1 0 91776 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_217
timestamp 1679581782
transform 1 0 92448 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_224
timestamp 1679581782
transform 1 0 93120 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_231
timestamp 1679581782
transform 1 0 93792 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_238
timestamp 1679581782
transform 1 0 94464 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_245
timestamp 1679581782
transform 1 0 95136 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_252
timestamp 1679581782
transform 1 0 95808 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_259
timestamp 1679581782
transform 1 0 96480 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_266
timestamp 1679581782
transform 1 0 97152 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_273
timestamp 1679581782
transform 1 0 97824 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_280
timestamp 1679581782
transform 1 0 98496 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_287
timestamp 1679581782
transform 1 0 99168 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_294
timestamp 1679581782
transform 1 0 99840 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_301
timestamp 1679581782
transform 1 0 100512 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_308
timestamp 1679581782
transform 1 0 101184 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_315
timestamp 1679581782
transform 1 0 101856 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_322
timestamp 1679581782
transform 1 0 102528 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_329
timestamp 1679581782
transform 1 0 103200 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_336
timestamp 1679581782
transform 1 0 103872 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_343
timestamp 1679581782
transform 1 0 104544 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_350
timestamp 1679581782
transform 1 0 105216 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_357
timestamp 1679581782
transform 1 0 105888 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_364
timestamp 1679581782
transform 1 0 106560 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_371
timestamp 1679581782
transform 1 0 107232 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_378
timestamp 1679581782
transform 1 0 107904 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_385
timestamp 1679581782
transform 1 0 108576 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_392
timestamp 1679581782
transform 1 0 109248 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_399
timestamp 1679581782
transform 1 0 109920 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_406
timestamp 1679581782
transform 1 0 110592 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_413
timestamp 1679581782
transform 1 0 111264 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_420
timestamp 1679581782
transform 1 0 111936 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_427
timestamp 1679581782
transform 1 0 112608 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_434
timestamp 1679581782
transform 1 0 113280 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_441
timestamp 1679581782
transform 1 0 113952 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_448
timestamp 1679581782
transform 1 0 114624 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_455
timestamp 1679581782
transform 1 0 115296 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_462
timestamp 1679581782
transform 1 0 115968 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_469
timestamp 1679581782
transform 1 0 116640 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_476
timestamp 1679581782
transform 1 0 117312 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_483
timestamp 1679581782
transform 1 0 117984 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_490
timestamp 1679581782
transform 1 0 118656 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_497
timestamp 1679581782
transform 1 0 119328 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_504
timestamp 1679581782
transform 1 0 120000 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_511
timestamp 1679581782
transform 1 0 120672 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_518
timestamp 1679581782
transform 1 0 121344 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_525
timestamp 1679581782
transform 1 0 122016 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_532
timestamp 1679581782
transform 1 0 122688 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_539
timestamp 1679581782
transform 1 0 123360 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_546
timestamp 1679581782
transform 1 0 124032 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_553
timestamp 1679581782
transform 1 0 124704 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_560
timestamp 1679581782
transform 1 0 125376 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_567
timestamp 1679581782
transform 1 0 126048 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_574
timestamp 1679581782
transform 1 0 126720 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_581
timestamp 1679581782
transform 1 0 127392 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_588
timestamp 1679581782
transform 1 0 128064 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_595
timestamp 1679581782
transform 1 0 128736 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_602
timestamp 1679581782
transform 1 0 129408 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_609
timestamp 1679581782
transform 1 0 130080 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_616
timestamp 1679581782
transform 1 0 130752 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_623
timestamp 1679581782
transform 1 0 131424 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_630
timestamp 1679581782
transform 1 0 132096 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_637
timestamp 1679581782
transform 1 0 132768 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_644
timestamp 1679581782
transform 1 0 133440 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_651
timestamp 1679581782
transform 1 0 134112 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_658
timestamp 1679581782
transform 1 0 134784 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_665
timestamp 1679581782
transform 1 0 135456 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_672
timestamp 1679581782
transform 1 0 136128 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_679
timestamp 1679581782
transform 1 0 136800 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_686
timestamp 1679581782
transform 1 0 137472 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_693
timestamp 1679581782
transform 1 0 138144 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_700
timestamp 1679581782
transform 1 0 138816 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_707
timestamp 1679581782
transform 1 0 139488 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_714
timestamp 1679581782
transform 1 0 140160 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_721
timestamp 1679581782
transform 1 0 140832 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_728
timestamp 1679581782
transform 1 0 141504 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_735
timestamp 1679581782
transform 1 0 142176 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_742
timestamp 1679581782
transform 1 0 142848 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_749
timestamp 1679581782
transform 1 0 143520 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_756
timestamp 1679581782
transform 1 0 144192 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_763
timestamp 1679581782
transform 1 0 144864 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_770
timestamp 1679581782
transform 1 0 145536 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_777
timestamp 1679581782
transform 1 0 146208 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_784
timestamp 1679581782
transform 1 0 146880 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_791
timestamp 1679581782
transform 1 0 147552 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_798
timestamp 1679581782
transform 1 0 148224 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_805
timestamp 1679581782
transform 1 0 148896 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_812
timestamp 1679581782
transform 1 0 149568 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_819
timestamp 1679581782
transform 1 0 150240 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_826
timestamp 1679581782
transform 1 0 150912 0 -1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_833
timestamp 1679581782
transform 1 0 151584 0 -1 109620
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_840
timestamp 1677579658
transform 1 0 152256 0 -1 109620
box -48 -56 144 834
use sg13g2_decap_8  FILLER_50_0
timestamp 1679581782
transform 1 0 71616 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_7
timestamp 1679581782
transform 1 0 72288 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_14
timestamp 1679581782
transform 1 0 72960 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_21
timestamp 1679581782
transform 1 0 73632 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_28
timestamp 1679581782
transform 1 0 74304 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_35
timestamp 1679581782
transform 1 0 74976 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_42
timestamp 1679581782
transform 1 0 75648 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_49
timestamp 1679581782
transform 1 0 76320 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_56
timestamp 1679581782
transform 1 0 76992 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_63
timestamp 1679581782
transform 1 0 77664 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_70
timestamp 1679581782
transform 1 0 78336 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_77
timestamp 1679581782
transform 1 0 79008 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_84
timestamp 1679581782
transform 1 0 79680 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_91
timestamp 1679581782
transform 1 0 80352 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_98
timestamp 1679581782
transform 1 0 81024 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_105
timestamp 1679581782
transform 1 0 81696 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_112
timestamp 1679581782
transform 1 0 82368 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_119
timestamp 1679581782
transform 1 0 83040 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_126
timestamp 1679581782
transform 1 0 83712 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_133
timestamp 1679581782
transform 1 0 84384 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_140
timestamp 1679581782
transform 1 0 85056 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_147
timestamp 1679581782
transform 1 0 85728 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_154
timestamp 1679581782
transform 1 0 86400 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_161
timestamp 1679581782
transform 1 0 87072 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_168
timestamp 1679581782
transform 1 0 87744 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_175
timestamp 1679581782
transform 1 0 88416 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_182
timestamp 1679581782
transform 1 0 89088 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_189
timestamp 1679581782
transform 1 0 89760 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_196
timestamp 1679581782
transform 1 0 90432 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_203
timestamp 1679581782
transform 1 0 91104 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_210
timestamp 1679581782
transform 1 0 91776 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_217
timestamp 1679581782
transform 1 0 92448 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_224
timestamp 1679581782
transform 1 0 93120 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_231
timestamp 1679581782
transform 1 0 93792 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_238
timestamp 1679581782
transform 1 0 94464 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_245
timestamp 1679581782
transform 1 0 95136 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_252
timestamp 1679581782
transform 1 0 95808 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_259
timestamp 1679581782
transform 1 0 96480 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_266
timestamp 1679581782
transform 1 0 97152 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_273
timestamp 1679581782
transform 1 0 97824 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_280
timestamp 1679581782
transform 1 0 98496 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_287
timestamp 1679581782
transform 1 0 99168 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_294
timestamp 1679581782
transform 1 0 99840 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_301
timestamp 1679581782
transform 1 0 100512 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_308
timestamp 1679581782
transform 1 0 101184 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_315
timestamp 1679581782
transform 1 0 101856 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_322
timestamp 1679581782
transform 1 0 102528 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_329
timestamp 1679581782
transform 1 0 103200 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_336
timestamp 1679581782
transform 1 0 103872 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_343
timestamp 1679581782
transform 1 0 104544 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_350
timestamp 1679581782
transform 1 0 105216 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_357
timestamp 1679581782
transform 1 0 105888 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_364
timestamp 1679581782
transform 1 0 106560 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_371
timestamp 1679581782
transform 1 0 107232 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_378
timestamp 1679581782
transform 1 0 107904 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_385
timestamp 1679581782
transform 1 0 108576 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_392
timestamp 1679581782
transform 1 0 109248 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_399
timestamp 1679581782
transform 1 0 109920 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_406
timestamp 1679581782
transform 1 0 110592 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_413
timestamp 1679581782
transform 1 0 111264 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_420
timestamp 1679581782
transform 1 0 111936 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_427
timestamp 1679581782
transform 1 0 112608 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_434
timestamp 1679581782
transform 1 0 113280 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_441
timestamp 1679581782
transform 1 0 113952 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_448
timestamp 1679581782
transform 1 0 114624 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_455
timestamp 1679581782
transform 1 0 115296 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_462
timestamp 1679581782
transform 1 0 115968 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_469
timestamp 1679581782
transform 1 0 116640 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_476
timestamp 1679581782
transform 1 0 117312 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_483
timestamp 1679581782
transform 1 0 117984 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_490
timestamp 1679581782
transform 1 0 118656 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_497
timestamp 1679581782
transform 1 0 119328 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_504
timestamp 1679581782
transform 1 0 120000 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_511
timestamp 1679581782
transform 1 0 120672 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_518
timestamp 1679581782
transform 1 0 121344 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_525
timestamp 1679581782
transform 1 0 122016 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_532
timestamp 1679581782
transform 1 0 122688 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_539
timestamp 1679581782
transform 1 0 123360 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_546
timestamp 1679581782
transform 1 0 124032 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_553
timestamp 1679581782
transform 1 0 124704 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_560
timestamp 1679581782
transform 1 0 125376 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_567
timestamp 1679581782
transform 1 0 126048 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_574
timestamp 1679581782
transform 1 0 126720 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_581
timestamp 1679581782
transform 1 0 127392 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_588
timestamp 1679581782
transform 1 0 128064 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_595
timestamp 1679581782
transform 1 0 128736 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_602
timestamp 1679581782
transform 1 0 129408 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_609
timestamp 1679581782
transform 1 0 130080 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_616
timestamp 1679581782
transform 1 0 130752 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_623
timestamp 1679581782
transform 1 0 131424 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_630
timestamp 1679581782
transform 1 0 132096 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_637
timestamp 1679581782
transform 1 0 132768 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_644
timestamp 1679581782
transform 1 0 133440 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_651
timestamp 1679581782
transform 1 0 134112 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_658
timestamp 1679581782
transform 1 0 134784 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_665
timestamp 1679581782
transform 1 0 135456 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_672
timestamp 1679581782
transform 1 0 136128 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_679
timestamp 1679581782
transform 1 0 136800 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_686
timestamp 1679581782
transform 1 0 137472 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_693
timestamp 1679581782
transform 1 0 138144 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_700
timestamp 1679581782
transform 1 0 138816 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_707
timestamp 1679581782
transform 1 0 139488 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_714
timestamp 1679581782
transform 1 0 140160 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_721
timestamp 1679581782
transform 1 0 140832 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_728
timestamp 1679581782
transform 1 0 141504 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_735
timestamp 1679581782
transform 1 0 142176 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_742
timestamp 1679581782
transform 1 0 142848 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_749
timestamp 1679581782
transform 1 0 143520 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_756
timestamp 1679581782
transform 1 0 144192 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_763
timestamp 1679581782
transform 1 0 144864 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_770
timestamp 1679581782
transform 1 0 145536 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_777
timestamp 1679581782
transform 1 0 146208 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_784
timestamp 1679581782
transform 1 0 146880 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_791
timestamp 1679581782
transform 1 0 147552 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_798
timestamp 1679581782
transform 1 0 148224 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_805
timestamp 1679581782
transform 1 0 148896 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_812
timestamp 1679581782
transform 1 0 149568 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_819
timestamp 1679581782
transform 1 0 150240 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_826
timestamp 1679581782
transform 1 0 150912 0 1 109620
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_833
timestamp 1679581782
transform 1 0 151584 0 1 109620
box -48 -56 720 834
use sg13g2_fill_1  FILLER_50_840
timestamp 1677579658
transform 1 0 152256 0 1 109620
box -48 -56 144 834
use sg13g2_decap_8  FILLER_51_0
timestamp 1679581782
transform 1 0 71616 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_7
timestamp 1679581782
transform 1 0 72288 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_14
timestamp 1679581782
transform 1 0 72960 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_21
timestamp 1679581782
transform 1 0 73632 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_28
timestamp 1679581782
transform 1 0 74304 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_35
timestamp 1679581782
transform 1 0 74976 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_42
timestamp 1679581782
transform 1 0 75648 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_49
timestamp 1679581782
transform 1 0 76320 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_56
timestamp 1679581782
transform 1 0 76992 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_63
timestamp 1679581782
transform 1 0 77664 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_70
timestamp 1679581782
transform 1 0 78336 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_77
timestamp 1679581782
transform 1 0 79008 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_84
timestamp 1679581782
transform 1 0 79680 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_91
timestamp 1679581782
transform 1 0 80352 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_98
timestamp 1679581782
transform 1 0 81024 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_105
timestamp 1679581782
transform 1 0 81696 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_112
timestamp 1679581782
transform 1 0 82368 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_119
timestamp 1679581782
transform 1 0 83040 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_126
timestamp 1679581782
transform 1 0 83712 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_133
timestamp 1679581782
transform 1 0 84384 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_140
timestamp 1679581782
transform 1 0 85056 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_147
timestamp 1679581782
transform 1 0 85728 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_154
timestamp 1679581782
transform 1 0 86400 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_161
timestamp 1679581782
transform 1 0 87072 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_168
timestamp 1679581782
transform 1 0 87744 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_175
timestamp 1679581782
transform 1 0 88416 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_182
timestamp 1679581782
transform 1 0 89088 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_189
timestamp 1679581782
transform 1 0 89760 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_196
timestamp 1679581782
transform 1 0 90432 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_203
timestamp 1679581782
transform 1 0 91104 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_210
timestamp 1679581782
transform 1 0 91776 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_217
timestamp 1679581782
transform 1 0 92448 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_224
timestamp 1679581782
transform 1 0 93120 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_231
timestamp 1679581782
transform 1 0 93792 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_238
timestamp 1679581782
transform 1 0 94464 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_245
timestamp 1679581782
transform 1 0 95136 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_252
timestamp 1679581782
transform 1 0 95808 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_259
timestamp 1679581782
transform 1 0 96480 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_266
timestamp 1679581782
transform 1 0 97152 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_273
timestamp 1679581782
transform 1 0 97824 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_280
timestamp 1679581782
transform 1 0 98496 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_287
timestamp 1679581782
transform 1 0 99168 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_294
timestamp 1679581782
transform 1 0 99840 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_301
timestamp 1679581782
transform 1 0 100512 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_308
timestamp 1679581782
transform 1 0 101184 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_315
timestamp 1679581782
transform 1 0 101856 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_322
timestamp 1679581782
transform 1 0 102528 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_329
timestamp 1679581782
transform 1 0 103200 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_336
timestamp 1679581782
transform 1 0 103872 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_343
timestamp 1679581782
transform 1 0 104544 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_350
timestamp 1679581782
transform 1 0 105216 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_357
timestamp 1679581782
transform 1 0 105888 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_364
timestamp 1679581782
transform 1 0 106560 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_371
timestamp 1679581782
transform 1 0 107232 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_378
timestamp 1679581782
transform 1 0 107904 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_385
timestamp 1679581782
transform 1 0 108576 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_392
timestamp 1679581782
transform 1 0 109248 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_399
timestamp 1679581782
transform 1 0 109920 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_406
timestamp 1679581782
transform 1 0 110592 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_413
timestamp 1679581782
transform 1 0 111264 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_420
timestamp 1679581782
transform 1 0 111936 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_427
timestamp 1679581782
transform 1 0 112608 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_434
timestamp 1679581782
transform 1 0 113280 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_441
timestamp 1679581782
transform 1 0 113952 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_448
timestamp 1679581782
transform 1 0 114624 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_455
timestamp 1679581782
transform 1 0 115296 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_462
timestamp 1679581782
transform 1 0 115968 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_469
timestamp 1679581782
transform 1 0 116640 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_476
timestamp 1679581782
transform 1 0 117312 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_483
timestamp 1679581782
transform 1 0 117984 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_490
timestamp 1679581782
transform 1 0 118656 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_497
timestamp 1679581782
transform 1 0 119328 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_504
timestamp 1679581782
transform 1 0 120000 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_511
timestamp 1679581782
transform 1 0 120672 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_518
timestamp 1679581782
transform 1 0 121344 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_525
timestamp 1679581782
transform 1 0 122016 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_532
timestamp 1679581782
transform 1 0 122688 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_539
timestamp 1679581782
transform 1 0 123360 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_546
timestamp 1679581782
transform 1 0 124032 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_553
timestamp 1679581782
transform 1 0 124704 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_560
timestamp 1679581782
transform 1 0 125376 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_567
timestamp 1679581782
transform 1 0 126048 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_574
timestamp 1679581782
transform 1 0 126720 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_581
timestamp 1679581782
transform 1 0 127392 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_588
timestamp 1679581782
transform 1 0 128064 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_595
timestamp 1679581782
transform 1 0 128736 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_602
timestamp 1679581782
transform 1 0 129408 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_609
timestamp 1679581782
transform 1 0 130080 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_616
timestamp 1679581782
transform 1 0 130752 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_623
timestamp 1679581782
transform 1 0 131424 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_630
timestamp 1679581782
transform 1 0 132096 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_637
timestamp 1679581782
transform 1 0 132768 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_644
timestamp 1679581782
transform 1 0 133440 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_651
timestamp 1679581782
transform 1 0 134112 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_658
timestamp 1679581782
transform 1 0 134784 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_665
timestamp 1679581782
transform 1 0 135456 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_672
timestamp 1679581782
transform 1 0 136128 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_679
timestamp 1679581782
transform 1 0 136800 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_686
timestamp 1679581782
transform 1 0 137472 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_693
timestamp 1679581782
transform 1 0 138144 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_700
timestamp 1679581782
transform 1 0 138816 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_707
timestamp 1679581782
transform 1 0 139488 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_714
timestamp 1679581782
transform 1 0 140160 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_721
timestamp 1679581782
transform 1 0 140832 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_728
timestamp 1679581782
transform 1 0 141504 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_735
timestamp 1679581782
transform 1 0 142176 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_742
timestamp 1679581782
transform 1 0 142848 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_749
timestamp 1679581782
transform 1 0 143520 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_756
timestamp 1679581782
transform 1 0 144192 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_763
timestamp 1679581782
transform 1 0 144864 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_770
timestamp 1679581782
transform 1 0 145536 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_777
timestamp 1679581782
transform 1 0 146208 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_784
timestamp 1679581782
transform 1 0 146880 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_791
timestamp 1679581782
transform 1 0 147552 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_798
timestamp 1679581782
transform 1 0 148224 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_805
timestamp 1679581782
transform 1 0 148896 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_812
timestamp 1679581782
transform 1 0 149568 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_819
timestamp 1679581782
transform 1 0 150240 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_826
timestamp 1679581782
transform 1 0 150912 0 -1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_833
timestamp 1679581782
transform 1 0 151584 0 -1 111132
box -48 -56 720 834
use sg13g2_fill_1  FILLER_51_840
timestamp 1677579658
transform 1 0 152256 0 -1 111132
box -48 -56 144 834
use sg13g2_decap_8  FILLER_52_0
timestamp 1679581782
transform 1 0 71616 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_7
timestamp 1679581782
transform 1 0 72288 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_14
timestamp 1679581782
transform 1 0 72960 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_21
timestamp 1679581782
transform 1 0 73632 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_28
timestamp 1679581782
transform 1 0 74304 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_35
timestamp 1679581782
transform 1 0 74976 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_42
timestamp 1679581782
transform 1 0 75648 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_49
timestamp 1679581782
transform 1 0 76320 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_56
timestamp 1679581782
transform 1 0 76992 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_63
timestamp 1679581782
transform 1 0 77664 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_70
timestamp 1679581782
transform 1 0 78336 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_77
timestamp 1679581782
transform 1 0 79008 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_84
timestamp 1679581782
transform 1 0 79680 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_91
timestamp 1679581782
transform 1 0 80352 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_98
timestamp 1679581782
transform 1 0 81024 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_105
timestamp 1679581782
transform 1 0 81696 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_112
timestamp 1679581782
transform 1 0 82368 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_119
timestamp 1679581782
transform 1 0 83040 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_126
timestamp 1679581782
transform 1 0 83712 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_133
timestamp 1679581782
transform 1 0 84384 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_140
timestamp 1679581782
transform 1 0 85056 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_147
timestamp 1679581782
transform 1 0 85728 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_154
timestamp 1679581782
transform 1 0 86400 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_161
timestamp 1679581782
transform 1 0 87072 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_168
timestamp 1679581782
transform 1 0 87744 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_175
timestamp 1679581782
transform 1 0 88416 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_182
timestamp 1679581782
transform 1 0 89088 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_189
timestamp 1679581782
transform 1 0 89760 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_196
timestamp 1679581782
transform 1 0 90432 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_203
timestamp 1679581782
transform 1 0 91104 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_210
timestamp 1679581782
transform 1 0 91776 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_217
timestamp 1679581782
transform 1 0 92448 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_224
timestamp 1679581782
transform 1 0 93120 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_231
timestamp 1679581782
transform 1 0 93792 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_238
timestamp 1679581782
transform 1 0 94464 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_245
timestamp 1679581782
transform 1 0 95136 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_252
timestamp 1679581782
transform 1 0 95808 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_259
timestamp 1679581782
transform 1 0 96480 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_266
timestamp 1679581782
transform 1 0 97152 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_273
timestamp 1679581782
transform 1 0 97824 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_280
timestamp 1679581782
transform 1 0 98496 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_287
timestamp 1679581782
transform 1 0 99168 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_294
timestamp 1679581782
transform 1 0 99840 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_301
timestamp 1679581782
transform 1 0 100512 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_308
timestamp 1679581782
transform 1 0 101184 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_315
timestamp 1679581782
transform 1 0 101856 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_322
timestamp 1679581782
transform 1 0 102528 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_329
timestamp 1679581782
transform 1 0 103200 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_336
timestamp 1679581782
transform 1 0 103872 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_343
timestamp 1679581782
transform 1 0 104544 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_350
timestamp 1679581782
transform 1 0 105216 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_357
timestamp 1679581782
transform 1 0 105888 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_364
timestamp 1679581782
transform 1 0 106560 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_371
timestamp 1679581782
transform 1 0 107232 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_378
timestamp 1679581782
transform 1 0 107904 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_385
timestamp 1679581782
transform 1 0 108576 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_392
timestamp 1679581782
transform 1 0 109248 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_399
timestamp 1679581782
transform 1 0 109920 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_406
timestamp 1679581782
transform 1 0 110592 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_413
timestamp 1679581782
transform 1 0 111264 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_420
timestamp 1679581782
transform 1 0 111936 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_427
timestamp 1679581782
transform 1 0 112608 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_434
timestamp 1679581782
transform 1 0 113280 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_441
timestamp 1679581782
transform 1 0 113952 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_448
timestamp 1679581782
transform 1 0 114624 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_455
timestamp 1679581782
transform 1 0 115296 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_462
timestamp 1679581782
transform 1 0 115968 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_469
timestamp 1679581782
transform 1 0 116640 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_476
timestamp 1679581782
transform 1 0 117312 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_483
timestamp 1679581782
transform 1 0 117984 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_490
timestamp 1679581782
transform 1 0 118656 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_497
timestamp 1679581782
transform 1 0 119328 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_504
timestamp 1679581782
transform 1 0 120000 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_511
timestamp 1679581782
transform 1 0 120672 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_518
timestamp 1679581782
transform 1 0 121344 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_525
timestamp 1679581782
transform 1 0 122016 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_532
timestamp 1679581782
transform 1 0 122688 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_539
timestamp 1679581782
transform 1 0 123360 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_546
timestamp 1679581782
transform 1 0 124032 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_553
timestamp 1679581782
transform 1 0 124704 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_560
timestamp 1679581782
transform 1 0 125376 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_567
timestamp 1679581782
transform 1 0 126048 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_574
timestamp 1679581782
transform 1 0 126720 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_581
timestamp 1679581782
transform 1 0 127392 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_588
timestamp 1679581782
transform 1 0 128064 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_595
timestamp 1679581782
transform 1 0 128736 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_602
timestamp 1679581782
transform 1 0 129408 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_609
timestamp 1679581782
transform 1 0 130080 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_616
timestamp 1679581782
transform 1 0 130752 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_623
timestamp 1679581782
transform 1 0 131424 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_630
timestamp 1679581782
transform 1 0 132096 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_637
timestamp 1679581782
transform 1 0 132768 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_644
timestamp 1679581782
transform 1 0 133440 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_651
timestamp 1679581782
transform 1 0 134112 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_658
timestamp 1679581782
transform 1 0 134784 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_665
timestamp 1679581782
transform 1 0 135456 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_672
timestamp 1679581782
transform 1 0 136128 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_679
timestamp 1679581782
transform 1 0 136800 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_686
timestamp 1679581782
transform 1 0 137472 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_693
timestamp 1679581782
transform 1 0 138144 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_700
timestamp 1679581782
transform 1 0 138816 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_707
timestamp 1679581782
transform 1 0 139488 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_714
timestamp 1679581782
transform 1 0 140160 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_721
timestamp 1679581782
transform 1 0 140832 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_728
timestamp 1679581782
transform 1 0 141504 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_735
timestamp 1679581782
transform 1 0 142176 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_742
timestamp 1679581782
transform 1 0 142848 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_749
timestamp 1679581782
transform 1 0 143520 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_756
timestamp 1679581782
transform 1 0 144192 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_763
timestamp 1679581782
transform 1 0 144864 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_770
timestamp 1679581782
transform 1 0 145536 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_777
timestamp 1679581782
transform 1 0 146208 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_784
timestamp 1679581782
transform 1 0 146880 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_791
timestamp 1679581782
transform 1 0 147552 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_798
timestamp 1679581782
transform 1 0 148224 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_805
timestamp 1679581782
transform 1 0 148896 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_812
timestamp 1679581782
transform 1 0 149568 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_819
timestamp 1679581782
transform 1 0 150240 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_826
timestamp 1679581782
transform 1 0 150912 0 1 111132
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_833
timestamp 1679581782
transform 1 0 151584 0 1 111132
box -48 -56 720 834
use sg13g2_fill_1  FILLER_52_840
timestamp 1677579658
transform 1 0 152256 0 1 111132
box -48 -56 144 834
use sg13g2_decap_8  FILLER_53_0
timestamp 1679581782
transform 1 0 71616 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_7
timestamp 1679581782
transform 1 0 72288 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_14
timestamp 1679581782
transform 1 0 72960 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_21
timestamp 1679581782
transform 1 0 73632 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_28
timestamp 1679581782
transform 1 0 74304 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_35
timestamp 1679581782
transform 1 0 74976 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_42
timestamp 1679581782
transform 1 0 75648 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_49
timestamp 1679581782
transform 1 0 76320 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_56
timestamp 1679581782
transform 1 0 76992 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_63
timestamp 1679581782
transform 1 0 77664 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_70
timestamp 1679581782
transform 1 0 78336 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_77
timestamp 1679581782
transform 1 0 79008 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_84
timestamp 1679581782
transform 1 0 79680 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_91
timestamp 1679581782
transform 1 0 80352 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_98
timestamp 1679581782
transform 1 0 81024 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_105
timestamp 1679581782
transform 1 0 81696 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_112
timestamp 1679581782
transform 1 0 82368 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_119
timestamp 1679581782
transform 1 0 83040 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_126
timestamp 1679581782
transform 1 0 83712 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_133
timestamp 1679581782
transform 1 0 84384 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_140
timestamp 1679581782
transform 1 0 85056 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_147
timestamp 1679581782
transform 1 0 85728 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_154
timestamp 1679581782
transform 1 0 86400 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_161
timestamp 1679581782
transform 1 0 87072 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_168
timestamp 1679581782
transform 1 0 87744 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_175
timestamp 1679581782
transform 1 0 88416 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_182
timestamp 1679581782
transform 1 0 89088 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_189
timestamp 1679581782
transform 1 0 89760 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_196
timestamp 1679581782
transform 1 0 90432 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_203
timestamp 1679581782
transform 1 0 91104 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_210
timestamp 1679581782
transform 1 0 91776 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_217
timestamp 1679581782
transform 1 0 92448 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_224
timestamp 1679581782
transform 1 0 93120 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_231
timestamp 1679581782
transform 1 0 93792 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_238
timestamp 1679581782
transform 1 0 94464 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_245
timestamp 1679581782
transform 1 0 95136 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_252
timestamp 1679581782
transform 1 0 95808 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_259
timestamp 1679581782
transform 1 0 96480 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_266
timestamp 1679581782
transform 1 0 97152 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_273
timestamp 1679581782
transform 1 0 97824 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_280
timestamp 1679581782
transform 1 0 98496 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_287
timestamp 1679581782
transform 1 0 99168 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_294
timestamp 1679581782
transform 1 0 99840 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_301
timestamp 1679581782
transform 1 0 100512 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_308
timestamp 1679581782
transform 1 0 101184 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_315
timestamp 1679581782
transform 1 0 101856 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_322
timestamp 1679581782
transform 1 0 102528 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_329
timestamp 1679581782
transform 1 0 103200 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_336
timestamp 1679581782
transform 1 0 103872 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_343
timestamp 1679581782
transform 1 0 104544 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_350
timestamp 1679581782
transform 1 0 105216 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_357
timestamp 1679581782
transform 1 0 105888 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_364
timestamp 1679581782
transform 1 0 106560 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_371
timestamp 1679581782
transform 1 0 107232 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_378
timestamp 1679581782
transform 1 0 107904 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_385
timestamp 1679581782
transform 1 0 108576 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_392
timestamp 1679581782
transform 1 0 109248 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_399
timestamp 1679581782
transform 1 0 109920 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_406
timestamp 1679581782
transform 1 0 110592 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_413
timestamp 1679581782
transform 1 0 111264 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_420
timestamp 1679581782
transform 1 0 111936 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_427
timestamp 1679581782
transform 1 0 112608 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_434
timestamp 1679581782
transform 1 0 113280 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_441
timestamp 1679581782
transform 1 0 113952 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_448
timestamp 1679581782
transform 1 0 114624 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_455
timestamp 1679581782
transform 1 0 115296 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_462
timestamp 1679581782
transform 1 0 115968 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_469
timestamp 1679581782
transform 1 0 116640 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_476
timestamp 1679581782
transform 1 0 117312 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_483
timestamp 1679581782
transform 1 0 117984 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_490
timestamp 1679581782
transform 1 0 118656 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_497
timestamp 1679581782
transform 1 0 119328 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_504
timestamp 1679581782
transform 1 0 120000 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_511
timestamp 1679581782
transform 1 0 120672 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_518
timestamp 1679581782
transform 1 0 121344 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_525
timestamp 1679581782
transform 1 0 122016 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_532
timestamp 1679581782
transform 1 0 122688 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_539
timestamp 1679581782
transform 1 0 123360 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_546
timestamp 1679581782
transform 1 0 124032 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_553
timestamp 1679581782
transform 1 0 124704 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_560
timestamp 1679581782
transform 1 0 125376 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_567
timestamp 1679581782
transform 1 0 126048 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_574
timestamp 1679581782
transform 1 0 126720 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_581
timestamp 1679581782
transform 1 0 127392 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_588
timestamp 1679581782
transform 1 0 128064 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_595
timestamp 1679581782
transform 1 0 128736 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_602
timestamp 1679581782
transform 1 0 129408 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_609
timestamp 1679581782
transform 1 0 130080 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_616
timestamp 1679581782
transform 1 0 130752 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_623
timestamp 1679581782
transform 1 0 131424 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_630
timestamp 1679581782
transform 1 0 132096 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_637
timestamp 1679581782
transform 1 0 132768 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_644
timestamp 1679581782
transform 1 0 133440 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_651
timestamp 1679581782
transform 1 0 134112 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_658
timestamp 1679581782
transform 1 0 134784 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_665
timestamp 1679581782
transform 1 0 135456 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_672
timestamp 1679581782
transform 1 0 136128 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_679
timestamp 1679581782
transform 1 0 136800 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_686
timestamp 1679581782
transform 1 0 137472 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_693
timestamp 1679581782
transform 1 0 138144 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_700
timestamp 1679581782
transform 1 0 138816 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_707
timestamp 1679581782
transform 1 0 139488 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_714
timestamp 1679581782
transform 1 0 140160 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_721
timestamp 1679581782
transform 1 0 140832 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_728
timestamp 1679581782
transform 1 0 141504 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_735
timestamp 1679581782
transform 1 0 142176 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_742
timestamp 1679581782
transform 1 0 142848 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_749
timestamp 1679581782
transform 1 0 143520 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_756
timestamp 1679581782
transform 1 0 144192 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_763
timestamp 1679581782
transform 1 0 144864 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_770
timestamp 1679581782
transform 1 0 145536 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_777
timestamp 1679581782
transform 1 0 146208 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_784
timestamp 1679581782
transform 1 0 146880 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_791
timestamp 1679581782
transform 1 0 147552 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_798
timestamp 1679581782
transform 1 0 148224 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_805
timestamp 1679581782
transform 1 0 148896 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_812
timestamp 1679581782
transform 1 0 149568 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_819
timestamp 1679581782
transform 1 0 150240 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_826
timestamp 1679581782
transform 1 0 150912 0 -1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_833
timestamp 1679581782
transform 1 0 151584 0 -1 112644
box -48 -56 720 834
use sg13g2_fill_1  FILLER_53_840
timestamp 1677579658
transform 1 0 152256 0 -1 112644
box -48 -56 144 834
use sg13g2_decap_8  FILLER_54_0
timestamp 1679581782
transform 1 0 71616 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_7
timestamp 1679581782
transform 1 0 72288 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_14
timestamp 1679581782
transform 1 0 72960 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_21
timestamp 1679581782
transform 1 0 73632 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_28
timestamp 1679581782
transform 1 0 74304 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_35
timestamp 1679581782
transform 1 0 74976 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_42
timestamp 1679581782
transform 1 0 75648 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_49
timestamp 1679581782
transform 1 0 76320 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_56
timestamp 1679581782
transform 1 0 76992 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_63
timestamp 1679581782
transform 1 0 77664 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_70
timestamp 1679581782
transform 1 0 78336 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_77
timestamp 1679581782
transform 1 0 79008 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_84
timestamp 1679581782
transform 1 0 79680 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_91
timestamp 1679581782
transform 1 0 80352 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_98
timestamp 1679581782
transform 1 0 81024 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_105
timestamp 1679581782
transform 1 0 81696 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_112
timestamp 1679581782
transform 1 0 82368 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_119
timestamp 1679581782
transform 1 0 83040 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_126
timestamp 1679581782
transform 1 0 83712 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_133
timestamp 1679581782
transform 1 0 84384 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_140
timestamp 1679581782
transform 1 0 85056 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_147
timestamp 1679581782
transform 1 0 85728 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_154
timestamp 1679581782
transform 1 0 86400 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_161
timestamp 1679581782
transform 1 0 87072 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_168
timestamp 1679581782
transform 1 0 87744 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_175
timestamp 1679581782
transform 1 0 88416 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_182
timestamp 1679581782
transform 1 0 89088 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_189
timestamp 1679581782
transform 1 0 89760 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_196
timestamp 1679581782
transform 1 0 90432 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_203
timestamp 1679581782
transform 1 0 91104 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_210
timestamp 1679581782
transform 1 0 91776 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_217
timestamp 1679581782
transform 1 0 92448 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_224
timestamp 1679581782
transform 1 0 93120 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_231
timestamp 1679581782
transform 1 0 93792 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_238
timestamp 1679581782
transform 1 0 94464 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_245
timestamp 1679581782
transform 1 0 95136 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_252
timestamp 1679581782
transform 1 0 95808 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_259
timestamp 1679581782
transform 1 0 96480 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_266
timestamp 1679581782
transform 1 0 97152 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_273
timestamp 1679581782
transform 1 0 97824 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_280
timestamp 1679581782
transform 1 0 98496 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_287
timestamp 1679581782
transform 1 0 99168 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_294
timestamp 1679581782
transform 1 0 99840 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_301
timestamp 1679581782
transform 1 0 100512 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_308
timestamp 1679581782
transform 1 0 101184 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_315
timestamp 1679581782
transform 1 0 101856 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_322
timestamp 1679581782
transform 1 0 102528 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_329
timestamp 1679581782
transform 1 0 103200 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_336
timestamp 1679581782
transform 1 0 103872 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_343
timestamp 1679581782
transform 1 0 104544 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_350
timestamp 1679581782
transform 1 0 105216 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_357
timestamp 1679581782
transform 1 0 105888 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_364
timestamp 1679581782
transform 1 0 106560 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_371
timestamp 1679581782
transform 1 0 107232 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_378
timestamp 1679581782
transform 1 0 107904 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_385
timestamp 1679581782
transform 1 0 108576 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_392
timestamp 1679581782
transform 1 0 109248 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_399
timestamp 1679581782
transform 1 0 109920 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_406
timestamp 1679581782
transform 1 0 110592 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_413
timestamp 1679581782
transform 1 0 111264 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_420
timestamp 1679581782
transform 1 0 111936 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_427
timestamp 1679581782
transform 1 0 112608 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_434
timestamp 1679581782
transform 1 0 113280 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_441
timestamp 1679581782
transform 1 0 113952 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_448
timestamp 1679581782
transform 1 0 114624 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_455
timestamp 1679581782
transform 1 0 115296 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_462
timestamp 1679581782
transform 1 0 115968 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_469
timestamp 1679581782
transform 1 0 116640 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_476
timestamp 1679581782
transform 1 0 117312 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_483
timestamp 1679581782
transform 1 0 117984 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_490
timestamp 1679581782
transform 1 0 118656 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_497
timestamp 1679581782
transform 1 0 119328 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_504
timestamp 1679581782
transform 1 0 120000 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_511
timestamp 1679581782
transform 1 0 120672 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_518
timestamp 1679581782
transform 1 0 121344 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_525
timestamp 1679581782
transform 1 0 122016 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_532
timestamp 1679581782
transform 1 0 122688 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_539
timestamp 1679581782
transform 1 0 123360 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_546
timestamp 1679581782
transform 1 0 124032 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_553
timestamp 1679581782
transform 1 0 124704 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_560
timestamp 1679581782
transform 1 0 125376 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_567
timestamp 1679581782
transform 1 0 126048 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_574
timestamp 1679581782
transform 1 0 126720 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_581
timestamp 1679581782
transform 1 0 127392 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_588
timestamp 1679581782
transform 1 0 128064 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_595
timestamp 1679581782
transform 1 0 128736 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_602
timestamp 1679581782
transform 1 0 129408 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_609
timestamp 1679581782
transform 1 0 130080 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_616
timestamp 1679581782
transform 1 0 130752 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_623
timestamp 1679581782
transform 1 0 131424 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_630
timestamp 1679581782
transform 1 0 132096 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_637
timestamp 1679581782
transform 1 0 132768 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_644
timestamp 1679581782
transform 1 0 133440 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_651
timestamp 1679581782
transform 1 0 134112 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_658
timestamp 1679581782
transform 1 0 134784 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_665
timestamp 1679581782
transform 1 0 135456 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_672
timestamp 1679581782
transform 1 0 136128 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_679
timestamp 1679581782
transform 1 0 136800 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_686
timestamp 1679581782
transform 1 0 137472 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_693
timestamp 1679581782
transform 1 0 138144 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_700
timestamp 1679581782
transform 1 0 138816 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_707
timestamp 1679581782
transform 1 0 139488 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_714
timestamp 1679581782
transform 1 0 140160 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_721
timestamp 1679581782
transform 1 0 140832 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_728
timestamp 1679581782
transform 1 0 141504 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_735
timestamp 1679581782
transform 1 0 142176 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_742
timestamp 1679581782
transform 1 0 142848 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_749
timestamp 1679581782
transform 1 0 143520 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_756
timestamp 1679581782
transform 1 0 144192 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_763
timestamp 1679581782
transform 1 0 144864 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_770
timestamp 1679581782
transform 1 0 145536 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_777
timestamp 1679581782
transform 1 0 146208 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_784
timestamp 1679581782
transform 1 0 146880 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_791
timestamp 1679581782
transform 1 0 147552 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_798
timestamp 1679581782
transform 1 0 148224 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_805
timestamp 1679581782
transform 1 0 148896 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_812
timestamp 1679581782
transform 1 0 149568 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_819
timestamp 1679581782
transform 1 0 150240 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_826
timestamp 1679581782
transform 1 0 150912 0 1 112644
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_833
timestamp 1679581782
transform 1 0 151584 0 1 112644
box -48 -56 720 834
use sg13g2_fill_1  FILLER_54_840
timestamp 1677579658
transform 1 0 152256 0 1 112644
box -48 -56 144 834
use sg13g2_decap_8  FILLER_55_0
timestamp 1679581782
transform 1 0 71616 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_7
timestamp 1679581782
transform 1 0 72288 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_14
timestamp 1679581782
transform 1 0 72960 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_21
timestamp 1679581782
transform 1 0 73632 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_28
timestamp 1679581782
transform 1 0 74304 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_35
timestamp 1679581782
transform 1 0 74976 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_42
timestamp 1679581782
transform 1 0 75648 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_49
timestamp 1679581782
transform 1 0 76320 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_56
timestamp 1679581782
transform 1 0 76992 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_63
timestamp 1679581782
transform 1 0 77664 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_70
timestamp 1679581782
transform 1 0 78336 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_77
timestamp 1679581782
transform 1 0 79008 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_84
timestamp 1679581782
transform 1 0 79680 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_91
timestamp 1679581782
transform 1 0 80352 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_98
timestamp 1679581782
transform 1 0 81024 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_105
timestamp 1679581782
transform 1 0 81696 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_112
timestamp 1679581782
transform 1 0 82368 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_119
timestamp 1679581782
transform 1 0 83040 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_126
timestamp 1679581782
transform 1 0 83712 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_133
timestamp 1679581782
transform 1 0 84384 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_140
timestamp 1679581782
transform 1 0 85056 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_147
timestamp 1679581782
transform 1 0 85728 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_154
timestamp 1679581782
transform 1 0 86400 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_161
timestamp 1679581782
transform 1 0 87072 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_168
timestamp 1679581782
transform 1 0 87744 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_175
timestamp 1679581782
transform 1 0 88416 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_182
timestamp 1679581782
transform 1 0 89088 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_189
timestamp 1679581782
transform 1 0 89760 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_196
timestamp 1679581782
transform 1 0 90432 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_203
timestamp 1679581782
transform 1 0 91104 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_210
timestamp 1679581782
transform 1 0 91776 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_217
timestamp 1679581782
transform 1 0 92448 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_224
timestamp 1679581782
transform 1 0 93120 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_231
timestamp 1679581782
transform 1 0 93792 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_238
timestamp 1679581782
transform 1 0 94464 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_245
timestamp 1679581782
transform 1 0 95136 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_252
timestamp 1679581782
transform 1 0 95808 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_259
timestamp 1679581782
transform 1 0 96480 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_266
timestamp 1679581782
transform 1 0 97152 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_273
timestamp 1679581782
transform 1 0 97824 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_280
timestamp 1679581782
transform 1 0 98496 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_287
timestamp 1679581782
transform 1 0 99168 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_294
timestamp 1679581782
transform 1 0 99840 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_301
timestamp 1679581782
transform 1 0 100512 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_308
timestamp 1679581782
transform 1 0 101184 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_315
timestamp 1679581782
transform 1 0 101856 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_322
timestamp 1679581782
transform 1 0 102528 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_329
timestamp 1679581782
transform 1 0 103200 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_336
timestamp 1679581782
transform 1 0 103872 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_343
timestamp 1679581782
transform 1 0 104544 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_350
timestamp 1679581782
transform 1 0 105216 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_357
timestamp 1679581782
transform 1 0 105888 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_364
timestamp 1679581782
transform 1 0 106560 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_371
timestamp 1679581782
transform 1 0 107232 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_378
timestamp 1679581782
transform 1 0 107904 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_385
timestamp 1679581782
transform 1 0 108576 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_392
timestamp 1679581782
transform 1 0 109248 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_399
timestamp 1679581782
transform 1 0 109920 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_406
timestamp 1679581782
transform 1 0 110592 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_413
timestamp 1679581782
transform 1 0 111264 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_420
timestamp 1679581782
transform 1 0 111936 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_427
timestamp 1679581782
transform 1 0 112608 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_434
timestamp 1679581782
transform 1 0 113280 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_441
timestamp 1679581782
transform 1 0 113952 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_448
timestamp 1679581782
transform 1 0 114624 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_455
timestamp 1679581782
transform 1 0 115296 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_462
timestamp 1679581782
transform 1 0 115968 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_469
timestamp 1679581782
transform 1 0 116640 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_476
timestamp 1679581782
transform 1 0 117312 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_483
timestamp 1679581782
transform 1 0 117984 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_490
timestamp 1679581782
transform 1 0 118656 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_497
timestamp 1679581782
transform 1 0 119328 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_504
timestamp 1679581782
transform 1 0 120000 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_511
timestamp 1679581782
transform 1 0 120672 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_518
timestamp 1679581782
transform 1 0 121344 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_525
timestamp 1679581782
transform 1 0 122016 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_532
timestamp 1679581782
transform 1 0 122688 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_539
timestamp 1679581782
transform 1 0 123360 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_546
timestamp 1679581782
transform 1 0 124032 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_553
timestamp 1679581782
transform 1 0 124704 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_560
timestamp 1679581782
transform 1 0 125376 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_567
timestamp 1679581782
transform 1 0 126048 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_574
timestamp 1679581782
transform 1 0 126720 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_581
timestamp 1679581782
transform 1 0 127392 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_588
timestamp 1679581782
transform 1 0 128064 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_595
timestamp 1679581782
transform 1 0 128736 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_602
timestamp 1679581782
transform 1 0 129408 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_609
timestamp 1679581782
transform 1 0 130080 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_616
timestamp 1679581782
transform 1 0 130752 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_623
timestamp 1679581782
transform 1 0 131424 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_630
timestamp 1679581782
transform 1 0 132096 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_637
timestamp 1679581782
transform 1 0 132768 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_644
timestamp 1679581782
transform 1 0 133440 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_651
timestamp 1679581782
transform 1 0 134112 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_658
timestamp 1679581782
transform 1 0 134784 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_665
timestamp 1679581782
transform 1 0 135456 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_672
timestamp 1679581782
transform 1 0 136128 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_679
timestamp 1679581782
transform 1 0 136800 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_686
timestamp 1679581782
transform 1 0 137472 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_693
timestamp 1679581782
transform 1 0 138144 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_700
timestamp 1679581782
transform 1 0 138816 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_707
timestamp 1679581782
transform 1 0 139488 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_714
timestamp 1679581782
transform 1 0 140160 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_721
timestamp 1679581782
transform 1 0 140832 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_728
timestamp 1679581782
transform 1 0 141504 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_735
timestamp 1679581782
transform 1 0 142176 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_742
timestamp 1679581782
transform 1 0 142848 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_749
timestamp 1679581782
transform 1 0 143520 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_756
timestamp 1679581782
transform 1 0 144192 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_763
timestamp 1679581782
transform 1 0 144864 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_770
timestamp 1679581782
transform 1 0 145536 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_777
timestamp 1679581782
transform 1 0 146208 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_784
timestamp 1679581782
transform 1 0 146880 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_791
timestamp 1679581782
transform 1 0 147552 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_798
timestamp 1679581782
transform 1 0 148224 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_805
timestamp 1679581782
transform 1 0 148896 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_812
timestamp 1679581782
transform 1 0 149568 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_819
timestamp 1679581782
transform 1 0 150240 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_826
timestamp 1679581782
transform 1 0 150912 0 -1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_833
timestamp 1679581782
transform 1 0 151584 0 -1 114156
box -48 -56 720 834
use sg13g2_fill_1  FILLER_55_840
timestamp 1677579658
transform 1 0 152256 0 -1 114156
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_0
timestamp 1679581782
transform 1 0 71616 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_7
timestamp 1679581782
transform 1 0 72288 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_14
timestamp 1679581782
transform 1 0 72960 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_21
timestamp 1679581782
transform 1 0 73632 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_28
timestamp 1679581782
transform 1 0 74304 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_35
timestamp 1679581782
transform 1 0 74976 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_42
timestamp 1679581782
transform 1 0 75648 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_49
timestamp 1679581782
transform 1 0 76320 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_56
timestamp 1679581782
transform 1 0 76992 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_63
timestamp 1679581782
transform 1 0 77664 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_70
timestamp 1679581782
transform 1 0 78336 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_77
timestamp 1679581782
transform 1 0 79008 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_84
timestamp 1679581782
transform 1 0 79680 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_91
timestamp 1679581782
transform 1 0 80352 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_98
timestamp 1679581782
transform 1 0 81024 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_105
timestamp 1679581782
transform 1 0 81696 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_112
timestamp 1679581782
transform 1 0 82368 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_119
timestamp 1679581782
transform 1 0 83040 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_126
timestamp 1679581782
transform 1 0 83712 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_133
timestamp 1679581782
transform 1 0 84384 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_140
timestamp 1679581782
transform 1 0 85056 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_147
timestamp 1679581782
transform 1 0 85728 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_154
timestamp 1679581782
transform 1 0 86400 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_161
timestamp 1679581782
transform 1 0 87072 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_168
timestamp 1679581782
transform 1 0 87744 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_175
timestamp 1679581782
transform 1 0 88416 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_182
timestamp 1679581782
transform 1 0 89088 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_189
timestamp 1679581782
transform 1 0 89760 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_196
timestamp 1679581782
transform 1 0 90432 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_203
timestamp 1679581782
transform 1 0 91104 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_210
timestamp 1679581782
transform 1 0 91776 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_217
timestamp 1679581782
transform 1 0 92448 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_224
timestamp 1679581782
transform 1 0 93120 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_231
timestamp 1679581782
transform 1 0 93792 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_238
timestamp 1679581782
transform 1 0 94464 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_245
timestamp 1679581782
transform 1 0 95136 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_252
timestamp 1679581782
transform 1 0 95808 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_259
timestamp 1679581782
transform 1 0 96480 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_266
timestamp 1679581782
transform 1 0 97152 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_273
timestamp 1679581782
transform 1 0 97824 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_280
timestamp 1679581782
transform 1 0 98496 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_287
timestamp 1679581782
transform 1 0 99168 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_294
timestamp 1679581782
transform 1 0 99840 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_301
timestamp 1679581782
transform 1 0 100512 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_308
timestamp 1679581782
transform 1 0 101184 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_315
timestamp 1679581782
transform 1 0 101856 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_322
timestamp 1679581782
transform 1 0 102528 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_329
timestamp 1679581782
transform 1 0 103200 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_336
timestamp 1679581782
transform 1 0 103872 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_343
timestamp 1679581782
transform 1 0 104544 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_350
timestamp 1679581782
transform 1 0 105216 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_357
timestamp 1679581782
transform 1 0 105888 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_364
timestamp 1679581782
transform 1 0 106560 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_371
timestamp 1679581782
transform 1 0 107232 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_378
timestamp 1679581782
transform 1 0 107904 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_385
timestamp 1679581782
transform 1 0 108576 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_392
timestamp 1679581782
transform 1 0 109248 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_399
timestamp 1679581782
transform 1 0 109920 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_406
timestamp 1679581782
transform 1 0 110592 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_413
timestamp 1679581782
transform 1 0 111264 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_420
timestamp 1679581782
transform 1 0 111936 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_427
timestamp 1679581782
transform 1 0 112608 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_434
timestamp 1679581782
transform 1 0 113280 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_441
timestamp 1679581782
transform 1 0 113952 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_448
timestamp 1679581782
transform 1 0 114624 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_455
timestamp 1679581782
transform 1 0 115296 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_462
timestamp 1679581782
transform 1 0 115968 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_469
timestamp 1679581782
transform 1 0 116640 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_476
timestamp 1679581782
transform 1 0 117312 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_483
timestamp 1679581782
transform 1 0 117984 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_490
timestamp 1679581782
transform 1 0 118656 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_497
timestamp 1679581782
transform 1 0 119328 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_504
timestamp 1679581782
transform 1 0 120000 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_511
timestamp 1679581782
transform 1 0 120672 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_518
timestamp 1679581782
transform 1 0 121344 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_525
timestamp 1679581782
transform 1 0 122016 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_532
timestamp 1679581782
transform 1 0 122688 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_539
timestamp 1679581782
transform 1 0 123360 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_546
timestamp 1679581782
transform 1 0 124032 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_553
timestamp 1679581782
transform 1 0 124704 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_560
timestamp 1679581782
transform 1 0 125376 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_567
timestamp 1679581782
transform 1 0 126048 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_574
timestamp 1679581782
transform 1 0 126720 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_581
timestamp 1679581782
transform 1 0 127392 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_588
timestamp 1679581782
transform 1 0 128064 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_595
timestamp 1679581782
transform 1 0 128736 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_602
timestamp 1679581782
transform 1 0 129408 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_609
timestamp 1679581782
transform 1 0 130080 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_616
timestamp 1679581782
transform 1 0 130752 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_623
timestamp 1679581782
transform 1 0 131424 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_630
timestamp 1679581782
transform 1 0 132096 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_637
timestamp 1679581782
transform 1 0 132768 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_644
timestamp 1679581782
transform 1 0 133440 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_651
timestamp 1679581782
transform 1 0 134112 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_658
timestamp 1679581782
transform 1 0 134784 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_665
timestamp 1679581782
transform 1 0 135456 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_672
timestamp 1679581782
transform 1 0 136128 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_679
timestamp 1679581782
transform 1 0 136800 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_686
timestamp 1679581782
transform 1 0 137472 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_693
timestamp 1679581782
transform 1 0 138144 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_700
timestamp 1679581782
transform 1 0 138816 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_707
timestamp 1679581782
transform 1 0 139488 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_714
timestamp 1679581782
transform 1 0 140160 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_721
timestamp 1679581782
transform 1 0 140832 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_728
timestamp 1679581782
transform 1 0 141504 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_735
timestamp 1679581782
transform 1 0 142176 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_742
timestamp 1679581782
transform 1 0 142848 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_749
timestamp 1679581782
transform 1 0 143520 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_756
timestamp 1679581782
transform 1 0 144192 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_763
timestamp 1679581782
transform 1 0 144864 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_770
timestamp 1679581782
transform 1 0 145536 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_777
timestamp 1679581782
transform 1 0 146208 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_784
timestamp 1679581782
transform 1 0 146880 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_791
timestamp 1679581782
transform 1 0 147552 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_798
timestamp 1679581782
transform 1 0 148224 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_805
timestamp 1679581782
transform 1 0 148896 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_812
timestamp 1679581782
transform 1 0 149568 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_819
timestamp 1679581782
transform 1 0 150240 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_826
timestamp 1679581782
transform 1 0 150912 0 1 114156
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_833
timestamp 1679581782
transform 1 0 151584 0 1 114156
box -48 -56 720 834
use sg13g2_fill_1  FILLER_56_840
timestamp 1677579658
transform 1 0 152256 0 1 114156
box -48 -56 144 834
use sg13g2_decap_8  FILLER_57_0
timestamp 1679581782
transform 1 0 71616 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_7
timestamp 1679581782
transform 1 0 72288 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_14
timestamp 1679581782
transform 1 0 72960 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_21
timestamp 1679581782
transform 1 0 73632 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_28
timestamp 1679581782
transform 1 0 74304 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_35
timestamp 1679581782
transform 1 0 74976 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_42
timestamp 1679581782
transform 1 0 75648 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_49
timestamp 1679581782
transform 1 0 76320 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_56
timestamp 1679581782
transform 1 0 76992 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_63
timestamp 1679581782
transform 1 0 77664 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_70
timestamp 1679581782
transform 1 0 78336 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_77
timestamp 1679581782
transform 1 0 79008 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_84
timestamp 1679581782
transform 1 0 79680 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_91
timestamp 1679581782
transform 1 0 80352 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_98
timestamp 1679581782
transform 1 0 81024 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_105
timestamp 1679581782
transform 1 0 81696 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_112
timestamp 1679581782
transform 1 0 82368 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_119
timestamp 1679581782
transform 1 0 83040 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_126
timestamp 1679581782
transform 1 0 83712 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_133
timestamp 1679581782
transform 1 0 84384 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_140
timestamp 1679581782
transform 1 0 85056 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_147
timestamp 1679581782
transform 1 0 85728 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_154
timestamp 1679581782
transform 1 0 86400 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_161
timestamp 1679581782
transform 1 0 87072 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_168
timestamp 1679581782
transform 1 0 87744 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_175
timestamp 1679581782
transform 1 0 88416 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_182
timestamp 1679581782
transform 1 0 89088 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_189
timestamp 1679581782
transform 1 0 89760 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_196
timestamp 1679581782
transform 1 0 90432 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_203
timestamp 1679581782
transform 1 0 91104 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_210
timestamp 1679581782
transform 1 0 91776 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_217
timestamp 1679581782
transform 1 0 92448 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_224
timestamp 1679581782
transform 1 0 93120 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_231
timestamp 1679581782
transform 1 0 93792 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_238
timestamp 1679581782
transform 1 0 94464 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_245
timestamp 1679581782
transform 1 0 95136 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_252
timestamp 1679581782
transform 1 0 95808 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_259
timestamp 1679581782
transform 1 0 96480 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_266
timestamp 1679581782
transform 1 0 97152 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_273
timestamp 1679581782
transform 1 0 97824 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_280
timestamp 1679581782
transform 1 0 98496 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_287
timestamp 1679581782
transform 1 0 99168 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_294
timestamp 1679581782
transform 1 0 99840 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_301
timestamp 1679581782
transform 1 0 100512 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_308
timestamp 1679581782
transform 1 0 101184 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_315
timestamp 1679581782
transform 1 0 101856 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_322
timestamp 1679581782
transform 1 0 102528 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_329
timestamp 1679581782
transform 1 0 103200 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_336
timestamp 1679581782
transform 1 0 103872 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_343
timestamp 1679581782
transform 1 0 104544 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_350
timestamp 1679581782
transform 1 0 105216 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_357
timestamp 1679581782
transform 1 0 105888 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_364
timestamp 1679581782
transform 1 0 106560 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_371
timestamp 1679581782
transform 1 0 107232 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_378
timestamp 1679581782
transform 1 0 107904 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_385
timestamp 1679581782
transform 1 0 108576 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_392
timestamp 1679581782
transform 1 0 109248 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_399
timestamp 1679581782
transform 1 0 109920 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_406
timestamp 1679581782
transform 1 0 110592 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_413
timestamp 1679581782
transform 1 0 111264 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_420
timestamp 1679581782
transform 1 0 111936 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_427
timestamp 1679581782
transform 1 0 112608 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_434
timestamp 1679581782
transform 1 0 113280 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_441
timestamp 1679581782
transform 1 0 113952 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_448
timestamp 1679581782
transform 1 0 114624 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_455
timestamp 1679581782
transform 1 0 115296 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_462
timestamp 1679581782
transform 1 0 115968 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_469
timestamp 1679581782
transform 1 0 116640 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_476
timestamp 1679581782
transform 1 0 117312 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_483
timestamp 1679581782
transform 1 0 117984 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_490
timestamp 1679581782
transform 1 0 118656 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_497
timestamp 1679581782
transform 1 0 119328 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_504
timestamp 1679581782
transform 1 0 120000 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_511
timestamp 1679581782
transform 1 0 120672 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_518
timestamp 1679581782
transform 1 0 121344 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_525
timestamp 1679581782
transform 1 0 122016 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_532
timestamp 1679581782
transform 1 0 122688 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_539
timestamp 1679581782
transform 1 0 123360 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_546
timestamp 1679581782
transform 1 0 124032 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_553
timestamp 1679581782
transform 1 0 124704 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_560
timestamp 1679581782
transform 1 0 125376 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_567
timestamp 1679581782
transform 1 0 126048 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_574
timestamp 1679581782
transform 1 0 126720 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_581
timestamp 1679581782
transform 1 0 127392 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_588
timestamp 1679581782
transform 1 0 128064 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_595
timestamp 1679581782
transform 1 0 128736 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_602
timestamp 1679581782
transform 1 0 129408 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_609
timestamp 1679581782
transform 1 0 130080 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_616
timestamp 1679581782
transform 1 0 130752 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_623
timestamp 1679581782
transform 1 0 131424 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_630
timestamp 1679581782
transform 1 0 132096 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_637
timestamp 1679581782
transform 1 0 132768 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_644
timestamp 1679581782
transform 1 0 133440 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_651
timestamp 1679581782
transform 1 0 134112 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_658
timestamp 1679581782
transform 1 0 134784 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_665
timestamp 1679581782
transform 1 0 135456 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_672
timestamp 1679581782
transform 1 0 136128 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_679
timestamp 1679581782
transform 1 0 136800 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_686
timestamp 1679581782
transform 1 0 137472 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_693
timestamp 1679581782
transform 1 0 138144 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_700
timestamp 1679581782
transform 1 0 138816 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_707
timestamp 1679581782
transform 1 0 139488 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_714
timestamp 1679581782
transform 1 0 140160 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_721
timestamp 1679581782
transform 1 0 140832 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_728
timestamp 1679581782
transform 1 0 141504 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_735
timestamp 1679581782
transform 1 0 142176 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_742
timestamp 1679581782
transform 1 0 142848 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_749
timestamp 1679581782
transform 1 0 143520 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_756
timestamp 1679581782
transform 1 0 144192 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_763
timestamp 1679581782
transform 1 0 144864 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_770
timestamp 1679581782
transform 1 0 145536 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_777
timestamp 1679581782
transform 1 0 146208 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_784
timestamp 1679581782
transform 1 0 146880 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_791
timestamp 1679581782
transform 1 0 147552 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_798
timestamp 1679581782
transform 1 0 148224 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_805
timestamp 1679581782
transform 1 0 148896 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_812
timestamp 1679581782
transform 1 0 149568 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_819
timestamp 1679581782
transform 1 0 150240 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_826
timestamp 1679581782
transform 1 0 150912 0 -1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_833
timestamp 1679581782
transform 1 0 151584 0 -1 115668
box -48 -56 720 834
use sg13g2_fill_1  FILLER_57_840
timestamp 1677579658
transform 1 0 152256 0 -1 115668
box -48 -56 144 834
use sg13g2_decap_8  FILLER_58_0
timestamp 1679581782
transform 1 0 71616 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_7
timestamp 1679581782
transform 1 0 72288 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_14
timestamp 1679581782
transform 1 0 72960 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_21
timestamp 1679581782
transform 1 0 73632 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_28
timestamp 1679581782
transform 1 0 74304 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_35
timestamp 1679581782
transform 1 0 74976 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_42
timestamp 1679581782
transform 1 0 75648 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_49
timestamp 1679581782
transform 1 0 76320 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_56
timestamp 1679581782
transform 1 0 76992 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_63
timestamp 1679581782
transform 1 0 77664 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_70
timestamp 1679581782
transform 1 0 78336 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_77
timestamp 1679581782
transform 1 0 79008 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_84
timestamp 1679581782
transform 1 0 79680 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_91
timestamp 1679581782
transform 1 0 80352 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_98
timestamp 1679581782
transform 1 0 81024 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_105
timestamp 1679581782
transform 1 0 81696 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_112
timestamp 1679581782
transform 1 0 82368 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_119
timestamp 1679581782
transform 1 0 83040 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_126
timestamp 1679581782
transform 1 0 83712 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_133
timestamp 1679581782
transform 1 0 84384 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_140
timestamp 1679581782
transform 1 0 85056 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_147
timestamp 1679581782
transform 1 0 85728 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_154
timestamp 1679581782
transform 1 0 86400 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_161
timestamp 1679581782
transform 1 0 87072 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_168
timestamp 1679581782
transform 1 0 87744 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_175
timestamp 1679581782
transform 1 0 88416 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_182
timestamp 1679581782
transform 1 0 89088 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_189
timestamp 1679581782
transform 1 0 89760 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_196
timestamp 1679581782
transform 1 0 90432 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_203
timestamp 1679581782
transform 1 0 91104 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_210
timestamp 1679581782
transform 1 0 91776 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_217
timestamp 1679581782
transform 1 0 92448 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_224
timestamp 1679581782
transform 1 0 93120 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_231
timestamp 1679581782
transform 1 0 93792 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_238
timestamp 1679581782
transform 1 0 94464 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_245
timestamp 1679581782
transform 1 0 95136 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_252
timestamp 1679581782
transform 1 0 95808 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_259
timestamp 1679581782
transform 1 0 96480 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_266
timestamp 1679581782
transform 1 0 97152 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_273
timestamp 1679581782
transform 1 0 97824 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_280
timestamp 1679581782
transform 1 0 98496 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_287
timestamp 1679581782
transform 1 0 99168 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_294
timestamp 1679581782
transform 1 0 99840 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_301
timestamp 1679581782
transform 1 0 100512 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_308
timestamp 1679581782
transform 1 0 101184 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_315
timestamp 1679581782
transform 1 0 101856 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_322
timestamp 1679581782
transform 1 0 102528 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_329
timestamp 1679581782
transform 1 0 103200 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_336
timestamp 1679581782
transform 1 0 103872 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_343
timestamp 1679581782
transform 1 0 104544 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_350
timestamp 1679581782
transform 1 0 105216 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_357
timestamp 1679581782
transform 1 0 105888 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_364
timestamp 1679581782
transform 1 0 106560 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_371
timestamp 1679581782
transform 1 0 107232 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_378
timestamp 1679581782
transform 1 0 107904 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_385
timestamp 1679581782
transform 1 0 108576 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_392
timestamp 1679581782
transform 1 0 109248 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_399
timestamp 1679581782
transform 1 0 109920 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_406
timestamp 1679581782
transform 1 0 110592 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_413
timestamp 1679581782
transform 1 0 111264 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_420
timestamp 1679581782
transform 1 0 111936 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_427
timestamp 1679581782
transform 1 0 112608 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_434
timestamp 1679581782
transform 1 0 113280 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_441
timestamp 1679581782
transform 1 0 113952 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_448
timestamp 1679581782
transform 1 0 114624 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_455
timestamp 1679581782
transform 1 0 115296 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_462
timestamp 1679581782
transform 1 0 115968 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_469
timestamp 1679581782
transform 1 0 116640 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_476
timestamp 1679581782
transform 1 0 117312 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_483
timestamp 1679581782
transform 1 0 117984 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_490
timestamp 1679581782
transform 1 0 118656 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_497
timestamp 1679581782
transform 1 0 119328 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_504
timestamp 1679581782
transform 1 0 120000 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_511
timestamp 1679581782
transform 1 0 120672 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_518
timestamp 1679581782
transform 1 0 121344 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_525
timestamp 1679581782
transform 1 0 122016 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_532
timestamp 1679581782
transform 1 0 122688 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_539
timestamp 1679581782
transform 1 0 123360 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_546
timestamp 1679581782
transform 1 0 124032 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_553
timestamp 1679581782
transform 1 0 124704 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_560
timestamp 1679581782
transform 1 0 125376 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_567
timestamp 1679581782
transform 1 0 126048 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_574
timestamp 1679581782
transform 1 0 126720 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_581
timestamp 1679581782
transform 1 0 127392 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_588
timestamp 1679581782
transform 1 0 128064 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_595
timestamp 1679581782
transform 1 0 128736 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_602
timestamp 1679581782
transform 1 0 129408 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_609
timestamp 1679581782
transform 1 0 130080 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_616
timestamp 1679581782
transform 1 0 130752 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_623
timestamp 1679581782
transform 1 0 131424 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_630
timestamp 1679581782
transform 1 0 132096 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_637
timestamp 1679581782
transform 1 0 132768 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_644
timestamp 1679581782
transform 1 0 133440 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_651
timestamp 1679581782
transform 1 0 134112 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_658
timestamp 1679581782
transform 1 0 134784 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_665
timestamp 1679581782
transform 1 0 135456 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_672
timestamp 1679581782
transform 1 0 136128 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_679
timestamp 1679581782
transform 1 0 136800 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_686
timestamp 1679581782
transform 1 0 137472 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_693
timestamp 1679581782
transform 1 0 138144 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_700
timestamp 1679581782
transform 1 0 138816 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_707
timestamp 1679581782
transform 1 0 139488 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_714
timestamp 1679581782
transform 1 0 140160 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_721
timestamp 1679581782
transform 1 0 140832 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_728
timestamp 1679581782
transform 1 0 141504 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_735
timestamp 1679581782
transform 1 0 142176 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_742
timestamp 1679581782
transform 1 0 142848 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_749
timestamp 1679581782
transform 1 0 143520 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_756
timestamp 1679581782
transform 1 0 144192 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_763
timestamp 1679581782
transform 1 0 144864 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_770
timestamp 1679581782
transform 1 0 145536 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_777
timestamp 1679581782
transform 1 0 146208 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_784
timestamp 1679581782
transform 1 0 146880 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_791
timestamp 1679581782
transform 1 0 147552 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_798
timestamp 1679581782
transform 1 0 148224 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_805
timestamp 1679581782
transform 1 0 148896 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_812
timestamp 1679581782
transform 1 0 149568 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_819
timestamp 1679581782
transform 1 0 150240 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_826
timestamp 1679581782
transform 1 0 150912 0 1 115668
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_833
timestamp 1679581782
transform 1 0 151584 0 1 115668
box -48 -56 720 834
use sg13g2_fill_1  FILLER_58_840
timestamp 1677579658
transform 1 0 152256 0 1 115668
box -48 -56 144 834
use sg13g2_decap_8  FILLER_59_0
timestamp 1679581782
transform 1 0 71616 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_7
timestamp 1679581782
transform 1 0 72288 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_14
timestamp 1679581782
transform 1 0 72960 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_21
timestamp 1679581782
transform 1 0 73632 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_28
timestamp 1679581782
transform 1 0 74304 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_35
timestamp 1679581782
transform 1 0 74976 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_42
timestamp 1679581782
transform 1 0 75648 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_49
timestamp 1679581782
transform 1 0 76320 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_56
timestamp 1679581782
transform 1 0 76992 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_63
timestamp 1679581782
transform 1 0 77664 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_70
timestamp 1679581782
transform 1 0 78336 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_77
timestamp 1679581782
transform 1 0 79008 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_84
timestamp 1679581782
transform 1 0 79680 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_91
timestamp 1679581782
transform 1 0 80352 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_98
timestamp 1679581782
transform 1 0 81024 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_105
timestamp 1679581782
transform 1 0 81696 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_112
timestamp 1679581782
transform 1 0 82368 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_119
timestamp 1679581782
transform 1 0 83040 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_126
timestamp 1679581782
transform 1 0 83712 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_133
timestamp 1679581782
transform 1 0 84384 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_140
timestamp 1679581782
transform 1 0 85056 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_147
timestamp 1679581782
transform 1 0 85728 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_154
timestamp 1679581782
transform 1 0 86400 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_161
timestamp 1679581782
transform 1 0 87072 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_168
timestamp 1679581782
transform 1 0 87744 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_175
timestamp 1679581782
transform 1 0 88416 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_182
timestamp 1679581782
transform 1 0 89088 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_189
timestamp 1679581782
transform 1 0 89760 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_196
timestamp 1679581782
transform 1 0 90432 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_203
timestamp 1679581782
transform 1 0 91104 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_210
timestamp 1679581782
transform 1 0 91776 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_217
timestamp 1679581782
transform 1 0 92448 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_224
timestamp 1679581782
transform 1 0 93120 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_231
timestamp 1679581782
transform 1 0 93792 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_238
timestamp 1679581782
transform 1 0 94464 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_245
timestamp 1679581782
transform 1 0 95136 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_252
timestamp 1679581782
transform 1 0 95808 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_259
timestamp 1679581782
transform 1 0 96480 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_266
timestamp 1679581782
transform 1 0 97152 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_273
timestamp 1679581782
transform 1 0 97824 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_280
timestamp 1679581782
transform 1 0 98496 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_287
timestamp 1679581782
transform 1 0 99168 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_294
timestamp 1679581782
transform 1 0 99840 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_301
timestamp 1679581782
transform 1 0 100512 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_308
timestamp 1679581782
transform 1 0 101184 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_315
timestamp 1679581782
transform 1 0 101856 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_322
timestamp 1679581782
transform 1 0 102528 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_329
timestamp 1679581782
transform 1 0 103200 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_336
timestamp 1679581782
transform 1 0 103872 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_343
timestamp 1679581782
transform 1 0 104544 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_350
timestamp 1679581782
transform 1 0 105216 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_357
timestamp 1679581782
transform 1 0 105888 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_364
timestamp 1679581782
transform 1 0 106560 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_371
timestamp 1679581782
transform 1 0 107232 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_378
timestamp 1679581782
transform 1 0 107904 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_385
timestamp 1679581782
transform 1 0 108576 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_392
timestamp 1679581782
transform 1 0 109248 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_399
timestamp 1679581782
transform 1 0 109920 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_406
timestamp 1679581782
transform 1 0 110592 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_413
timestamp 1679581782
transform 1 0 111264 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_420
timestamp 1679581782
transform 1 0 111936 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_427
timestamp 1679581782
transform 1 0 112608 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_434
timestamp 1679581782
transform 1 0 113280 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_441
timestamp 1679581782
transform 1 0 113952 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_448
timestamp 1679581782
transform 1 0 114624 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_455
timestamp 1679581782
transform 1 0 115296 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_462
timestamp 1679581782
transform 1 0 115968 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_469
timestamp 1679581782
transform 1 0 116640 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_476
timestamp 1679581782
transform 1 0 117312 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_483
timestamp 1679581782
transform 1 0 117984 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_490
timestamp 1679581782
transform 1 0 118656 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_497
timestamp 1679581782
transform 1 0 119328 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_504
timestamp 1679581782
transform 1 0 120000 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_511
timestamp 1679581782
transform 1 0 120672 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_518
timestamp 1679581782
transform 1 0 121344 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_525
timestamp 1679581782
transform 1 0 122016 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_532
timestamp 1679581782
transform 1 0 122688 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_539
timestamp 1679581782
transform 1 0 123360 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_546
timestamp 1679581782
transform 1 0 124032 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_553
timestamp 1679581782
transform 1 0 124704 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_560
timestamp 1679581782
transform 1 0 125376 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_567
timestamp 1679581782
transform 1 0 126048 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_574
timestamp 1679581782
transform 1 0 126720 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_581
timestamp 1679581782
transform 1 0 127392 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_588
timestamp 1679581782
transform 1 0 128064 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_595
timestamp 1679581782
transform 1 0 128736 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_602
timestamp 1679581782
transform 1 0 129408 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_609
timestamp 1679581782
transform 1 0 130080 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_616
timestamp 1679581782
transform 1 0 130752 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_623
timestamp 1679581782
transform 1 0 131424 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_630
timestamp 1679581782
transform 1 0 132096 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_637
timestamp 1679581782
transform 1 0 132768 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_644
timestamp 1679581782
transform 1 0 133440 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_651
timestamp 1679581782
transform 1 0 134112 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_658
timestamp 1679581782
transform 1 0 134784 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_665
timestamp 1679581782
transform 1 0 135456 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_672
timestamp 1679581782
transform 1 0 136128 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_679
timestamp 1679581782
transform 1 0 136800 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_686
timestamp 1679581782
transform 1 0 137472 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_693
timestamp 1679581782
transform 1 0 138144 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_700
timestamp 1679581782
transform 1 0 138816 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_707
timestamp 1679581782
transform 1 0 139488 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_714
timestamp 1679581782
transform 1 0 140160 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_721
timestamp 1679581782
transform 1 0 140832 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_728
timestamp 1679581782
transform 1 0 141504 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_735
timestamp 1679581782
transform 1 0 142176 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_742
timestamp 1679581782
transform 1 0 142848 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_749
timestamp 1679581782
transform 1 0 143520 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_756
timestamp 1679581782
transform 1 0 144192 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_763
timestamp 1679581782
transform 1 0 144864 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_770
timestamp 1679581782
transform 1 0 145536 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_777
timestamp 1679581782
transform 1 0 146208 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_784
timestamp 1679581782
transform 1 0 146880 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_791
timestamp 1679581782
transform 1 0 147552 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_798
timestamp 1679581782
transform 1 0 148224 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_805
timestamp 1679581782
transform 1 0 148896 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_812
timestamp 1679581782
transform 1 0 149568 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_819
timestamp 1679581782
transform 1 0 150240 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_826
timestamp 1679581782
transform 1 0 150912 0 -1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_833
timestamp 1679581782
transform 1 0 151584 0 -1 117180
box -48 -56 720 834
use sg13g2_fill_1  FILLER_59_840
timestamp 1677579658
transform 1 0 152256 0 -1 117180
box -48 -56 144 834
use sg13g2_decap_8  FILLER_60_0
timestamp 1679581782
transform 1 0 71616 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_7
timestamp 1679581782
transform 1 0 72288 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_14
timestamp 1679581782
transform 1 0 72960 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_21
timestamp 1679581782
transform 1 0 73632 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_28
timestamp 1679581782
transform 1 0 74304 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_35
timestamp 1679581782
transform 1 0 74976 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_42
timestamp 1679581782
transform 1 0 75648 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_49
timestamp 1679581782
transform 1 0 76320 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_56
timestamp 1679581782
transform 1 0 76992 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_63
timestamp 1679581782
transform 1 0 77664 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_70
timestamp 1679581782
transform 1 0 78336 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_77
timestamp 1679581782
transform 1 0 79008 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_84
timestamp 1679581782
transform 1 0 79680 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_91
timestamp 1679581782
transform 1 0 80352 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_98
timestamp 1679581782
transform 1 0 81024 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_105
timestamp 1679581782
transform 1 0 81696 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_112
timestamp 1679581782
transform 1 0 82368 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_119
timestamp 1679581782
transform 1 0 83040 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_126
timestamp 1679581782
transform 1 0 83712 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_133
timestamp 1679581782
transform 1 0 84384 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_140
timestamp 1679581782
transform 1 0 85056 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_147
timestamp 1679581782
transform 1 0 85728 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_154
timestamp 1679581782
transform 1 0 86400 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_161
timestamp 1679581782
transform 1 0 87072 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_168
timestamp 1679581782
transform 1 0 87744 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_175
timestamp 1679581782
transform 1 0 88416 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_182
timestamp 1679581782
transform 1 0 89088 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_189
timestamp 1679581782
transform 1 0 89760 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_196
timestamp 1679581782
transform 1 0 90432 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_203
timestamp 1679581782
transform 1 0 91104 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_210
timestamp 1679581782
transform 1 0 91776 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_217
timestamp 1679581782
transform 1 0 92448 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_224
timestamp 1679581782
transform 1 0 93120 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_231
timestamp 1679581782
transform 1 0 93792 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_238
timestamp 1679581782
transform 1 0 94464 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_245
timestamp 1679581782
transform 1 0 95136 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_252
timestamp 1679581782
transform 1 0 95808 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_259
timestamp 1679581782
transform 1 0 96480 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_266
timestamp 1679581782
transform 1 0 97152 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_273
timestamp 1679581782
transform 1 0 97824 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_280
timestamp 1679581782
transform 1 0 98496 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_287
timestamp 1679581782
transform 1 0 99168 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_294
timestamp 1679581782
transform 1 0 99840 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_301
timestamp 1679581782
transform 1 0 100512 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_308
timestamp 1679581782
transform 1 0 101184 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_315
timestamp 1679581782
transform 1 0 101856 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_322
timestamp 1679581782
transform 1 0 102528 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_329
timestamp 1679581782
transform 1 0 103200 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_336
timestamp 1679581782
transform 1 0 103872 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_343
timestamp 1679581782
transform 1 0 104544 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_350
timestamp 1679581782
transform 1 0 105216 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_357
timestamp 1679581782
transform 1 0 105888 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_364
timestamp 1679581782
transform 1 0 106560 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_371
timestamp 1679581782
transform 1 0 107232 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_378
timestamp 1679581782
transform 1 0 107904 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_385
timestamp 1679581782
transform 1 0 108576 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_392
timestamp 1679581782
transform 1 0 109248 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_399
timestamp 1679581782
transform 1 0 109920 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_406
timestamp 1679581782
transform 1 0 110592 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_413
timestamp 1679581782
transform 1 0 111264 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_420
timestamp 1679581782
transform 1 0 111936 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_427
timestamp 1679581782
transform 1 0 112608 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_434
timestamp 1679581782
transform 1 0 113280 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_441
timestamp 1679581782
transform 1 0 113952 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_448
timestamp 1679581782
transform 1 0 114624 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_455
timestamp 1679581782
transform 1 0 115296 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_462
timestamp 1679581782
transform 1 0 115968 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_469
timestamp 1679581782
transform 1 0 116640 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_476
timestamp 1679581782
transform 1 0 117312 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_483
timestamp 1679581782
transform 1 0 117984 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_490
timestamp 1679581782
transform 1 0 118656 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_497
timestamp 1679581782
transform 1 0 119328 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_504
timestamp 1679581782
transform 1 0 120000 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_511
timestamp 1679581782
transform 1 0 120672 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_518
timestamp 1679581782
transform 1 0 121344 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_525
timestamp 1679581782
transform 1 0 122016 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_532
timestamp 1679581782
transform 1 0 122688 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_539
timestamp 1679581782
transform 1 0 123360 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_546
timestamp 1679581782
transform 1 0 124032 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_553
timestamp 1679581782
transform 1 0 124704 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_560
timestamp 1679581782
transform 1 0 125376 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_567
timestamp 1679581782
transform 1 0 126048 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_574
timestamp 1679581782
transform 1 0 126720 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_581
timestamp 1679581782
transform 1 0 127392 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_588
timestamp 1679581782
transform 1 0 128064 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_595
timestamp 1679581782
transform 1 0 128736 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_602
timestamp 1679581782
transform 1 0 129408 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_609
timestamp 1679581782
transform 1 0 130080 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_616
timestamp 1679581782
transform 1 0 130752 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_623
timestamp 1679581782
transform 1 0 131424 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_630
timestamp 1679581782
transform 1 0 132096 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_637
timestamp 1679581782
transform 1 0 132768 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_644
timestamp 1679581782
transform 1 0 133440 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_651
timestamp 1679581782
transform 1 0 134112 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_658
timestamp 1679581782
transform 1 0 134784 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_665
timestamp 1679581782
transform 1 0 135456 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_672
timestamp 1679581782
transform 1 0 136128 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_679
timestamp 1679581782
transform 1 0 136800 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_686
timestamp 1679581782
transform 1 0 137472 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_693
timestamp 1679581782
transform 1 0 138144 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_700
timestamp 1679581782
transform 1 0 138816 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_707
timestamp 1679581782
transform 1 0 139488 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_714
timestamp 1679581782
transform 1 0 140160 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_721
timestamp 1679581782
transform 1 0 140832 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_728
timestamp 1679581782
transform 1 0 141504 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_735
timestamp 1679581782
transform 1 0 142176 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_742
timestamp 1679581782
transform 1 0 142848 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_749
timestamp 1679581782
transform 1 0 143520 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_756
timestamp 1679581782
transform 1 0 144192 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_763
timestamp 1679581782
transform 1 0 144864 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_770
timestamp 1679581782
transform 1 0 145536 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_777
timestamp 1679581782
transform 1 0 146208 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_784
timestamp 1679581782
transform 1 0 146880 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_791
timestamp 1679581782
transform 1 0 147552 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_798
timestamp 1679581782
transform 1 0 148224 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_805
timestamp 1679581782
transform 1 0 148896 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_812
timestamp 1679581782
transform 1 0 149568 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_819
timestamp 1679581782
transform 1 0 150240 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_826
timestamp 1679581782
transform 1 0 150912 0 1 117180
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_833
timestamp 1679581782
transform 1 0 151584 0 1 117180
box -48 -56 720 834
use sg13g2_fill_1  FILLER_60_840
timestamp 1677579658
transform 1 0 152256 0 1 117180
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_0
timestamp 1679581782
transform 1 0 71616 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_7
timestamp 1679581782
transform 1 0 72288 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_14
timestamp 1679581782
transform 1 0 72960 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_21
timestamp 1679581782
transform 1 0 73632 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_28
timestamp 1679581782
transform 1 0 74304 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_35
timestamp 1679581782
transform 1 0 74976 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_42
timestamp 1679581782
transform 1 0 75648 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_49
timestamp 1679581782
transform 1 0 76320 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_56
timestamp 1679581782
transform 1 0 76992 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_63
timestamp 1679581782
transform 1 0 77664 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_70
timestamp 1679581782
transform 1 0 78336 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_77
timestamp 1679581782
transform 1 0 79008 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_84
timestamp 1679581782
transform 1 0 79680 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_91
timestamp 1679581782
transform 1 0 80352 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_98
timestamp 1679581782
transform 1 0 81024 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_105
timestamp 1679581782
transform 1 0 81696 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_112
timestamp 1679581782
transform 1 0 82368 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_119
timestamp 1679581782
transform 1 0 83040 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_126
timestamp 1679581782
transform 1 0 83712 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_133
timestamp 1679581782
transform 1 0 84384 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_140
timestamp 1679581782
transform 1 0 85056 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_147
timestamp 1679581782
transform 1 0 85728 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_154
timestamp 1679581782
transform 1 0 86400 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_161
timestamp 1679581782
transform 1 0 87072 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_168
timestamp 1679581782
transform 1 0 87744 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_175
timestamp 1679581782
transform 1 0 88416 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_182
timestamp 1679581782
transform 1 0 89088 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_189
timestamp 1679581782
transform 1 0 89760 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_196
timestamp 1679581782
transform 1 0 90432 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_203
timestamp 1679581782
transform 1 0 91104 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_210
timestamp 1679581782
transform 1 0 91776 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_217
timestamp 1679581782
transform 1 0 92448 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_224
timestamp 1679581782
transform 1 0 93120 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_231
timestamp 1679581782
transform 1 0 93792 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_238
timestamp 1679581782
transform 1 0 94464 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_245
timestamp 1679581782
transform 1 0 95136 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_252
timestamp 1679581782
transform 1 0 95808 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_259
timestamp 1679581782
transform 1 0 96480 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_266
timestamp 1679581782
transform 1 0 97152 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_273
timestamp 1679581782
transform 1 0 97824 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_280
timestamp 1679581782
transform 1 0 98496 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_287
timestamp 1679581782
transform 1 0 99168 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_294
timestamp 1679581782
transform 1 0 99840 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_301
timestamp 1679581782
transform 1 0 100512 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_308
timestamp 1679581782
transform 1 0 101184 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_315
timestamp 1679581782
transform 1 0 101856 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_322
timestamp 1679581782
transform 1 0 102528 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_329
timestamp 1679581782
transform 1 0 103200 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_336
timestamp 1679581782
transform 1 0 103872 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_343
timestamp 1679581782
transform 1 0 104544 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_350
timestamp 1679581782
transform 1 0 105216 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_357
timestamp 1679581782
transform 1 0 105888 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_364
timestamp 1679581782
transform 1 0 106560 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_371
timestamp 1679581782
transform 1 0 107232 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_378
timestamp 1679581782
transform 1 0 107904 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_385
timestamp 1679581782
transform 1 0 108576 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_392
timestamp 1679581782
transform 1 0 109248 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_399
timestamp 1679581782
transform 1 0 109920 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_406
timestamp 1679581782
transform 1 0 110592 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_413
timestamp 1679581782
transform 1 0 111264 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_420
timestamp 1679581782
transform 1 0 111936 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_427
timestamp 1679581782
transform 1 0 112608 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_434
timestamp 1679581782
transform 1 0 113280 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_441
timestamp 1679581782
transform 1 0 113952 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_448
timestamp 1679581782
transform 1 0 114624 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_455
timestamp 1679581782
transform 1 0 115296 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_462
timestamp 1679581782
transform 1 0 115968 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_469
timestamp 1679581782
transform 1 0 116640 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_476
timestamp 1679581782
transform 1 0 117312 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_483
timestamp 1679581782
transform 1 0 117984 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_490
timestamp 1679581782
transform 1 0 118656 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_497
timestamp 1679581782
transform 1 0 119328 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_504
timestamp 1679581782
transform 1 0 120000 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_511
timestamp 1679581782
transform 1 0 120672 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_518
timestamp 1679581782
transform 1 0 121344 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_525
timestamp 1679581782
transform 1 0 122016 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_532
timestamp 1679581782
transform 1 0 122688 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_539
timestamp 1679581782
transform 1 0 123360 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_546
timestamp 1679581782
transform 1 0 124032 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_553
timestamp 1679581782
transform 1 0 124704 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_560
timestamp 1679581782
transform 1 0 125376 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_567
timestamp 1679581782
transform 1 0 126048 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_574
timestamp 1679581782
transform 1 0 126720 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_581
timestamp 1679581782
transform 1 0 127392 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_588
timestamp 1679581782
transform 1 0 128064 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_595
timestamp 1679581782
transform 1 0 128736 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_602
timestamp 1679581782
transform 1 0 129408 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_609
timestamp 1679581782
transform 1 0 130080 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_616
timestamp 1679581782
transform 1 0 130752 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_623
timestamp 1679581782
transform 1 0 131424 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_630
timestamp 1679581782
transform 1 0 132096 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_637
timestamp 1679581782
transform 1 0 132768 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_644
timestamp 1679581782
transform 1 0 133440 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_651
timestamp 1679581782
transform 1 0 134112 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_658
timestamp 1679581782
transform 1 0 134784 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_665
timestamp 1679581782
transform 1 0 135456 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_672
timestamp 1679581782
transform 1 0 136128 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_679
timestamp 1679581782
transform 1 0 136800 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_686
timestamp 1679581782
transform 1 0 137472 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_693
timestamp 1679581782
transform 1 0 138144 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_700
timestamp 1679581782
transform 1 0 138816 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_707
timestamp 1679581782
transform 1 0 139488 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_714
timestamp 1679581782
transform 1 0 140160 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_721
timestamp 1679581782
transform 1 0 140832 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_728
timestamp 1679581782
transform 1 0 141504 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_735
timestamp 1679581782
transform 1 0 142176 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_742
timestamp 1679581782
transform 1 0 142848 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_749
timestamp 1679581782
transform 1 0 143520 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_756
timestamp 1679581782
transform 1 0 144192 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_763
timestamp 1679581782
transform 1 0 144864 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_770
timestamp 1679581782
transform 1 0 145536 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_777
timestamp 1679581782
transform 1 0 146208 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_784
timestamp 1679581782
transform 1 0 146880 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_791
timestamp 1679581782
transform 1 0 147552 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_798
timestamp 1679581782
transform 1 0 148224 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_805
timestamp 1679581782
transform 1 0 148896 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_812
timestamp 1679581782
transform 1 0 149568 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_819
timestamp 1679581782
transform 1 0 150240 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_826
timestamp 1679581782
transform 1 0 150912 0 -1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_833
timestamp 1679581782
transform 1 0 151584 0 -1 118692
box -48 -56 720 834
use sg13g2_fill_1  FILLER_61_840
timestamp 1677579658
transform 1 0 152256 0 -1 118692
box -48 -56 144 834
use sg13g2_decap_8  FILLER_62_0
timestamp 1679581782
transform 1 0 71616 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_7
timestamp 1679581782
transform 1 0 72288 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_14
timestamp 1679581782
transform 1 0 72960 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_21
timestamp 1679581782
transform 1 0 73632 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_28
timestamp 1679581782
transform 1 0 74304 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_35
timestamp 1679581782
transform 1 0 74976 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_42
timestamp 1679581782
transform 1 0 75648 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_49
timestamp 1679581782
transform 1 0 76320 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_56
timestamp 1679581782
transform 1 0 76992 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_63
timestamp 1679581782
transform 1 0 77664 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_70
timestamp 1679581782
transform 1 0 78336 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_77
timestamp 1679581782
transform 1 0 79008 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_84
timestamp 1679581782
transform 1 0 79680 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_91
timestamp 1679581782
transform 1 0 80352 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_98
timestamp 1679581782
transform 1 0 81024 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_105
timestamp 1679581782
transform 1 0 81696 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_112
timestamp 1679581782
transform 1 0 82368 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_119
timestamp 1679581782
transform 1 0 83040 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_126
timestamp 1679581782
transform 1 0 83712 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_133
timestamp 1679581782
transform 1 0 84384 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_140
timestamp 1679581782
transform 1 0 85056 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_147
timestamp 1679581782
transform 1 0 85728 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_154
timestamp 1679581782
transform 1 0 86400 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_161
timestamp 1679581782
transform 1 0 87072 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_168
timestamp 1679581782
transform 1 0 87744 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_175
timestamp 1679581782
transform 1 0 88416 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_182
timestamp 1679581782
transform 1 0 89088 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_189
timestamp 1679581782
transform 1 0 89760 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_196
timestamp 1679581782
transform 1 0 90432 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_203
timestamp 1679581782
transform 1 0 91104 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_210
timestamp 1679581782
transform 1 0 91776 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_217
timestamp 1679581782
transform 1 0 92448 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_224
timestamp 1679581782
transform 1 0 93120 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_231
timestamp 1679581782
transform 1 0 93792 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_238
timestamp 1679581782
transform 1 0 94464 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_245
timestamp 1679581782
transform 1 0 95136 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_252
timestamp 1679581782
transform 1 0 95808 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_259
timestamp 1679581782
transform 1 0 96480 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_266
timestamp 1679581782
transform 1 0 97152 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_273
timestamp 1679581782
transform 1 0 97824 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_280
timestamp 1679581782
transform 1 0 98496 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_287
timestamp 1679581782
transform 1 0 99168 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_294
timestamp 1679581782
transform 1 0 99840 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_301
timestamp 1679581782
transform 1 0 100512 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_308
timestamp 1679581782
transform 1 0 101184 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_315
timestamp 1679581782
transform 1 0 101856 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_322
timestamp 1679581782
transform 1 0 102528 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_329
timestamp 1679581782
transform 1 0 103200 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_336
timestamp 1679581782
transform 1 0 103872 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_343
timestamp 1679581782
transform 1 0 104544 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_350
timestamp 1679581782
transform 1 0 105216 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_357
timestamp 1679581782
transform 1 0 105888 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_364
timestamp 1679581782
transform 1 0 106560 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_371
timestamp 1679581782
transform 1 0 107232 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_378
timestamp 1679581782
transform 1 0 107904 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_385
timestamp 1679581782
transform 1 0 108576 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_392
timestamp 1679581782
transform 1 0 109248 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_399
timestamp 1679581782
transform 1 0 109920 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_406
timestamp 1679581782
transform 1 0 110592 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_413
timestamp 1679581782
transform 1 0 111264 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_420
timestamp 1679581782
transform 1 0 111936 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_427
timestamp 1679581782
transform 1 0 112608 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_434
timestamp 1679581782
transform 1 0 113280 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_441
timestamp 1679581782
transform 1 0 113952 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_448
timestamp 1679581782
transform 1 0 114624 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_455
timestamp 1679581782
transform 1 0 115296 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_462
timestamp 1679581782
transform 1 0 115968 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_469
timestamp 1679581782
transform 1 0 116640 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_476
timestamp 1679581782
transform 1 0 117312 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_483
timestamp 1679581782
transform 1 0 117984 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_490
timestamp 1679581782
transform 1 0 118656 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_497
timestamp 1679581782
transform 1 0 119328 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_504
timestamp 1679581782
transform 1 0 120000 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_511
timestamp 1679581782
transform 1 0 120672 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_518
timestamp 1679581782
transform 1 0 121344 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_525
timestamp 1679581782
transform 1 0 122016 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_532
timestamp 1679581782
transform 1 0 122688 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_539
timestamp 1679581782
transform 1 0 123360 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_546
timestamp 1679581782
transform 1 0 124032 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_553
timestamp 1679581782
transform 1 0 124704 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_560
timestamp 1679581782
transform 1 0 125376 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_567
timestamp 1679581782
transform 1 0 126048 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_574
timestamp 1679581782
transform 1 0 126720 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_581
timestamp 1679581782
transform 1 0 127392 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_588
timestamp 1679581782
transform 1 0 128064 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_595
timestamp 1679581782
transform 1 0 128736 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_602
timestamp 1679581782
transform 1 0 129408 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_609
timestamp 1679581782
transform 1 0 130080 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_616
timestamp 1679581782
transform 1 0 130752 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_623
timestamp 1679581782
transform 1 0 131424 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_630
timestamp 1679581782
transform 1 0 132096 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_637
timestamp 1679581782
transform 1 0 132768 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_644
timestamp 1679581782
transform 1 0 133440 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_651
timestamp 1679581782
transform 1 0 134112 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_658
timestamp 1679581782
transform 1 0 134784 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_665
timestamp 1679581782
transform 1 0 135456 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_672
timestamp 1679581782
transform 1 0 136128 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_679
timestamp 1679581782
transform 1 0 136800 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_686
timestamp 1679581782
transform 1 0 137472 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_693
timestamp 1679581782
transform 1 0 138144 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_700
timestamp 1679581782
transform 1 0 138816 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_707
timestamp 1679581782
transform 1 0 139488 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_714
timestamp 1679581782
transform 1 0 140160 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_721
timestamp 1679581782
transform 1 0 140832 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_728
timestamp 1679581782
transform 1 0 141504 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_735
timestamp 1679581782
transform 1 0 142176 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_742
timestamp 1679581782
transform 1 0 142848 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_749
timestamp 1679581782
transform 1 0 143520 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_756
timestamp 1679581782
transform 1 0 144192 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_763
timestamp 1679581782
transform 1 0 144864 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_770
timestamp 1679581782
transform 1 0 145536 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_777
timestamp 1679581782
transform 1 0 146208 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_784
timestamp 1679581782
transform 1 0 146880 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_791
timestamp 1679581782
transform 1 0 147552 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_798
timestamp 1679581782
transform 1 0 148224 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_805
timestamp 1679581782
transform 1 0 148896 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_812
timestamp 1679581782
transform 1 0 149568 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_819
timestamp 1679581782
transform 1 0 150240 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_826
timestamp 1679581782
transform 1 0 150912 0 1 118692
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_833
timestamp 1679581782
transform 1 0 151584 0 1 118692
box -48 -56 720 834
use sg13g2_fill_1  FILLER_62_840
timestamp 1677579658
transform 1 0 152256 0 1 118692
box -48 -56 144 834
use sg13g2_decap_8  FILLER_63_0
timestamp 1679581782
transform 1 0 71616 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_7
timestamp 1679581782
transform 1 0 72288 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_14
timestamp 1679581782
transform 1 0 72960 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_21
timestamp 1679581782
transform 1 0 73632 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_28
timestamp 1679581782
transform 1 0 74304 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_35
timestamp 1679581782
transform 1 0 74976 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_42
timestamp 1679581782
transform 1 0 75648 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_49
timestamp 1679581782
transform 1 0 76320 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_56
timestamp 1679581782
transform 1 0 76992 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_63
timestamp 1679581782
transform 1 0 77664 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_70
timestamp 1679581782
transform 1 0 78336 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_77
timestamp 1679581782
transform 1 0 79008 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_84
timestamp 1679581782
transform 1 0 79680 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_91
timestamp 1679581782
transform 1 0 80352 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_98
timestamp 1679581782
transform 1 0 81024 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_105
timestamp 1679581782
transform 1 0 81696 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_112
timestamp 1679581782
transform 1 0 82368 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_119
timestamp 1679581782
transform 1 0 83040 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_126
timestamp 1679581782
transform 1 0 83712 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_133
timestamp 1679581782
transform 1 0 84384 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_140
timestamp 1679581782
transform 1 0 85056 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_147
timestamp 1679581782
transform 1 0 85728 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_154
timestamp 1679581782
transform 1 0 86400 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_161
timestamp 1679581782
transform 1 0 87072 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_168
timestamp 1679581782
transform 1 0 87744 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_175
timestamp 1679581782
transform 1 0 88416 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_182
timestamp 1679581782
transform 1 0 89088 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_189
timestamp 1679581782
transform 1 0 89760 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_196
timestamp 1679581782
transform 1 0 90432 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_203
timestamp 1679581782
transform 1 0 91104 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_210
timestamp 1679581782
transform 1 0 91776 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_217
timestamp 1679581782
transform 1 0 92448 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_224
timestamp 1679581782
transform 1 0 93120 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_231
timestamp 1679581782
transform 1 0 93792 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_238
timestamp 1679581782
transform 1 0 94464 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_245
timestamp 1679581782
transform 1 0 95136 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_252
timestamp 1679581782
transform 1 0 95808 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_259
timestamp 1679581782
transform 1 0 96480 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_266
timestamp 1679581782
transform 1 0 97152 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_273
timestamp 1679581782
transform 1 0 97824 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_280
timestamp 1679581782
transform 1 0 98496 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_287
timestamp 1679581782
transform 1 0 99168 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_294
timestamp 1679581782
transform 1 0 99840 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_301
timestamp 1679581782
transform 1 0 100512 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_308
timestamp 1679581782
transform 1 0 101184 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_315
timestamp 1679581782
transform 1 0 101856 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_322
timestamp 1679581782
transform 1 0 102528 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_329
timestamp 1679581782
transform 1 0 103200 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_336
timestamp 1679581782
transform 1 0 103872 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_343
timestamp 1679581782
transform 1 0 104544 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_350
timestamp 1679581782
transform 1 0 105216 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_357
timestamp 1679581782
transform 1 0 105888 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_364
timestamp 1679581782
transform 1 0 106560 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_371
timestamp 1679581782
transform 1 0 107232 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_378
timestamp 1679581782
transform 1 0 107904 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_385
timestamp 1679581782
transform 1 0 108576 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_392
timestamp 1679581782
transform 1 0 109248 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_399
timestamp 1679581782
transform 1 0 109920 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_406
timestamp 1679581782
transform 1 0 110592 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_413
timestamp 1679581782
transform 1 0 111264 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_420
timestamp 1679581782
transform 1 0 111936 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_427
timestamp 1679581782
transform 1 0 112608 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_434
timestamp 1679581782
transform 1 0 113280 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_441
timestamp 1679581782
transform 1 0 113952 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_448
timestamp 1679581782
transform 1 0 114624 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_455
timestamp 1679581782
transform 1 0 115296 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_462
timestamp 1679581782
transform 1 0 115968 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_469
timestamp 1679581782
transform 1 0 116640 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_476
timestamp 1679581782
transform 1 0 117312 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_483
timestamp 1679581782
transform 1 0 117984 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_490
timestamp 1679581782
transform 1 0 118656 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_497
timestamp 1679581782
transform 1 0 119328 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_504
timestamp 1679581782
transform 1 0 120000 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_511
timestamp 1679581782
transform 1 0 120672 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_518
timestamp 1679581782
transform 1 0 121344 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_525
timestamp 1679581782
transform 1 0 122016 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_532
timestamp 1679581782
transform 1 0 122688 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_539
timestamp 1679581782
transform 1 0 123360 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_546
timestamp 1679581782
transform 1 0 124032 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_553
timestamp 1679581782
transform 1 0 124704 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_560
timestamp 1679581782
transform 1 0 125376 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_567
timestamp 1679581782
transform 1 0 126048 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_574
timestamp 1679581782
transform 1 0 126720 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_581
timestamp 1679581782
transform 1 0 127392 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_588
timestamp 1679581782
transform 1 0 128064 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_595
timestamp 1679581782
transform 1 0 128736 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_602
timestamp 1679581782
transform 1 0 129408 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_609
timestamp 1679581782
transform 1 0 130080 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_616
timestamp 1679581782
transform 1 0 130752 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_623
timestamp 1679581782
transform 1 0 131424 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_630
timestamp 1679581782
transform 1 0 132096 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_637
timestamp 1679581782
transform 1 0 132768 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_644
timestamp 1679581782
transform 1 0 133440 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_651
timestamp 1679581782
transform 1 0 134112 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_658
timestamp 1679581782
transform 1 0 134784 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_665
timestamp 1679581782
transform 1 0 135456 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_672
timestamp 1679581782
transform 1 0 136128 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_679
timestamp 1679581782
transform 1 0 136800 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_686
timestamp 1679581782
transform 1 0 137472 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_693
timestamp 1679581782
transform 1 0 138144 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_700
timestamp 1679581782
transform 1 0 138816 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_707
timestamp 1679581782
transform 1 0 139488 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_714
timestamp 1679581782
transform 1 0 140160 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_721
timestamp 1679581782
transform 1 0 140832 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_728
timestamp 1679581782
transform 1 0 141504 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_735
timestamp 1679581782
transform 1 0 142176 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_742
timestamp 1679581782
transform 1 0 142848 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_749
timestamp 1679581782
transform 1 0 143520 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_756
timestamp 1679581782
transform 1 0 144192 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_763
timestamp 1679581782
transform 1 0 144864 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_770
timestamp 1679581782
transform 1 0 145536 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_777
timestamp 1679581782
transform 1 0 146208 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_784
timestamp 1679581782
transform 1 0 146880 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_791
timestamp 1679581782
transform 1 0 147552 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_798
timestamp 1679581782
transform 1 0 148224 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_805
timestamp 1679581782
transform 1 0 148896 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_812
timestamp 1679581782
transform 1 0 149568 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_819
timestamp 1679581782
transform 1 0 150240 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_826
timestamp 1679581782
transform 1 0 150912 0 -1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_833
timestamp 1679581782
transform 1 0 151584 0 -1 120204
box -48 -56 720 834
use sg13g2_fill_1  FILLER_63_840
timestamp 1677579658
transform 1 0 152256 0 -1 120204
box -48 -56 144 834
use sg13g2_decap_8  FILLER_64_0
timestamp 1679581782
transform 1 0 71616 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_7
timestamp 1679581782
transform 1 0 72288 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_14
timestamp 1679581782
transform 1 0 72960 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_21
timestamp 1679581782
transform 1 0 73632 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_28
timestamp 1679581782
transform 1 0 74304 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_35
timestamp 1679581782
transform 1 0 74976 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_42
timestamp 1679581782
transform 1 0 75648 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_49
timestamp 1679581782
transform 1 0 76320 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_56
timestamp 1679581782
transform 1 0 76992 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_63
timestamp 1679581782
transform 1 0 77664 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_70
timestamp 1679581782
transform 1 0 78336 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_77
timestamp 1679581782
transform 1 0 79008 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_84
timestamp 1679581782
transform 1 0 79680 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_91
timestamp 1679581782
transform 1 0 80352 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_98
timestamp 1679581782
transform 1 0 81024 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_105
timestamp 1679581782
transform 1 0 81696 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_112
timestamp 1679581782
transform 1 0 82368 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_119
timestamp 1679581782
transform 1 0 83040 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_126
timestamp 1679581782
transform 1 0 83712 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_133
timestamp 1679581782
transform 1 0 84384 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_140
timestamp 1679581782
transform 1 0 85056 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_147
timestamp 1679581782
transform 1 0 85728 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_154
timestamp 1679581782
transform 1 0 86400 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_161
timestamp 1679581782
transform 1 0 87072 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_168
timestamp 1679581782
transform 1 0 87744 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_175
timestamp 1679581782
transform 1 0 88416 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_182
timestamp 1679581782
transform 1 0 89088 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_189
timestamp 1679581782
transform 1 0 89760 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_196
timestamp 1679581782
transform 1 0 90432 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_203
timestamp 1679581782
transform 1 0 91104 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_210
timestamp 1679581782
transform 1 0 91776 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_217
timestamp 1679581782
transform 1 0 92448 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_224
timestamp 1679581782
transform 1 0 93120 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_231
timestamp 1679581782
transform 1 0 93792 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_238
timestamp 1679581782
transform 1 0 94464 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_245
timestamp 1679581782
transform 1 0 95136 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_252
timestamp 1679581782
transform 1 0 95808 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_259
timestamp 1679581782
transform 1 0 96480 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_266
timestamp 1679581782
transform 1 0 97152 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_273
timestamp 1679581782
transform 1 0 97824 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_280
timestamp 1679581782
transform 1 0 98496 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_287
timestamp 1679581782
transform 1 0 99168 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_294
timestamp 1679581782
transform 1 0 99840 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_301
timestamp 1679581782
transform 1 0 100512 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_308
timestamp 1679581782
transform 1 0 101184 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_315
timestamp 1679581782
transform 1 0 101856 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_322
timestamp 1679581782
transform 1 0 102528 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_329
timestamp 1679581782
transform 1 0 103200 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_336
timestamp 1679581782
transform 1 0 103872 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_343
timestamp 1679581782
transform 1 0 104544 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_350
timestamp 1679581782
transform 1 0 105216 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_357
timestamp 1679581782
transform 1 0 105888 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_364
timestamp 1679581782
transform 1 0 106560 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_371
timestamp 1679581782
transform 1 0 107232 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_378
timestamp 1679581782
transform 1 0 107904 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_385
timestamp 1679581782
transform 1 0 108576 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_392
timestamp 1679581782
transform 1 0 109248 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_399
timestamp 1679581782
transform 1 0 109920 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_406
timestamp 1679581782
transform 1 0 110592 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_413
timestamp 1679581782
transform 1 0 111264 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_420
timestamp 1679581782
transform 1 0 111936 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_427
timestamp 1679581782
transform 1 0 112608 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_434
timestamp 1679581782
transform 1 0 113280 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_441
timestamp 1679581782
transform 1 0 113952 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_448
timestamp 1679581782
transform 1 0 114624 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_455
timestamp 1679581782
transform 1 0 115296 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_462
timestamp 1679581782
transform 1 0 115968 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_469
timestamp 1679581782
transform 1 0 116640 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_476
timestamp 1679581782
transform 1 0 117312 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_483
timestamp 1679581782
transform 1 0 117984 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_490
timestamp 1679581782
transform 1 0 118656 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_497
timestamp 1679581782
transform 1 0 119328 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_504
timestamp 1679581782
transform 1 0 120000 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_511
timestamp 1679581782
transform 1 0 120672 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_518
timestamp 1679581782
transform 1 0 121344 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_525
timestamp 1679581782
transform 1 0 122016 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_532
timestamp 1679581782
transform 1 0 122688 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_539
timestamp 1679581782
transform 1 0 123360 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_546
timestamp 1679581782
transform 1 0 124032 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_553
timestamp 1679581782
transform 1 0 124704 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_560
timestamp 1679581782
transform 1 0 125376 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_567
timestamp 1679581782
transform 1 0 126048 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_574
timestamp 1679581782
transform 1 0 126720 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_581
timestamp 1679581782
transform 1 0 127392 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_588
timestamp 1679581782
transform 1 0 128064 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_595
timestamp 1679581782
transform 1 0 128736 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_602
timestamp 1679581782
transform 1 0 129408 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_609
timestamp 1679581782
transform 1 0 130080 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_616
timestamp 1679581782
transform 1 0 130752 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_623
timestamp 1679581782
transform 1 0 131424 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_630
timestamp 1679581782
transform 1 0 132096 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_637
timestamp 1679581782
transform 1 0 132768 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_644
timestamp 1679581782
transform 1 0 133440 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_651
timestamp 1679581782
transform 1 0 134112 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_658
timestamp 1679581782
transform 1 0 134784 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_665
timestamp 1679581782
transform 1 0 135456 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_672
timestamp 1679581782
transform 1 0 136128 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_679
timestamp 1679581782
transform 1 0 136800 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_686
timestamp 1679581782
transform 1 0 137472 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_693
timestamp 1679581782
transform 1 0 138144 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_700
timestamp 1679581782
transform 1 0 138816 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_707
timestamp 1679581782
transform 1 0 139488 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_714
timestamp 1679581782
transform 1 0 140160 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_721
timestamp 1679581782
transform 1 0 140832 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_728
timestamp 1679581782
transform 1 0 141504 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_735
timestamp 1679581782
transform 1 0 142176 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_742
timestamp 1679581782
transform 1 0 142848 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_749
timestamp 1679581782
transform 1 0 143520 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_756
timestamp 1679581782
transform 1 0 144192 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_763
timestamp 1679581782
transform 1 0 144864 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_770
timestamp 1679581782
transform 1 0 145536 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_777
timestamp 1679581782
transform 1 0 146208 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_784
timestamp 1679581782
transform 1 0 146880 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_791
timestamp 1679581782
transform 1 0 147552 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_798
timestamp 1679581782
transform 1 0 148224 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_805
timestamp 1679581782
transform 1 0 148896 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_812
timestamp 1679581782
transform 1 0 149568 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_819
timestamp 1679581782
transform 1 0 150240 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_826
timestamp 1679581782
transform 1 0 150912 0 1 120204
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_833
timestamp 1679581782
transform 1 0 151584 0 1 120204
box -48 -56 720 834
use sg13g2_fill_1  FILLER_64_840
timestamp 1677579658
transform 1 0 152256 0 1 120204
box -48 -56 144 834
use sg13g2_decap_8  FILLER_65_0
timestamp 1679581782
transform 1 0 71616 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_7
timestamp 1679581782
transform 1 0 72288 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_14
timestamp 1679581782
transform 1 0 72960 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_21
timestamp 1679581782
transform 1 0 73632 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_28
timestamp 1679581782
transform 1 0 74304 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_35
timestamp 1679581782
transform 1 0 74976 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_42
timestamp 1679581782
transform 1 0 75648 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_49
timestamp 1679581782
transform 1 0 76320 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_56
timestamp 1679581782
transform 1 0 76992 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_63
timestamp 1679581782
transform 1 0 77664 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_70
timestamp 1679581782
transform 1 0 78336 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_77
timestamp 1679581782
transform 1 0 79008 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_84
timestamp 1679581782
transform 1 0 79680 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_91
timestamp 1679581782
transform 1 0 80352 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_98
timestamp 1679581782
transform 1 0 81024 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_105
timestamp 1679581782
transform 1 0 81696 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_112
timestamp 1679581782
transform 1 0 82368 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_119
timestamp 1679581782
transform 1 0 83040 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_126
timestamp 1679581782
transform 1 0 83712 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_133
timestamp 1679581782
transform 1 0 84384 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_140
timestamp 1679581782
transform 1 0 85056 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_147
timestamp 1679581782
transform 1 0 85728 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_154
timestamp 1679581782
transform 1 0 86400 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_161
timestamp 1679581782
transform 1 0 87072 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_168
timestamp 1679581782
transform 1 0 87744 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_175
timestamp 1679581782
transform 1 0 88416 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_182
timestamp 1679581782
transform 1 0 89088 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_189
timestamp 1679581782
transform 1 0 89760 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_196
timestamp 1679581782
transform 1 0 90432 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_203
timestamp 1679581782
transform 1 0 91104 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_210
timestamp 1679581782
transform 1 0 91776 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_217
timestamp 1679581782
transform 1 0 92448 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_224
timestamp 1679581782
transform 1 0 93120 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_231
timestamp 1679581782
transform 1 0 93792 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_238
timestamp 1679581782
transform 1 0 94464 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_245
timestamp 1679581782
transform 1 0 95136 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_252
timestamp 1679581782
transform 1 0 95808 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_259
timestamp 1679581782
transform 1 0 96480 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_266
timestamp 1679581782
transform 1 0 97152 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_273
timestamp 1679581782
transform 1 0 97824 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_280
timestamp 1679581782
transform 1 0 98496 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_287
timestamp 1679581782
transform 1 0 99168 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_294
timestamp 1679581782
transform 1 0 99840 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_301
timestamp 1679581782
transform 1 0 100512 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_308
timestamp 1679581782
transform 1 0 101184 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_315
timestamp 1679581782
transform 1 0 101856 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_322
timestamp 1679581782
transform 1 0 102528 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_329
timestamp 1679581782
transform 1 0 103200 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_336
timestamp 1679581782
transform 1 0 103872 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_343
timestamp 1679581782
transform 1 0 104544 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_350
timestamp 1679581782
transform 1 0 105216 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_357
timestamp 1679581782
transform 1 0 105888 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_364
timestamp 1679581782
transform 1 0 106560 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_371
timestamp 1679581782
transform 1 0 107232 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_378
timestamp 1679581782
transform 1 0 107904 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_385
timestamp 1679581782
transform 1 0 108576 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_392
timestamp 1679581782
transform 1 0 109248 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_399
timestamp 1679581782
transform 1 0 109920 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_406
timestamp 1679581782
transform 1 0 110592 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_413
timestamp 1679581782
transform 1 0 111264 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_420
timestamp 1679581782
transform 1 0 111936 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_427
timestamp 1679581782
transform 1 0 112608 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_434
timestamp 1679581782
transform 1 0 113280 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_441
timestamp 1679581782
transform 1 0 113952 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_448
timestamp 1679581782
transform 1 0 114624 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_455
timestamp 1679581782
transform 1 0 115296 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_462
timestamp 1679581782
transform 1 0 115968 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_469
timestamp 1679581782
transform 1 0 116640 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_476
timestamp 1679581782
transform 1 0 117312 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_483
timestamp 1679581782
transform 1 0 117984 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_490
timestamp 1679581782
transform 1 0 118656 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_497
timestamp 1679581782
transform 1 0 119328 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_504
timestamp 1679581782
transform 1 0 120000 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_511
timestamp 1679581782
transform 1 0 120672 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_518
timestamp 1679581782
transform 1 0 121344 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_525
timestamp 1679581782
transform 1 0 122016 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_532
timestamp 1679581782
transform 1 0 122688 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_539
timestamp 1679581782
transform 1 0 123360 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_546
timestamp 1679581782
transform 1 0 124032 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_553
timestamp 1679581782
transform 1 0 124704 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_560
timestamp 1679581782
transform 1 0 125376 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_567
timestamp 1679581782
transform 1 0 126048 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_574
timestamp 1679581782
transform 1 0 126720 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_581
timestamp 1679581782
transform 1 0 127392 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_588
timestamp 1679581782
transform 1 0 128064 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_595
timestamp 1679581782
transform 1 0 128736 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_602
timestamp 1679581782
transform 1 0 129408 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_609
timestamp 1679581782
transform 1 0 130080 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_616
timestamp 1679581782
transform 1 0 130752 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_623
timestamp 1679581782
transform 1 0 131424 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_630
timestamp 1679581782
transform 1 0 132096 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_637
timestamp 1679581782
transform 1 0 132768 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_644
timestamp 1679581782
transform 1 0 133440 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_651
timestamp 1679581782
transform 1 0 134112 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_658
timestamp 1679581782
transform 1 0 134784 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_665
timestamp 1679581782
transform 1 0 135456 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_672
timestamp 1679581782
transform 1 0 136128 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_679
timestamp 1679581782
transform 1 0 136800 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_686
timestamp 1679581782
transform 1 0 137472 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_693
timestamp 1679581782
transform 1 0 138144 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_700
timestamp 1679581782
transform 1 0 138816 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_707
timestamp 1679581782
transform 1 0 139488 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_714
timestamp 1679581782
transform 1 0 140160 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_721
timestamp 1679581782
transform 1 0 140832 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_728
timestamp 1679581782
transform 1 0 141504 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_735
timestamp 1679581782
transform 1 0 142176 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_742
timestamp 1679581782
transform 1 0 142848 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_749
timestamp 1679581782
transform 1 0 143520 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_756
timestamp 1679581782
transform 1 0 144192 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_763
timestamp 1679581782
transform 1 0 144864 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_770
timestamp 1679581782
transform 1 0 145536 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_777
timestamp 1679581782
transform 1 0 146208 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_784
timestamp 1679581782
transform 1 0 146880 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_791
timestamp 1679581782
transform 1 0 147552 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_798
timestamp 1679581782
transform 1 0 148224 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_805
timestamp 1679581782
transform 1 0 148896 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_812
timestamp 1679581782
transform 1 0 149568 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_819
timestamp 1679581782
transform 1 0 150240 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_826
timestamp 1679581782
transform 1 0 150912 0 -1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_833
timestamp 1679581782
transform 1 0 151584 0 -1 121716
box -48 -56 720 834
use sg13g2_fill_1  FILLER_65_840
timestamp 1677579658
transform 1 0 152256 0 -1 121716
box -48 -56 144 834
use sg13g2_decap_8  FILLER_66_0
timestamp 1679581782
transform 1 0 71616 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_7
timestamp 1679581782
transform 1 0 72288 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_14
timestamp 1679581782
transform 1 0 72960 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_21
timestamp 1679581782
transform 1 0 73632 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_28
timestamp 1679581782
transform 1 0 74304 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_35
timestamp 1679581782
transform 1 0 74976 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_42
timestamp 1679581782
transform 1 0 75648 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_49
timestamp 1679581782
transform 1 0 76320 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_56
timestamp 1679581782
transform 1 0 76992 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_63
timestamp 1679581782
transform 1 0 77664 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_70
timestamp 1679581782
transform 1 0 78336 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_77
timestamp 1679581782
transform 1 0 79008 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_84
timestamp 1679581782
transform 1 0 79680 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_91
timestamp 1679581782
transform 1 0 80352 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_98
timestamp 1679581782
transform 1 0 81024 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_105
timestamp 1679581782
transform 1 0 81696 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_112
timestamp 1679581782
transform 1 0 82368 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_119
timestamp 1679581782
transform 1 0 83040 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_126
timestamp 1679581782
transform 1 0 83712 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_133
timestamp 1679581782
transform 1 0 84384 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_140
timestamp 1679581782
transform 1 0 85056 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_147
timestamp 1679581782
transform 1 0 85728 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_154
timestamp 1679581782
transform 1 0 86400 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_161
timestamp 1679581782
transform 1 0 87072 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_168
timestamp 1679581782
transform 1 0 87744 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_175
timestamp 1679581782
transform 1 0 88416 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_182
timestamp 1679581782
transform 1 0 89088 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_189
timestamp 1679581782
transform 1 0 89760 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_196
timestamp 1679581782
transform 1 0 90432 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_203
timestamp 1679581782
transform 1 0 91104 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_210
timestamp 1679581782
transform 1 0 91776 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_217
timestamp 1679581782
transform 1 0 92448 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_224
timestamp 1679581782
transform 1 0 93120 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_231
timestamp 1679581782
transform 1 0 93792 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_238
timestamp 1679581782
transform 1 0 94464 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_245
timestamp 1679581782
transform 1 0 95136 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_252
timestamp 1679581782
transform 1 0 95808 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_259
timestamp 1679581782
transform 1 0 96480 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_266
timestamp 1679581782
transform 1 0 97152 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_273
timestamp 1679581782
transform 1 0 97824 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_280
timestamp 1679581782
transform 1 0 98496 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_287
timestamp 1679581782
transform 1 0 99168 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_294
timestamp 1679581782
transform 1 0 99840 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_301
timestamp 1679581782
transform 1 0 100512 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_308
timestamp 1679581782
transform 1 0 101184 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_315
timestamp 1679581782
transform 1 0 101856 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_322
timestamp 1679581782
transform 1 0 102528 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_329
timestamp 1679581782
transform 1 0 103200 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_336
timestamp 1679581782
transform 1 0 103872 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_343
timestamp 1679581782
transform 1 0 104544 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_350
timestamp 1679581782
transform 1 0 105216 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_357
timestamp 1679581782
transform 1 0 105888 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_364
timestamp 1679581782
transform 1 0 106560 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_371
timestamp 1679581782
transform 1 0 107232 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_378
timestamp 1679581782
transform 1 0 107904 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_385
timestamp 1679581782
transform 1 0 108576 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_392
timestamp 1679581782
transform 1 0 109248 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_399
timestamp 1679581782
transform 1 0 109920 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_406
timestamp 1679581782
transform 1 0 110592 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_413
timestamp 1679581782
transform 1 0 111264 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_420
timestamp 1679581782
transform 1 0 111936 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_427
timestamp 1679581782
transform 1 0 112608 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_434
timestamp 1679581782
transform 1 0 113280 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_441
timestamp 1679581782
transform 1 0 113952 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_448
timestamp 1679581782
transform 1 0 114624 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_455
timestamp 1679581782
transform 1 0 115296 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_462
timestamp 1679581782
transform 1 0 115968 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_469
timestamp 1679581782
transform 1 0 116640 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_476
timestamp 1679581782
transform 1 0 117312 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_483
timestamp 1679581782
transform 1 0 117984 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_490
timestamp 1679581782
transform 1 0 118656 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_497
timestamp 1679581782
transform 1 0 119328 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_504
timestamp 1679581782
transform 1 0 120000 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_511
timestamp 1679581782
transform 1 0 120672 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_518
timestamp 1679581782
transform 1 0 121344 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_525
timestamp 1679581782
transform 1 0 122016 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_532
timestamp 1679581782
transform 1 0 122688 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_539
timestamp 1679581782
transform 1 0 123360 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_546
timestamp 1679581782
transform 1 0 124032 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_553
timestamp 1679581782
transform 1 0 124704 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_560
timestamp 1679581782
transform 1 0 125376 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_567
timestamp 1679581782
transform 1 0 126048 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_574
timestamp 1679581782
transform 1 0 126720 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_581
timestamp 1679581782
transform 1 0 127392 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_588
timestamp 1679581782
transform 1 0 128064 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_595
timestamp 1679581782
transform 1 0 128736 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_602
timestamp 1679581782
transform 1 0 129408 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_609
timestamp 1679581782
transform 1 0 130080 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_616
timestamp 1679581782
transform 1 0 130752 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_623
timestamp 1679581782
transform 1 0 131424 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_630
timestamp 1679581782
transform 1 0 132096 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_637
timestamp 1679581782
transform 1 0 132768 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_644
timestamp 1679581782
transform 1 0 133440 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_651
timestamp 1679581782
transform 1 0 134112 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_658
timestamp 1679581782
transform 1 0 134784 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_665
timestamp 1679581782
transform 1 0 135456 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_672
timestamp 1679581782
transform 1 0 136128 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_679
timestamp 1679581782
transform 1 0 136800 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_686
timestamp 1679581782
transform 1 0 137472 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_693
timestamp 1679581782
transform 1 0 138144 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_700
timestamp 1679581782
transform 1 0 138816 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_707
timestamp 1679581782
transform 1 0 139488 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_714
timestamp 1679581782
transform 1 0 140160 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_721
timestamp 1679581782
transform 1 0 140832 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_728
timestamp 1679581782
transform 1 0 141504 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_735
timestamp 1679581782
transform 1 0 142176 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_742
timestamp 1679581782
transform 1 0 142848 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_749
timestamp 1679581782
transform 1 0 143520 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_756
timestamp 1679581782
transform 1 0 144192 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_763
timestamp 1679581782
transform 1 0 144864 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_770
timestamp 1679581782
transform 1 0 145536 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_777
timestamp 1679581782
transform 1 0 146208 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_784
timestamp 1679581782
transform 1 0 146880 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_791
timestamp 1679581782
transform 1 0 147552 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_798
timestamp 1679581782
transform 1 0 148224 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_805
timestamp 1679581782
transform 1 0 148896 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_812
timestamp 1679581782
transform 1 0 149568 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_819
timestamp 1679581782
transform 1 0 150240 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_826
timestamp 1679581782
transform 1 0 150912 0 1 121716
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_833
timestamp 1679581782
transform 1 0 151584 0 1 121716
box -48 -56 720 834
use sg13g2_fill_1  FILLER_66_840
timestamp 1677579658
transform 1 0 152256 0 1 121716
box -48 -56 144 834
use sg13g2_decap_8  FILLER_67_0
timestamp 1679581782
transform 1 0 71616 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_7
timestamp 1679581782
transform 1 0 72288 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_14
timestamp 1679581782
transform 1 0 72960 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_21
timestamp 1679581782
transform 1 0 73632 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_28
timestamp 1679581782
transform 1 0 74304 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_35
timestamp 1679581782
transform 1 0 74976 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_42
timestamp 1679581782
transform 1 0 75648 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_49
timestamp 1679581782
transform 1 0 76320 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_56
timestamp 1679581782
transform 1 0 76992 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_63
timestamp 1679581782
transform 1 0 77664 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_70
timestamp 1679581782
transform 1 0 78336 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_77
timestamp 1679581782
transform 1 0 79008 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_84
timestamp 1679581782
transform 1 0 79680 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_91
timestamp 1679581782
transform 1 0 80352 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_98
timestamp 1679581782
transform 1 0 81024 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_105
timestamp 1679581782
transform 1 0 81696 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_112
timestamp 1679581782
transform 1 0 82368 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_119
timestamp 1679581782
transform 1 0 83040 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_126
timestamp 1679581782
transform 1 0 83712 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_133
timestamp 1679581782
transform 1 0 84384 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_140
timestamp 1679581782
transform 1 0 85056 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_147
timestamp 1679581782
transform 1 0 85728 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_154
timestamp 1679581782
transform 1 0 86400 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_161
timestamp 1679581782
transform 1 0 87072 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_168
timestamp 1679581782
transform 1 0 87744 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_175
timestamp 1679581782
transform 1 0 88416 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_182
timestamp 1679581782
transform 1 0 89088 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_189
timestamp 1679581782
transform 1 0 89760 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_196
timestamp 1679581782
transform 1 0 90432 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_203
timestamp 1679581782
transform 1 0 91104 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_210
timestamp 1679581782
transform 1 0 91776 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_217
timestamp 1679581782
transform 1 0 92448 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_224
timestamp 1679581782
transform 1 0 93120 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_231
timestamp 1679581782
transform 1 0 93792 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_238
timestamp 1679581782
transform 1 0 94464 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_245
timestamp 1679581782
transform 1 0 95136 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_252
timestamp 1679581782
transform 1 0 95808 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_259
timestamp 1679581782
transform 1 0 96480 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_266
timestamp 1679581782
transform 1 0 97152 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_273
timestamp 1679581782
transform 1 0 97824 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_280
timestamp 1679581782
transform 1 0 98496 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_287
timestamp 1679581782
transform 1 0 99168 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_294
timestamp 1679581782
transform 1 0 99840 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_301
timestamp 1679581782
transform 1 0 100512 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_308
timestamp 1679581782
transform 1 0 101184 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_315
timestamp 1679581782
transform 1 0 101856 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_322
timestamp 1679581782
transform 1 0 102528 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_329
timestamp 1679581782
transform 1 0 103200 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_336
timestamp 1679581782
transform 1 0 103872 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_343
timestamp 1679581782
transform 1 0 104544 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_350
timestamp 1679581782
transform 1 0 105216 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_357
timestamp 1679581782
transform 1 0 105888 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_364
timestamp 1679581782
transform 1 0 106560 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_371
timestamp 1679581782
transform 1 0 107232 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_378
timestamp 1679581782
transform 1 0 107904 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_385
timestamp 1679581782
transform 1 0 108576 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_392
timestamp 1679581782
transform 1 0 109248 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_399
timestamp 1679581782
transform 1 0 109920 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_406
timestamp 1679581782
transform 1 0 110592 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_413
timestamp 1679581782
transform 1 0 111264 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_420
timestamp 1679581782
transform 1 0 111936 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_427
timestamp 1679581782
transform 1 0 112608 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_434
timestamp 1679581782
transform 1 0 113280 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_441
timestamp 1679581782
transform 1 0 113952 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_448
timestamp 1679581782
transform 1 0 114624 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_455
timestamp 1679581782
transform 1 0 115296 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_462
timestamp 1679581782
transform 1 0 115968 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_469
timestamp 1679581782
transform 1 0 116640 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_476
timestamp 1679581782
transform 1 0 117312 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_483
timestamp 1679581782
transform 1 0 117984 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_490
timestamp 1679581782
transform 1 0 118656 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_497
timestamp 1679581782
transform 1 0 119328 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_504
timestamp 1679581782
transform 1 0 120000 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_511
timestamp 1679581782
transform 1 0 120672 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_518
timestamp 1679581782
transform 1 0 121344 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_525
timestamp 1679581782
transform 1 0 122016 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_532
timestamp 1679581782
transform 1 0 122688 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_539
timestamp 1679581782
transform 1 0 123360 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_546
timestamp 1679581782
transform 1 0 124032 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_553
timestamp 1679581782
transform 1 0 124704 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_560
timestamp 1679581782
transform 1 0 125376 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_567
timestamp 1679581782
transform 1 0 126048 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_574
timestamp 1679581782
transform 1 0 126720 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_581
timestamp 1679581782
transform 1 0 127392 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_588
timestamp 1679581782
transform 1 0 128064 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_595
timestamp 1679581782
transform 1 0 128736 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_602
timestamp 1679581782
transform 1 0 129408 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_609
timestamp 1679581782
transform 1 0 130080 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_616
timestamp 1679581782
transform 1 0 130752 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_623
timestamp 1679581782
transform 1 0 131424 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_630
timestamp 1679581782
transform 1 0 132096 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_637
timestamp 1679581782
transform 1 0 132768 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_644
timestamp 1679581782
transform 1 0 133440 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_651
timestamp 1679581782
transform 1 0 134112 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_658
timestamp 1679581782
transform 1 0 134784 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_665
timestamp 1679581782
transform 1 0 135456 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_672
timestamp 1679581782
transform 1 0 136128 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_679
timestamp 1679581782
transform 1 0 136800 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_686
timestamp 1679581782
transform 1 0 137472 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_693
timestamp 1679581782
transform 1 0 138144 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_700
timestamp 1679581782
transform 1 0 138816 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_707
timestamp 1679581782
transform 1 0 139488 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_714
timestamp 1679581782
transform 1 0 140160 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_721
timestamp 1679581782
transform 1 0 140832 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_728
timestamp 1679581782
transform 1 0 141504 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_735
timestamp 1679581782
transform 1 0 142176 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_742
timestamp 1679581782
transform 1 0 142848 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_749
timestamp 1679581782
transform 1 0 143520 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_756
timestamp 1679581782
transform 1 0 144192 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_763
timestamp 1679581782
transform 1 0 144864 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_770
timestamp 1679581782
transform 1 0 145536 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_777
timestamp 1679581782
transform 1 0 146208 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_784
timestamp 1679581782
transform 1 0 146880 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_791
timestamp 1679581782
transform 1 0 147552 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_798
timestamp 1679581782
transform 1 0 148224 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_805
timestamp 1679581782
transform 1 0 148896 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_812
timestamp 1679581782
transform 1 0 149568 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_819
timestamp 1679581782
transform 1 0 150240 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_826
timestamp 1679581782
transform 1 0 150912 0 -1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_833
timestamp 1679581782
transform 1 0 151584 0 -1 123228
box -48 -56 720 834
use sg13g2_fill_1  FILLER_67_840
timestamp 1677579658
transform 1 0 152256 0 -1 123228
box -48 -56 144 834
use sg13g2_decap_8  FILLER_68_0
timestamp 1679581782
transform 1 0 71616 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_7
timestamp 1679581782
transform 1 0 72288 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_14
timestamp 1679581782
transform 1 0 72960 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_21
timestamp 1679581782
transform 1 0 73632 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_28
timestamp 1679581782
transform 1 0 74304 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_35
timestamp 1679581782
transform 1 0 74976 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_42
timestamp 1679581782
transform 1 0 75648 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_49
timestamp 1679581782
transform 1 0 76320 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_56
timestamp 1679581782
transform 1 0 76992 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_63
timestamp 1679581782
transform 1 0 77664 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_70
timestamp 1679581782
transform 1 0 78336 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_77
timestamp 1679581782
transform 1 0 79008 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_84
timestamp 1679581782
transform 1 0 79680 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_91
timestamp 1679581782
transform 1 0 80352 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_98
timestamp 1679581782
transform 1 0 81024 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_105
timestamp 1679581782
transform 1 0 81696 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_112
timestamp 1679581782
transform 1 0 82368 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_119
timestamp 1679581782
transform 1 0 83040 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_126
timestamp 1679581782
transform 1 0 83712 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_133
timestamp 1679581782
transform 1 0 84384 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_140
timestamp 1679581782
transform 1 0 85056 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_147
timestamp 1679581782
transform 1 0 85728 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_154
timestamp 1679581782
transform 1 0 86400 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_161
timestamp 1679581782
transform 1 0 87072 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_168
timestamp 1679581782
transform 1 0 87744 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_175
timestamp 1679581782
transform 1 0 88416 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_182
timestamp 1679581782
transform 1 0 89088 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_189
timestamp 1679581782
transform 1 0 89760 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_196
timestamp 1679581782
transform 1 0 90432 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_203
timestamp 1679581782
transform 1 0 91104 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_210
timestamp 1679581782
transform 1 0 91776 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_217
timestamp 1679581782
transform 1 0 92448 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_224
timestamp 1679581782
transform 1 0 93120 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_231
timestamp 1679581782
transform 1 0 93792 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_238
timestamp 1679581782
transform 1 0 94464 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_245
timestamp 1679581782
transform 1 0 95136 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_252
timestamp 1679581782
transform 1 0 95808 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_259
timestamp 1679581782
transform 1 0 96480 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_266
timestamp 1679581782
transform 1 0 97152 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_273
timestamp 1679581782
transform 1 0 97824 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_280
timestamp 1679581782
transform 1 0 98496 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_287
timestamp 1679581782
transform 1 0 99168 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_294
timestamp 1679581782
transform 1 0 99840 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_301
timestamp 1679581782
transform 1 0 100512 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_308
timestamp 1679581782
transform 1 0 101184 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_315
timestamp 1679581782
transform 1 0 101856 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_322
timestamp 1679581782
transform 1 0 102528 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_329
timestamp 1679581782
transform 1 0 103200 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_336
timestamp 1679581782
transform 1 0 103872 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_343
timestamp 1679581782
transform 1 0 104544 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_350
timestamp 1679581782
transform 1 0 105216 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_357
timestamp 1679581782
transform 1 0 105888 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_364
timestamp 1679581782
transform 1 0 106560 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_371
timestamp 1679581782
transform 1 0 107232 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_378
timestamp 1679581782
transform 1 0 107904 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_385
timestamp 1679581782
transform 1 0 108576 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_392
timestamp 1679581782
transform 1 0 109248 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_399
timestamp 1679581782
transform 1 0 109920 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_406
timestamp 1679581782
transform 1 0 110592 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_413
timestamp 1679581782
transform 1 0 111264 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_420
timestamp 1679581782
transform 1 0 111936 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_427
timestamp 1679581782
transform 1 0 112608 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_434
timestamp 1679581782
transform 1 0 113280 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_441
timestamp 1679581782
transform 1 0 113952 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_448
timestamp 1679581782
transform 1 0 114624 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_455
timestamp 1679581782
transform 1 0 115296 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_462
timestamp 1679581782
transform 1 0 115968 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_469
timestamp 1679581782
transform 1 0 116640 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_476
timestamp 1679581782
transform 1 0 117312 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_483
timestamp 1679581782
transform 1 0 117984 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_490
timestamp 1679581782
transform 1 0 118656 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_497
timestamp 1679581782
transform 1 0 119328 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_504
timestamp 1679581782
transform 1 0 120000 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_511
timestamp 1679581782
transform 1 0 120672 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_518
timestamp 1679581782
transform 1 0 121344 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_525
timestamp 1679581782
transform 1 0 122016 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_532
timestamp 1679581782
transform 1 0 122688 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_539
timestamp 1679581782
transform 1 0 123360 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_546
timestamp 1679581782
transform 1 0 124032 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_553
timestamp 1679581782
transform 1 0 124704 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_560
timestamp 1679581782
transform 1 0 125376 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_567
timestamp 1679581782
transform 1 0 126048 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_574
timestamp 1679581782
transform 1 0 126720 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_581
timestamp 1679581782
transform 1 0 127392 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_588
timestamp 1679581782
transform 1 0 128064 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_595
timestamp 1679581782
transform 1 0 128736 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_602
timestamp 1679581782
transform 1 0 129408 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_609
timestamp 1679581782
transform 1 0 130080 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_616
timestamp 1679581782
transform 1 0 130752 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_623
timestamp 1679581782
transform 1 0 131424 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_630
timestamp 1679581782
transform 1 0 132096 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_637
timestamp 1679581782
transform 1 0 132768 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_644
timestamp 1679581782
transform 1 0 133440 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_651
timestamp 1679581782
transform 1 0 134112 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_658
timestamp 1679581782
transform 1 0 134784 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_665
timestamp 1679581782
transform 1 0 135456 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_672
timestamp 1679581782
transform 1 0 136128 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_679
timestamp 1679581782
transform 1 0 136800 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_686
timestamp 1679581782
transform 1 0 137472 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_693
timestamp 1679581782
transform 1 0 138144 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_700
timestamp 1679581782
transform 1 0 138816 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_707
timestamp 1679581782
transform 1 0 139488 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_714
timestamp 1679581782
transform 1 0 140160 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_721
timestamp 1679581782
transform 1 0 140832 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_728
timestamp 1679581782
transform 1 0 141504 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_735
timestamp 1679581782
transform 1 0 142176 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_742
timestamp 1679581782
transform 1 0 142848 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_749
timestamp 1679581782
transform 1 0 143520 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_756
timestamp 1679581782
transform 1 0 144192 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_763
timestamp 1679581782
transform 1 0 144864 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_770
timestamp 1679581782
transform 1 0 145536 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_777
timestamp 1679581782
transform 1 0 146208 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_784
timestamp 1679581782
transform 1 0 146880 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_791
timestamp 1679581782
transform 1 0 147552 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_798
timestamp 1679581782
transform 1 0 148224 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_805
timestamp 1679581782
transform 1 0 148896 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_812
timestamp 1679581782
transform 1 0 149568 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_819
timestamp 1679581782
transform 1 0 150240 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_826
timestamp 1679581782
transform 1 0 150912 0 1 123228
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_833
timestamp 1679581782
transform 1 0 151584 0 1 123228
box -48 -56 720 834
use sg13g2_fill_1  FILLER_68_840
timestamp 1677579658
transform 1 0 152256 0 1 123228
box -48 -56 144 834
use sg13g2_decap_8  FILLER_69_0
timestamp 1679581782
transform 1 0 71616 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_7
timestamp 1679581782
transform 1 0 72288 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_14
timestamp 1679581782
transform 1 0 72960 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_21
timestamp 1679581782
transform 1 0 73632 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_28
timestamp 1679581782
transform 1 0 74304 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_35
timestamp 1679581782
transform 1 0 74976 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_42
timestamp 1679581782
transform 1 0 75648 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_49
timestamp 1679581782
transform 1 0 76320 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_56
timestamp 1679581782
transform 1 0 76992 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_63
timestamp 1679581782
transform 1 0 77664 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_70
timestamp 1679581782
transform 1 0 78336 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_77
timestamp 1679581782
transform 1 0 79008 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_84
timestamp 1679581782
transform 1 0 79680 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_91
timestamp 1679581782
transform 1 0 80352 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_98
timestamp 1679581782
transform 1 0 81024 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_105
timestamp 1679581782
transform 1 0 81696 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_112
timestamp 1679581782
transform 1 0 82368 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_119
timestamp 1679581782
transform 1 0 83040 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_126
timestamp 1679581782
transform 1 0 83712 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_133
timestamp 1679581782
transform 1 0 84384 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_140
timestamp 1679581782
transform 1 0 85056 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_147
timestamp 1679581782
transform 1 0 85728 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_154
timestamp 1679581782
transform 1 0 86400 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_161
timestamp 1679581782
transform 1 0 87072 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_168
timestamp 1679581782
transform 1 0 87744 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_175
timestamp 1679581782
transform 1 0 88416 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_182
timestamp 1679581782
transform 1 0 89088 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_189
timestamp 1679581782
transform 1 0 89760 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_196
timestamp 1679581782
transform 1 0 90432 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_203
timestamp 1679581782
transform 1 0 91104 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_210
timestamp 1679581782
transform 1 0 91776 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_217
timestamp 1679581782
transform 1 0 92448 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_224
timestamp 1679581782
transform 1 0 93120 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_231
timestamp 1679581782
transform 1 0 93792 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_238
timestamp 1679581782
transform 1 0 94464 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_245
timestamp 1679581782
transform 1 0 95136 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_252
timestamp 1679581782
transform 1 0 95808 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_259
timestamp 1679581782
transform 1 0 96480 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_266
timestamp 1679581782
transform 1 0 97152 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_273
timestamp 1679581782
transform 1 0 97824 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_280
timestamp 1679581782
transform 1 0 98496 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_287
timestamp 1679581782
transform 1 0 99168 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_294
timestamp 1679581782
transform 1 0 99840 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_301
timestamp 1679581782
transform 1 0 100512 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_308
timestamp 1679581782
transform 1 0 101184 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_315
timestamp 1679581782
transform 1 0 101856 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_322
timestamp 1679581782
transform 1 0 102528 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_329
timestamp 1679581782
transform 1 0 103200 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_336
timestamp 1679581782
transform 1 0 103872 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_343
timestamp 1679581782
transform 1 0 104544 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_350
timestamp 1679581782
transform 1 0 105216 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_357
timestamp 1679581782
transform 1 0 105888 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_364
timestamp 1679581782
transform 1 0 106560 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_371
timestamp 1679581782
transform 1 0 107232 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_378
timestamp 1679581782
transform 1 0 107904 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_385
timestamp 1679581782
transform 1 0 108576 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_392
timestamp 1679581782
transform 1 0 109248 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_399
timestamp 1679581782
transform 1 0 109920 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_406
timestamp 1679581782
transform 1 0 110592 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_413
timestamp 1679581782
transform 1 0 111264 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_420
timestamp 1679581782
transform 1 0 111936 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_427
timestamp 1679581782
transform 1 0 112608 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_434
timestamp 1679581782
transform 1 0 113280 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_441
timestamp 1679581782
transform 1 0 113952 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_448
timestamp 1679581782
transform 1 0 114624 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_455
timestamp 1679581782
transform 1 0 115296 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_462
timestamp 1679581782
transform 1 0 115968 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_469
timestamp 1679581782
transform 1 0 116640 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_476
timestamp 1679581782
transform 1 0 117312 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_483
timestamp 1679581782
transform 1 0 117984 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_490
timestamp 1679581782
transform 1 0 118656 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_497
timestamp 1679581782
transform 1 0 119328 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_504
timestamp 1679581782
transform 1 0 120000 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_511
timestamp 1679581782
transform 1 0 120672 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_518
timestamp 1679581782
transform 1 0 121344 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_525
timestamp 1679581782
transform 1 0 122016 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_532
timestamp 1679581782
transform 1 0 122688 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_539
timestamp 1679581782
transform 1 0 123360 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_546
timestamp 1679581782
transform 1 0 124032 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_553
timestamp 1679581782
transform 1 0 124704 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_560
timestamp 1679581782
transform 1 0 125376 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_567
timestamp 1679581782
transform 1 0 126048 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_574
timestamp 1679581782
transform 1 0 126720 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_581
timestamp 1679581782
transform 1 0 127392 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_588
timestamp 1679581782
transform 1 0 128064 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_595
timestamp 1679581782
transform 1 0 128736 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_602
timestamp 1679581782
transform 1 0 129408 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_609
timestamp 1679581782
transform 1 0 130080 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_616
timestamp 1679581782
transform 1 0 130752 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_623
timestamp 1679581782
transform 1 0 131424 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_630
timestamp 1679581782
transform 1 0 132096 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_637
timestamp 1679581782
transform 1 0 132768 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_644
timestamp 1679581782
transform 1 0 133440 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_651
timestamp 1679581782
transform 1 0 134112 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_658
timestamp 1679581782
transform 1 0 134784 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_665
timestamp 1679581782
transform 1 0 135456 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_672
timestamp 1679581782
transform 1 0 136128 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_679
timestamp 1679581782
transform 1 0 136800 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_686
timestamp 1679581782
transform 1 0 137472 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_693
timestamp 1679581782
transform 1 0 138144 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_700
timestamp 1679581782
transform 1 0 138816 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_707
timestamp 1679581782
transform 1 0 139488 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_714
timestamp 1679581782
transform 1 0 140160 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_721
timestamp 1679581782
transform 1 0 140832 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_728
timestamp 1679581782
transform 1 0 141504 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_735
timestamp 1679581782
transform 1 0 142176 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_742
timestamp 1679581782
transform 1 0 142848 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_749
timestamp 1679581782
transform 1 0 143520 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_756
timestamp 1679581782
transform 1 0 144192 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_763
timestamp 1679581782
transform 1 0 144864 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_770
timestamp 1679581782
transform 1 0 145536 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_777
timestamp 1679581782
transform 1 0 146208 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_784
timestamp 1679581782
transform 1 0 146880 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_791
timestamp 1679581782
transform 1 0 147552 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_798
timestamp 1679581782
transform 1 0 148224 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_805
timestamp 1679581782
transform 1 0 148896 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_812
timestamp 1679581782
transform 1 0 149568 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_819
timestamp 1679581782
transform 1 0 150240 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_826
timestamp 1679581782
transform 1 0 150912 0 -1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_833
timestamp 1679581782
transform 1 0 151584 0 -1 124740
box -48 -56 720 834
use sg13g2_fill_1  FILLER_69_840
timestamp 1677579658
transform 1 0 152256 0 -1 124740
box -48 -56 144 834
use sg13g2_decap_8  FILLER_70_0
timestamp 1679581782
transform 1 0 71616 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_7
timestamp 1679581782
transform 1 0 72288 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_14
timestamp 1679581782
transform 1 0 72960 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_21
timestamp 1679581782
transform 1 0 73632 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_28
timestamp 1679581782
transform 1 0 74304 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_35
timestamp 1679581782
transform 1 0 74976 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_42
timestamp 1679581782
transform 1 0 75648 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_49
timestamp 1679581782
transform 1 0 76320 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_56
timestamp 1679581782
transform 1 0 76992 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_63
timestamp 1679581782
transform 1 0 77664 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_70
timestamp 1679581782
transform 1 0 78336 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_77
timestamp 1679581782
transform 1 0 79008 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_84
timestamp 1679581782
transform 1 0 79680 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_91
timestamp 1679581782
transform 1 0 80352 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_98
timestamp 1679581782
transform 1 0 81024 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_105
timestamp 1679581782
transform 1 0 81696 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_112
timestamp 1679581782
transform 1 0 82368 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_119
timestamp 1679581782
transform 1 0 83040 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_126
timestamp 1679581782
transform 1 0 83712 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_133
timestamp 1679581782
transform 1 0 84384 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_140
timestamp 1679581782
transform 1 0 85056 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_147
timestamp 1679581782
transform 1 0 85728 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_154
timestamp 1679581782
transform 1 0 86400 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_161
timestamp 1679581782
transform 1 0 87072 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_168
timestamp 1679581782
transform 1 0 87744 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_175
timestamp 1679581782
transform 1 0 88416 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_182
timestamp 1679581782
transform 1 0 89088 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_189
timestamp 1679581782
transform 1 0 89760 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_196
timestamp 1679581782
transform 1 0 90432 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_203
timestamp 1679581782
transform 1 0 91104 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_210
timestamp 1679581782
transform 1 0 91776 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_217
timestamp 1679581782
transform 1 0 92448 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_224
timestamp 1679581782
transform 1 0 93120 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_231
timestamp 1679581782
transform 1 0 93792 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_238
timestamp 1679581782
transform 1 0 94464 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_245
timestamp 1679581782
transform 1 0 95136 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_252
timestamp 1679581782
transform 1 0 95808 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_259
timestamp 1679581782
transform 1 0 96480 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_266
timestamp 1679581782
transform 1 0 97152 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_273
timestamp 1679581782
transform 1 0 97824 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_280
timestamp 1679581782
transform 1 0 98496 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_287
timestamp 1679581782
transform 1 0 99168 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_294
timestamp 1679581782
transform 1 0 99840 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_301
timestamp 1679581782
transform 1 0 100512 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_308
timestamp 1679581782
transform 1 0 101184 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_315
timestamp 1679581782
transform 1 0 101856 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_322
timestamp 1679581782
transform 1 0 102528 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_329
timestamp 1679581782
transform 1 0 103200 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_336
timestamp 1679581782
transform 1 0 103872 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_343
timestamp 1679581782
transform 1 0 104544 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_350
timestamp 1679581782
transform 1 0 105216 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_357
timestamp 1679581782
transform 1 0 105888 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_364
timestamp 1679581782
transform 1 0 106560 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_371
timestamp 1679581782
transform 1 0 107232 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_378
timestamp 1679581782
transform 1 0 107904 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_385
timestamp 1679581782
transform 1 0 108576 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_392
timestamp 1679581782
transform 1 0 109248 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_399
timestamp 1679581782
transform 1 0 109920 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_406
timestamp 1679581782
transform 1 0 110592 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_413
timestamp 1679581782
transform 1 0 111264 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_420
timestamp 1679581782
transform 1 0 111936 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_427
timestamp 1679581782
transform 1 0 112608 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_434
timestamp 1679581782
transform 1 0 113280 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_441
timestamp 1679581782
transform 1 0 113952 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_448
timestamp 1679581782
transform 1 0 114624 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_455
timestamp 1679581782
transform 1 0 115296 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_462
timestamp 1679581782
transform 1 0 115968 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_469
timestamp 1679581782
transform 1 0 116640 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_476
timestamp 1679581782
transform 1 0 117312 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_483
timestamp 1679581782
transform 1 0 117984 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_490
timestamp 1679581782
transform 1 0 118656 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_497
timestamp 1679581782
transform 1 0 119328 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_504
timestamp 1679581782
transform 1 0 120000 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_511
timestamp 1679581782
transform 1 0 120672 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_518
timestamp 1679581782
transform 1 0 121344 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_525
timestamp 1679581782
transform 1 0 122016 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_532
timestamp 1679581782
transform 1 0 122688 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_539
timestamp 1679581782
transform 1 0 123360 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_546
timestamp 1679581782
transform 1 0 124032 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_553
timestamp 1679581782
transform 1 0 124704 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_560
timestamp 1679581782
transform 1 0 125376 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_567
timestamp 1679581782
transform 1 0 126048 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_574
timestamp 1679581782
transform 1 0 126720 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_581
timestamp 1679581782
transform 1 0 127392 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_588
timestamp 1679581782
transform 1 0 128064 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_595
timestamp 1679581782
transform 1 0 128736 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_602
timestamp 1679581782
transform 1 0 129408 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_609
timestamp 1679581782
transform 1 0 130080 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_616
timestamp 1679581782
transform 1 0 130752 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_623
timestamp 1679581782
transform 1 0 131424 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_630
timestamp 1679581782
transform 1 0 132096 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_637
timestamp 1679581782
transform 1 0 132768 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_644
timestamp 1679581782
transform 1 0 133440 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_651
timestamp 1679581782
transform 1 0 134112 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_658
timestamp 1679581782
transform 1 0 134784 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_665
timestamp 1679581782
transform 1 0 135456 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_672
timestamp 1679581782
transform 1 0 136128 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_679
timestamp 1679581782
transform 1 0 136800 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_686
timestamp 1679581782
transform 1 0 137472 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_693
timestamp 1679581782
transform 1 0 138144 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_700
timestamp 1679581782
transform 1 0 138816 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_707
timestamp 1679581782
transform 1 0 139488 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_714
timestamp 1679581782
transform 1 0 140160 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_721
timestamp 1679581782
transform 1 0 140832 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_728
timestamp 1679581782
transform 1 0 141504 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_735
timestamp 1679581782
transform 1 0 142176 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_742
timestamp 1679581782
transform 1 0 142848 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_749
timestamp 1679581782
transform 1 0 143520 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_756
timestamp 1679581782
transform 1 0 144192 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_763
timestamp 1679581782
transform 1 0 144864 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_770
timestamp 1679581782
transform 1 0 145536 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_777
timestamp 1679581782
transform 1 0 146208 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_784
timestamp 1679581782
transform 1 0 146880 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_791
timestamp 1679581782
transform 1 0 147552 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_798
timestamp 1679581782
transform 1 0 148224 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_805
timestamp 1679581782
transform 1 0 148896 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_812
timestamp 1679581782
transform 1 0 149568 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_819
timestamp 1679581782
transform 1 0 150240 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_826
timestamp 1679581782
transform 1 0 150912 0 1 124740
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_833
timestamp 1679581782
transform 1 0 151584 0 1 124740
box -48 -56 720 834
use sg13g2_fill_1  FILLER_70_840
timestamp 1677579658
transform 1 0 152256 0 1 124740
box -48 -56 144 834
use sg13g2_decap_8  FILLER_71_0
timestamp 1679581782
transform 1 0 71616 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_7
timestamp 1679581782
transform 1 0 72288 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_14
timestamp 1679581782
transform 1 0 72960 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_21
timestamp 1679581782
transform 1 0 73632 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_28
timestamp 1679581782
transform 1 0 74304 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_35
timestamp 1679581782
transform 1 0 74976 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_42
timestamp 1679581782
transform 1 0 75648 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_49
timestamp 1679581782
transform 1 0 76320 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_56
timestamp 1679581782
transform 1 0 76992 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_63
timestamp 1679581782
transform 1 0 77664 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_70
timestamp 1679581782
transform 1 0 78336 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_77
timestamp 1679581782
transform 1 0 79008 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_84
timestamp 1679581782
transform 1 0 79680 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_91
timestamp 1679581782
transform 1 0 80352 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_98
timestamp 1679581782
transform 1 0 81024 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_105
timestamp 1679581782
transform 1 0 81696 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_112
timestamp 1679581782
transform 1 0 82368 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_119
timestamp 1679581782
transform 1 0 83040 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_126
timestamp 1679581782
transform 1 0 83712 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_133
timestamp 1679581782
transform 1 0 84384 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_140
timestamp 1679581782
transform 1 0 85056 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_147
timestamp 1679581782
transform 1 0 85728 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_154
timestamp 1679581782
transform 1 0 86400 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_161
timestamp 1679581782
transform 1 0 87072 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_168
timestamp 1679581782
transform 1 0 87744 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_175
timestamp 1679581782
transform 1 0 88416 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_182
timestamp 1679581782
transform 1 0 89088 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_189
timestamp 1679581782
transform 1 0 89760 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_196
timestamp 1679581782
transform 1 0 90432 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_203
timestamp 1679581782
transform 1 0 91104 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_210
timestamp 1679581782
transform 1 0 91776 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_217
timestamp 1679581782
transform 1 0 92448 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_224
timestamp 1679581782
transform 1 0 93120 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_231
timestamp 1679581782
transform 1 0 93792 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_238
timestamp 1679581782
transform 1 0 94464 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_245
timestamp 1679581782
transform 1 0 95136 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_252
timestamp 1679581782
transform 1 0 95808 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_259
timestamp 1679581782
transform 1 0 96480 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_266
timestamp 1679581782
transform 1 0 97152 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_273
timestamp 1679581782
transform 1 0 97824 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_280
timestamp 1679581782
transform 1 0 98496 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_287
timestamp 1679581782
transform 1 0 99168 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_294
timestamp 1679581782
transform 1 0 99840 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_301
timestamp 1679581782
transform 1 0 100512 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_308
timestamp 1679581782
transform 1 0 101184 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_315
timestamp 1679581782
transform 1 0 101856 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_322
timestamp 1679581782
transform 1 0 102528 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_329
timestamp 1679581782
transform 1 0 103200 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_336
timestamp 1679581782
transform 1 0 103872 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_343
timestamp 1679581782
transform 1 0 104544 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_350
timestamp 1679581782
transform 1 0 105216 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_357
timestamp 1679581782
transform 1 0 105888 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_364
timestamp 1679581782
transform 1 0 106560 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_371
timestamp 1679581782
transform 1 0 107232 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_378
timestamp 1679581782
transform 1 0 107904 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_385
timestamp 1679581782
transform 1 0 108576 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_392
timestamp 1679581782
transform 1 0 109248 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_399
timestamp 1679581782
transform 1 0 109920 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_406
timestamp 1679581782
transform 1 0 110592 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_413
timestamp 1679581782
transform 1 0 111264 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_420
timestamp 1679581782
transform 1 0 111936 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_427
timestamp 1679581782
transform 1 0 112608 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_434
timestamp 1679581782
transform 1 0 113280 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_441
timestamp 1679581782
transform 1 0 113952 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_448
timestamp 1679581782
transform 1 0 114624 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_455
timestamp 1679581782
transform 1 0 115296 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_462
timestamp 1679581782
transform 1 0 115968 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_469
timestamp 1679581782
transform 1 0 116640 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_476
timestamp 1679581782
transform 1 0 117312 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_483
timestamp 1679581782
transform 1 0 117984 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_490
timestamp 1679581782
transform 1 0 118656 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_497
timestamp 1679581782
transform 1 0 119328 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_504
timestamp 1679581782
transform 1 0 120000 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_511
timestamp 1679581782
transform 1 0 120672 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_518
timestamp 1679581782
transform 1 0 121344 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_525
timestamp 1679581782
transform 1 0 122016 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_532
timestamp 1679581782
transform 1 0 122688 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_539
timestamp 1679581782
transform 1 0 123360 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_546
timestamp 1679581782
transform 1 0 124032 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_553
timestamp 1679581782
transform 1 0 124704 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_560
timestamp 1679581782
transform 1 0 125376 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_567
timestamp 1679581782
transform 1 0 126048 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_574
timestamp 1679581782
transform 1 0 126720 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_581
timestamp 1679581782
transform 1 0 127392 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_588
timestamp 1679581782
transform 1 0 128064 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_595
timestamp 1679581782
transform 1 0 128736 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_602
timestamp 1679581782
transform 1 0 129408 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_609
timestamp 1679581782
transform 1 0 130080 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_616
timestamp 1679581782
transform 1 0 130752 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_623
timestamp 1679581782
transform 1 0 131424 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_630
timestamp 1679581782
transform 1 0 132096 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_637
timestamp 1679581782
transform 1 0 132768 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_644
timestamp 1679581782
transform 1 0 133440 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_651
timestamp 1679581782
transform 1 0 134112 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_658
timestamp 1679581782
transform 1 0 134784 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_665
timestamp 1679581782
transform 1 0 135456 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_672
timestamp 1679581782
transform 1 0 136128 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_679
timestamp 1679581782
transform 1 0 136800 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_686
timestamp 1679581782
transform 1 0 137472 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_693
timestamp 1679581782
transform 1 0 138144 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_700
timestamp 1679581782
transform 1 0 138816 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_707
timestamp 1679581782
transform 1 0 139488 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_714
timestamp 1679581782
transform 1 0 140160 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_721
timestamp 1679581782
transform 1 0 140832 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_728
timestamp 1679581782
transform 1 0 141504 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_735
timestamp 1679581782
transform 1 0 142176 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_742
timestamp 1679581782
transform 1 0 142848 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_749
timestamp 1679581782
transform 1 0 143520 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_756
timestamp 1679581782
transform 1 0 144192 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_763
timestamp 1679581782
transform 1 0 144864 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_770
timestamp 1679581782
transform 1 0 145536 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_777
timestamp 1679581782
transform 1 0 146208 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_784
timestamp 1679581782
transform 1 0 146880 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_791
timestamp 1679581782
transform 1 0 147552 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_798
timestamp 1679581782
transform 1 0 148224 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_805
timestamp 1679581782
transform 1 0 148896 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_812
timestamp 1679581782
transform 1 0 149568 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_819
timestamp 1679581782
transform 1 0 150240 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_826
timestamp 1679581782
transform 1 0 150912 0 -1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_833
timestamp 1679581782
transform 1 0 151584 0 -1 126252
box -48 -56 720 834
use sg13g2_fill_1  FILLER_71_840
timestamp 1677579658
transform 1 0 152256 0 -1 126252
box -48 -56 144 834
use sg13g2_decap_8  FILLER_72_0
timestamp 1679581782
transform 1 0 71616 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_7
timestamp 1679581782
transform 1 0 72288 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_14
timestamp 1679581782
transform 1 0 72960 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_21
timestamp 1679581782
transform 1 0 73632 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_28
timestamp 1679581782
transform 1 0 74304 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_35
timestamp 1679581782
transform 1 0 74976 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_42
timestamp 1679581782
transform 1 0 75648 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_49
timestamp 1679581782
transform 1 0 76320 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_56
timestamp 1679581782
transform 1 0 76992 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_63
timestamp 1679581782
transform 1 0 77664 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_70
timestamp 1679581782
transform 1 0 78336 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_77
timestamp 1679581782
transform 1 0 79008 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_84
timestamp 1679581782
transform 1 0 79680 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_91
timestamp 1679581782
transform 1 0 80352 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_98
timestamp 1679581782
transform 1 0 81024 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_105
timestamp 1679581782
transform 1 0 81696 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_112
timestamp 1679581782
transform 1 0 82368 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_119
timestamp 1679581782
transform 1 0 83040 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_126
timestamp 1679581782
transform 1 0 83712 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_133
timestamp 1679581782
transform 1 0 84384 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_140
timestamp 1679581782
transform 1 0 85056 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_147
timestamp 1679581782
transform 1 0 85728 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_154
timestamp 1679581782
transform 1 0 86400 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_161
timestamp 1679581782
transform 1 0 87072 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_168
timestamp 1679581782
transform 1 0 87744 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_175
timestamp 1679581782
transform 1 0 88416 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_182
timestamp 1679581782
transform 1 0 89088 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_189
timestamp 1679581782
transform 1 0 89760 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_196
timestamp 1679581782
transform 1 0 90432 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_203
timestamp 1679581782
transform 1 0 91104 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_210
timestamp 1679581782
transform 1 0 91776 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_217
timestamp 1679581782
transform 1 0 92448 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_224
timestamp 1679581782
transform 1 0 93120 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_231
timestamp 1679581782
transform 1 0 93792 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_238
timestamp 1679581782
transform 1 0 94464 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_245
timestamp 1679581782
transform 1 0 95136 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_252
timestamp 1679581782
transform 1 0 95808 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_259
timestamp 1679581782
transform 1 0 96480 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_266
timestamp 1679581782
transform 1 0 97152 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_273
timestamp 1679581782
transform 1 0 97824 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_280
timestamp 1679581782
transform 1 0 98496 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_287
timestamp 1679581782
transform 1 0 99168 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_294
timestamp 1679581782
transform 1 0 99840 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_301
timestamp 1679581782
transform 1 0 100512 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_308
timestamp 1679581782
transform 1 0 101184 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_315
timestamp 1679581782
transform 1 0 101856 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_322
timestamp 1679581782
transform 1 0 102528 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_329
timestamp 1679581782
transform 1 0 103200 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_336
timestamp 1679581782
transform 1 0 103872 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_343
timestamp 1679581782
transform 1 0 104544 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_350
timestamp 1679581782
transform 1 0 105216 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_357
timestamp 1679581782
transform 1 0 105888 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_364
timestamp 1679581782
transform 1 0 106560 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_371
timestamp 1679581782
transform 1 0 107232 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_378
timestamp 1679581782
transform 1 0 107904 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_385
timestamp 1679581782
transform 1 0 108576 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_392
timestamp 1679581782
transform 1 0 109248 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_399
timestamp 1679581782
transform 1 0 109920 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_406
timestamp 1679581782
transform 1 0 110592 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_413
timestamp 1679581782
transform 1 0 111264 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_420
timestamp 1679581782
transform 1 0 111936 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_427
timestamp 1679581782
transform 1 0 112608 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_434
timestamp 1679581782
transform 1 0 113280 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_441
timestamp 1679581782
transform 1 0 113952 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_448
timestamp 1679581782
transform 1 0 114624 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_455
timestamp 1679581782
transform 1 0 115296 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_462
timestamp 1679581782
transform 1 0 115968 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_469
timestamp 1679581782
transform 1 0 116640 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_476
timestamp 1679581782
transform 1 0 117312 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_483
timestamp 1679581782
transform 1 0 117984 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_490
timestamp 1679581782
transform 1 0 118656 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_497
timestamp 1679581782
transform 1 0 119328 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_504
timestamp 1679581782
transform 1 0 120000 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_511
timestamp 1679581782
transform 1 0 120672 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_518
timestamp 1679581782
transform 1 0 121344 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_525
timestamp 1679581782
transform 1 0 122016 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_532
timestamp 1679581782
transform 1 0 122688 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_539
timestamp 1679581782
transform 1 0 123360 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_546
timestamp 1679581782
transform 1 0 124032 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_553
timestamp 1679581782
transform 1 0 124704 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_560
timestamp 1679581782
transform 1 0 125376 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_567
timestamp 1679581782
transform 1 0 126048 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_574
timestamp 1679581782
transform 1 0 126720 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_581
timestamp 1679581782
transform 1 0 127392 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_588
timestamp 1679581782
transform 1 0 128064 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_595
timestamp 1679581782
transform 1 0 128736 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_602
timestamp 1679581782
transform 1 0 129408 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_609
timestamp 1679581782
transform 1 0 130080 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_616
timestamp 1679581782
transform 1 0 130752 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_623
timestamp 1679581782
transform 1 0 131424 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_630
timestamp 1679581782
transform 1 0 132096 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_637
timestamp 1679581782
transform 1 0 132768 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_644
timestamp 1679581782
transform 1 0 133440 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_651
timestamp 1679581782
transform 1 0 134112 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_658
timestamp 1679581782
transform 1 0 134784 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_665
timestamp 1679581782
transform 1 0 135456 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_672
timestamp 1679581782
transform 1 0 136128 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_679
timestamp 1679581782
transform 1 0 136800 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_686
timestamp 1679581782
transform 1 0 137472 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_693
timestamp 1679581782
transform 1 0 138144 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_700
timestamp 1679581782
transform 1 0 138816 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_707
timestamp 1679581782
transform 1 0 139488 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_714
timestamp 1679581782
transform 1 0 140160 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_721
timestamp 1679581782
transform 1 0 140832 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_728
timestamp 1679581782
transform 1 0 141504 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_735
timestamp 1679581782
transform 1 0 142176 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_742
timestamp 1679581782
transform 1 0 142848 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_749
timestamp 1679581782
transform 1 0 143520 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_756
timestamp 1679581782
transform 1 0 144192 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_763
timestamp 1679581782
transform 1 0 144864 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_770
timestamp 1679581782
transform 1 0 145536 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_777
timestamp 1679581782
transform 1 0 146208 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_784
timestamp 1679581782
transform 1 0 146880 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_791
timestamp 1679581782
transform 1 0 147552 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_798
timestamp 1679581782
transform 1 0 148224 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_805
timestamp 1679581782
transform 1 0 148896 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_812
timestamp 1679581782
transform 1 0 149568 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_819
timestamp 1679581782
transform 1 0 150240 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_826
timestamp 1679581782
transform 1 0 150912 0 1 126252
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_833
timestamp 1679581782
transform 1 0 151584 0 1 126252
box -48 -56 720 834
use sg13g2_fill_1  FILLER_72_840
timestamp 1677579658
transform 1 0 152256 0 1 126252
box -48 -56 144 834
use sg13g2_decap_8  FILLER_73_0
timestamp 1679581782
transform 1 0 71616 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_7
timestamp 1679581782
transform 1 0 72288 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_14
timestamp 1679581782
transform 1 0 72960 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_21
timestamp 1679581782
transform 1 0 73632 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_28
timestamp 1679581782
transform 1 0 74304 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_35
timestamp 1679581782
transform 1 0 74976 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_42
timestamp 1679581782
transform 1 0 75648 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_49
timestamp 1679581782
transform 1 0 76320 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_56
timestamp 1679581782
transform 1 0 76992 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_63
timestamp 1679581782
transform 1 0 77664 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_70
timestamp 1679581782
transform 1 0 78336 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_77
timestamp 1679581782
transform 1 0 79008 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_84
timestamp 1679581782
transform 1 0 79680 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_91
timestamp 1679581782
transform 1 0 80352 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_98
timestamp 1679581782
transform 1 0 81024 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_105
timestamp 1679581782
transform 1 0 81696 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_112
timestamp 1679581782
transform 1 0 82368 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_119
timestamp 1679581782
transform 1 0 83040 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_126
timestamp 1679581782
transform 1 0 83712 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_133
timestamp 1679581782
transform 1 0 84384 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_140
timestamp 1679581782
transform 1 0 85056 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_147
timestamp 1679581782
transform 1 0 85728 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_154
timestamp 1679581782
transform 1 0 86400 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_161
timestamp 1679581782
transform 1 0 87072 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_168
timestamp 1679581782
transform 1 0 87744 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_175
timestamp 1679581782
transform 1 0 88416 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_182
timestamp 1679581782
transform 1 0 89088 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_189
timestamp 1679581782
transform 1 0 89760 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_196
timestamp 1679581782
transform 1 0 90432 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_203
timestamp 1679581782
transform 1 0 91104 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_210
timestamp 1679581782
transform 1 0 91776 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_217
timestamp 1679581782
transform 1 0 92448 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_224
timestamp 1679581782
transform 1 0 93120 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_231
timestamp 1679581782
transform 1 0 93792 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_238
timestamp 1679581782
transform 1 0 94464 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_245
timestamp 1679581782
transform 1 0 95136 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_252
timestamp 1679581782
transform 1 0 95808 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_259
timestamp 1679581782
transform 1 0 96480 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_266
timestamp 1679581782
transform 1 0 97152 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_273
timestamp 1679581782
transform 1 0 97824 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_280
timestamp 1679581782
transform 1 0 98496 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_287
timestamp 1679581782
transform 1 0 99168 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_294
timestamp 1679581782
transform 1 0 99840 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_301
timestamp 1679581782
transform 1 0 100512 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_308
timestamp 1679581782
transform 1 0 101184 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_315
timestamp 1679581782
transform 1 0 101856 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_322
timestamp 1679581782
transform 1 0 102528 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_329
timestamp 1679581782
transform 1 0 103200 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_336
timestamp 1679581782
transform 1 0 103872 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_343
timestamp 1679581782
transform 1 0 104544 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_350
timestamp 1679581782
transform 1 0 105216 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_357
timestamp 1679581782
transform 1 0 105888 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_364
timestamp 1679581782
transform 1 0 106560 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_371
timestamp 1679581782
transform 1 0 107232 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_378
timestamp 1679581782
transform 1 0 107904 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_385
timestamp 1679581782
transform 1 0 108576 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_392
timestamp 1679581782
transform 1 0 109248 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_399
timestamp 1679581782
transform 1 0 109920 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_406
timestamp 1679581782
transform 1 0 110592 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_413
timestamp 1679581782
transform 1 0 111264 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_420
timestamp 1679581782
transform 1 0 111936 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_427
timestamp 1679581782
transform 1 0 112608 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_434
timestamp 1679581782
transform 1 0 113280 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_441
timestamp 1679581782
transform 1 0 113952 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_448
timestamp 1679581782
transform 1 0 114624 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_455
timestamp 1679581782
transform 1 0 115296 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_462
timestamp 1679581782
transform 1 0 115968 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_469
timestamp 1679581782
transform 1 0 116640 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_476
timestamp 1679581782
transform 1 0 117312 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_483
timestamp 1679581782
transform 1 0 117984 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_490
timestamp 1679581782
transform 1 0 118656 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_497
timestamp 1679581782
transform 1 0 119328 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_504
timestamp 1679581782
transform 1 0 120000 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_511
timestamp 1679581782
transform 1 0 120672 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_518
timestamp 1679581782
transform 1 0 121344 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_525
timestamp 1679581782
transform 1 0 122016 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_532
timestamp 1679581782
transform 1 0 122688 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_539
timestamp 1679581782
transform 1 0 123360 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_546
timestamp 1679581782
transform 1 0 124032 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_553
timestamp 1679581782
transform 1 0 124704 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_560
timestamp 1679581782
transform 1 0 125376 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_567
timestamp 1679581782
transform 1 0 126048 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_574
timestamp 1679581782
transform 1 0 126720 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_581
timestamp 1679581782
transform 1 0 127392 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_588
timestamp 1679581782
transform 1 0 128064 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_595
timestamp 1679581782
transform 1 0 128736 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_602
timestamp 1679581782
transform 1 0 129408 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_609
timestamp 1679581782
transform 1 0 130080 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_616
timestamp 1679581782
transform 1 0 130752 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_623
timestamp 1679581782
transform 1 0 131424 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_630
timestamp 1679581782
transform 1 0 132096 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_637
timestamp 1679581782
transform 1 0 132768 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_644
timestamp 1679581782
transform 1 0 133440 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_651
timestamp 1679581782
transform 1 0 134112 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_658
timestamp 1679581782
transform 1 0 134784 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_665
timestamp 1679581782
transform 1 0 135456 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_672
timestamp 1679581782
transform 1 0 136128 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_679
timestamp 1679581782
transform 1 0 136800 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_686
timestamp 1679581782
transform 1 0 137472 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_693
timestamp 1679581782
transform 1 0 138144 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_700
timestamp 1679581782
transform 1 0 138816 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_707
timestamp 1679581782
transform 1 0 139488 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_714
timestamp 1679581782
transform 1 0 140160 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_721
timestamp 1679581782
transform 1 0 140832 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_728
timestamp 1679581782
transform 1 0 141504 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_735
timestamp 1679581782
transform 1 0 142176 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_742
timestamp 1679581782
transform 1 0 142848 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_749
timestamp 1679581782
transform 1 0 143520 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_756
timestamp 1679581782
transform 1 0 144192 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_763
timestamp 1679581782
transform 1 0 144864 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_770
timestamp 1679581782
transform 1 0 145536 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_777
timestamp 1679581782
transform 1 0 146208 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_784
timestamp 1679581782
transform 1 0 146880 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_791
timestamp 1679581782
transform 1 0 147552 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_798
timestamp 1679581782
transform 1 0 148224 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_805
timestamp 1679581782
transform 1 0 148896 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_812
timestamp 1679581782
transform 1 0 149568 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_819
timestamp 1679581782
transform 1 0 150240 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_826
timestamp 1679581782
transform 1 0 150912 0 -1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_833
timestamp 1679581782
transform 1 0 151584 0 -1 127764
box -48 -56 720 834
use sg13g2_fill_1  FILLER_73_840
timestamp 1677579658
transform 1 0 152256 0 -1 127764
box -48 -56 144 834
use sg13g2_decap_8  FILLER_74_0
timestamp 1679581782
transform 1 0 71616 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_7
timestamp 1679581782
transform 1 0 72288 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_14
timestamp 1679581782
transform 1 0 72960 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_21
timestamp 1679581782
transform 1 0 73632 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_28
timestamp 1679581782
transform 1 0 74304 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_35
timestamp 1679581782
transform 1 0 74976 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_42
timestamp 1679581782
transform 1 0 75648 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_49
timestamp 1679581782
transform 1 0 76320 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_56
timestamp 1679581782
transform 1 0 76992 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_63
timestamp 1679581782
transform 1 0 77664 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_70
timestamp 1679581782
transform 1 0 78336 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_77
timestamp 1679581782
transform 1 0 79008 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_84
timestamp 1679581782
transform 1 0 79680 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_91
timestamp 1679581782
transform 1 0 80352 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_98
timestamp 1679581782
transform 1 0 81024 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_105
timestamp 1679581782
transform 1 0 81696 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_112
timestamp 1679581782
transform 1 0 82368 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_119
timestamp 1679581782
transform 1 0 83040 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_126
timestamp 1679581782
transform 1 0 83712 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_133
timestamp 1679581782
transform 1 0 84384 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_140
timestamp 1679581782
transform 1 0 85056 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_147
timestamp 1679581782
transform 1 0 85728 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_154
timestamp 1679581782
transform 1 0 86400 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_161
timestamp 1679581782
transform 1 0 87072 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_168
timestamp 1679581782
transform 1 0 87744 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_175
timestamp 1679581782
transform 1 0 88416 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_182
timestamp 1679581782
transform 1 0 89088 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_189
timestamp 1679581782
transform 1 0 89760 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_196
timestamp 1679581782
transform 1 0 90432 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_203
timestamp 1679581782
transform 1 0 91104 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_210
timestamp 1679581782
transform 1 0 91776 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_217
timestamp 1679581782
transform 1 0 92448 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_224
timestamp 1679581782
transform 1 0 93120 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_231
timestamp 1679581782
transform 1 0 93792 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_238
timestamp 1679581782
transform 1 0 94464 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_245
timestamp 1679581782
transform 1 0 95136 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_252
timestamp 1679581782
transform 1 0 95808 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_259
timestamp 1679581782
transform 1 0 96480 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_266
timestamp 1679581782
transform 1 0 97152 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_273
timestamp 1679581782
transform 1 0 97824 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_280
timestamp 1679581782
transform 1 0 98496 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_287
timestamp 1679581782
transform 1 0 99168 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_294
timestamp 1679581782
transform 1 0 99840 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_301
timestamp 1679581782
transform 1 0 100512 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_308
timestamp 1679581782
transform 1 0 101184 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_315
timestamp 1679581782
transform 1 0 101856 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_322
timestamp 1679581782
transform 1 0 102528 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_329
timestamp 1679581782
transform 1 0 103200 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_336
timestamp 1679581782
transform 1 0 103872 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_343
timestamp 1679581782
transform 1 0 104544 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_350
timestamp 1679581782
transform 1 0 105216 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_357
timestamp 1679581782
transform 1 0 105888 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_364
timestamp 1679581782
transform 1 0 106560 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_371
timestamp 1679581782
transform 1 0 107232 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_378
timestamp 1679581782
transform 1 0 107904 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_385
timestamp 1679581782
transform 1 0 108576 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_392
timestamp 1679581782
transform 1 0 109248 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_399
timestamp 1679581782
transform 1 0 109920 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_406
timestamp 1679581782
transform 1 0 110592 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_413
timestamp 1679581782
transform 1 0 111264 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_420
timestamp 1679581782
transform 1 0 111936 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_427
timestamp 1679581782
transform 1 0 112608 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_434
timestamp 1679581782
transform 1 0 113280 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_441
timestamp 1679581782
transform 1 0 113952 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_448
timestamp 1679581782
transform 1 0 114624 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_455
timestamp 1679581782
transform 1 0 115296 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_462
timestamp 1679581782
transform 1 0 115968 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_469
timestamp 1679581782
transform 1 0 116640 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_476
timestamp 1679581782
transform 1 0 117312 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_483
timestamp 1679581782
transform 1 0 117984 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_490
timestamp 1679581782
transform 1 0 118656 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_497
timestamp 1679581782
transform 1 0 119328 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_504
timestamp 1679581782
transform 1 0 120000 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_511
timestamp 1679581782
transform 1 0 120672 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_518
timestamp 1679581782
transform 1 0 121344 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_525
timestamp 1679581782
transform 1 0 122016 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_532
timestamp 1679581782
transform 1 0 122688 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_539
timestamp 1679581782
transform 1 0 123360 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_546
timestamp 1679581782
transform 1 0 124032 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_553
timestamp 1679581782
transform 1 0 124704 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_560
timestamp 1679581782
transform 1 0 125376 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_567
timestamp 1679581782
transform 1 0 126048 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_574
timestamp 1679581782
transform 1 0 126720 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_581
timestamp 1679581782
transform 1 0 127392 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_588
timestamp 1679581782
transform 1 0 128064 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_595
timestamp 1679581782
transform 1 0 128736 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_602
timestamp 1679581782
transform 1 0 129408 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_609
timestamp 1679581782
transform 1 0 130080 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_616
timestamp 1679581782
transform 1 0 130752 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_623
timestamp 1679581782
transform 1 0 131424 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_630
timestamp 1679581782
transform 1 0 132096 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_637
timestamp 1679581782
transform 1 0 132768 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_644
timestamp 1679581782
transform 1 0 133440 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_651
timestamp 1679581782
transform 1 0 134112 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_658
timestamp 1679581782
transform 1 0 134784 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_665
timestamp 1679581782
transform 1 0 135456 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_672
timestamp 1679581782
transform 1 0 136128 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_679
timestamp 1679581782
transform 1 0 136800 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_686
timestamp 1679581782
transform 1 0 137472 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_693
timestamp 1679581782
transform 1 0 138144 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_700
timestamp 1679581782
transform 1 0 138816 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_707
timestamp 1679581782
transform 1 0 139488 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_714
timestamp 1679581782
transform 1 0 140160 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_721
timestamp 1679581782
transform 1 0 140832 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_728
timestamp 1679581782
transform 1 0 141504 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_735
timestamp 1679581782
transform 1 0 142176 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_742
timestamp 1679581782
transform 1 0 142848 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_749
timestamp 1679581782
transform 1 0 143520 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_756
timestamp 1679581782
transform 1 0 144192 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_763
timestamp 1679581782
transform 1 0 144864 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_770
timestamp 1679581782
transform 1 0 145536 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_777
timestamp 1679581782
transform 1 0 146208 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_784
timestamp 1679581782
transform 1 0 146880 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_791
timestamp 1679581782
transform 1 0 147552 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_798
timestamp 1679581782
transform 1 0 148224 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_805
timestamp 1679581782
transform 1 0 148896 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_812
timestamp 1679581782
transform 1 0 149568 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_819
timestamp 1679581782
transform 1 0 150240 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_826
timestamp 1679581782
transform 1 0 150912 0 1 127764
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_833
timestamp 1679581782
transform 1 0 151584 0 1 127764
box -48 -56 720 834
use sg13g2_fill_1  FILLER_74_840
timestamp 1677579658
transform 1 0 152256 0 1 127764
box -48 -56 144 834
use sg13g2_decap_8  FILLER_75_0
timestamp 1679581782
transform 1 0 71616 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_7
timestamp 1679581782
transform 1 0 72288 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_14
timestamp 1679581782
transform 1 0 72960 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_21
timestamp 1679581782
transform 1 0 73632 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_28
timestamp 1679581782
transform 1 0 74304 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_35
timestamp 1679581782
transform 1 0 74976 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_42
timestamp 1679581782
transform 1 0 75648 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_49
timestamp 1679581782
transform 1 0 76320 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_56
timestamp 1679581782
transform 1 0 76992 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_63
timestamp 1679581782
transform 1 0 77664 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_70
timestamp 1679581782
transform 1 0 78336 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_77
timestamp 1679581782
transform 1 0 79008 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_84
timestamp 1679581782
transform 1 0 79680 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_91
timestamp 1679581782
transform 1 0 80352 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_98
timestamp 1679581782
transform 1 0 81024 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_105
timestamp 1679581782
transform 1 0 81696 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_112
timestamp 1679581782
transform 1 0 82368 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_119
timestamp 1679581782
transform 1 0 83040 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_126
timestamp 1679581782
transform 1 0 83712 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_133
timestamp 1679581782
transform 1 0 84384 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_140
timestamp 1679581782
transform 1 0 85056 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_147
timestamp 1679581782
transform 1 0 85728 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_154
timestamp 1679581782
transform 1 0 86400 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_161
timestamp 1679581782
transform 1 0 87072 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_168
timestamp 1679581782
transform 1 0 87744 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_175
timestamp 1679581782
transform 1 0 88416 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_182
timestamp 1679581782
transform 1 0 89088 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_189
timestamp 1679581782
transform 1 0 89760 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_196
timestamp 1679581782
transform 1 0 90432 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_203
timestamp 1679581782
transform 1 0 91104 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_210
timestamp 1679581782
transform 1 0 91776 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_217
timestamp 1679581782
transform 1 0 92448 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_224
timestamp 1679581782
transform 1 0 93120 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_231
timestamp 1679581782
transform 1 0 93792 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_238
timestamp 1679581782
transform 1 0 94464 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_245
timestamp 1679581782
transform 1 0 95136 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_252
timestamp 1679581782
transform 1 0 95808 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_259
timestamp 1679581782
transform 1 0 96480 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_266
timestamp 1679581782
transform 1 0 97152 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_273
timestamp 1679581782
transform 1 0 97824 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_280
timestamp 1679581782
transform 1 0 98496 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_287
timestamp 1679581782
transform 1 0 99168 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_294
timestamp 1679581782
transform 1 0 99840 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_301
timestamp 1679581782
transform 1 0 100512 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_308
timestamp 1679581782
transform 1 0 101184 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_315
timestamp 1679581782
transform 1 0 101856 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_322
timestamp 1679581782
transform 1 0 102528 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_329
timestamp 1679581782
transform 1 0 103200 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_336
timestamp 1679581782
transform 1 0 103872 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_343
timestamp 1679581782
transform 1 0 104544 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_350
timestamp 1679581782
transform 1 0 105216 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_357
timestamp 1679581782
transform 1 0 105888 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_364
timestamp 1679581782
transform 1 0 106560 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_371
timestamp 1679581782
transform 1 0 107232 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_378
timestamp 1679581782
transform 1 0 107904 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_385
timestamp 1679581782
transform 1 0 108576 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_392
timestamp 1679581782
transform 1 0 109248 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_399
timestamp 1679581782
transform 1 0 109920 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_406
timestamp 1679581782
transform 1 0 110592 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_413
timestamp 1679581782
transform 1 0 111264 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_420
timestamp 1679581782
transform 1 0 111936 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_427
timestamp 1679581782
transform 1 0 112608 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_434
timestamp 1679581782
transform 1 0 113280 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_441
timestamp 1679581782
transform 1 0 113952 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_448
timestamp 1679581782
transform 1 0 114624 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_455
timestamp 1679581782
transform 1 0 115296 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_462
timestamp 1679581782
transform 1 0 115968 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_469
timestamp 1679581782
transform 1 0 116640 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_476
timestamp 1679581782
transform 1 0 117312 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_483
timestamp 1679581782
transform 1 0 117984 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_490
timestamp 1679581782
transform 1 0 118656 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_497
timestamp 1679581782
transform 1 0 119328 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_504
timestamp 1679581782
transform 1 0 120000 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_511
timestamp 1679581782
transform 1 0 120672 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_518
timestamp 1679581782
transform 1 0 121344 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_525
timestamp 1679581782
transform 1 0 122016 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_532
timestamp 1679581782
transform 1 0 122688 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_539
timestamp 1679581782
transform 1 0 123360 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_546
timestamp 1679581782
transform 1 0 124032 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_553
timestamp 1679581782
transform 1 0 124704 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_560
timestamp 1679581782
transform 1 0 125376 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_567
timestamp 1679581782
transform 1 0 126048 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_574
timestamp 1679581782
transform 1 0 126720 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_581
timestamp 1679581782
transform 1 0 127392 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_588
timestamp 1679581782
transform 1 0 128064 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_595
timestamp 1679581782
transform 1 0 128736 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_602
timestamp 1679581782
transform 1 0 129408 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_609
timestamp 1679581782
transform 1 0 130080 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_616
timestamp 1679581782
transform 1 0 130752 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_623
timestamp 1679581782
transform 1 0 131424 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_630
timestamp 1679581782
transform 1 0 132096 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_637
timestamp 1679581782
transform 1 0 132768 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_644
timestamp 1679581782
transform 1 0 133440 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_651
timestamp 1679581782
transform 1 0 134112 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_658
timestamp 1679581782
transform 1 0 134784 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_665
timestamp 1679581782
transform 1 0 135456 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_672
timestamp 1679581782
transform 1 0 136128 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_679
timestamp 1679581782
transform 1 0 136800 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_686
timestamp 1679581782
transform 1 0 137472 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_693
timestamp 1679581782
transform 1 0 138144 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_700
timestamp 1679581782
transform 1 0 138816 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_707
timestamp 1679581782
transform 1 0 139488 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_714
timestamp 1679581782
transform 1 0 140160 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_721
timestamp 1679581782
transform 1 0 140832 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_728
timestamp 1679581782
transform 1 0 141504 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_735
timestamp 1679581782
transform 1 0 142176 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_742
timestamp 1679581782
transform 1 0 142848 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_749
timestamp 1679581782
transform 1 0 143520 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_756
timestamp 1679581782
transform 1 0 144192 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_763
timestamp 1679581782
transform 1 0 144864 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_770
timestamp 1679581782
transform 1 0 145536 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_777
timestamp 1679581782
transform 1 0 146208 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_784
timestamp 1679581782
transform 1 0 146880 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_791
timestamp 1679581782
transform 1 0 147552 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_798
timestamp 1679581782
transform 1 0 148224 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_805
timestamp 1679581782
transform 1 0 148896 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_812
timestamp 1679581782
transform 1 0 149568 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_819
timestamp 1679581782
transform 1 0 150240 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_826
timestamp 1679581782
transform 1 0 150912 0 -1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_833
timestamp 1679581782
transform 1 0 151584 0 -1 129276
box -48 -56 720 834
use sg13g2_fill_1  FILLER_75_840
timestamp 1677579658
transform 1 0 152256 0 -1 129276
box -48 -56 144 834
use sg13g2_decap_8  FILLER_76_0
timestamp 1679581782
transform 1 0 71616 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_7
timestamp 1679581782
transform 1 0 72288 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_14
timestamp 1679581782
transform 1 0 72960 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_21
timestamp 1679581782
transform 1 0 73632 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_28
timestamp 1679581782
transform 1 0 74304 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_35
timestamp 1679581782
transform 1 0 74976 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_42
timestamp 1679581782
transform 1 0 75648 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_49
timestamp 1679581782
transform 1 0 76320 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_56
timestamp 1679581782
transform 1 0 76992 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_63
timestamp 1679581782
transform 1 0 77664 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_70
timestamp 1679581782
transform 1 0 78336 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_77
timestamp 1679581782
transform 1 0 79008 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_84
timestamp 1679581782
transform 1 0 79680 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_91
timestamp 1679581782
transform 1 0 80352 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_98
timestamp 1679581782
transform 1 0 81024 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_105
timestamp 1679581782
transform 1 0 81696 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_112
timestamp 1679581782
transform 1 0 82368 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_119
timestamp 1679581782
transform 1 0 83040 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_126
timestamp 1679581782
transform 1 0 83712 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_133
timestamp 1679581782
transform 1 0 84384 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_140
timestamp 1679581782
transform 1 0 85056 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_147
timestamp 1679581782
transform 1 0 85728 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_154
timestamp 1679581782
transform 1 0 86400 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_161
timestamp 1679581782
transform 1 0 87072 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_168
timestamp 1679581782
transform 1 0 87744 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_175
timestamp 1679581782
transform 1 0 88416 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_182
timestamp 1679581782
transform 1 0 89088 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_189
timestamp 1679581782
transform 1 0 89760 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_196
timestamp 1679581782
transform 1 0 90432 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_203
timestamp 1679581782
transform 1 0 91104 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_210
timestamp 1679581782
transform 1 0 91776 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_217
timestamp 1679581782
transform 1 0 92448 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_224
timestamp 1679581782
transform 1 0 93120 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_231
timestamp 1679581782
transform 1 0 93792 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_238
timestamp 1679581782
transform 1 0 94464 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_245
timestamp 1679581782
transform 1 0 95136 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_252
timestamp 1679581782
transform 1 0 95808 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_259
timestamp 1679581782
transform 1 0 96480 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_266
timestamp 1679581782
transform 1 0 97152 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_273
timestamp 1679581782
transform 1 0 97824 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_280
timestamp 1679581782
transform 1 0 98496 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_287
timestamp 1679581782
transform 1 0 99168 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_294
timestamp 1679581782
transform 1 0 99840 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_301
timestamp 1679581782
transform 1 0 100512 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_308
timestamp 1679581782
transform 1 0 101184 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_315
timestamp 1679581782
transform 1 0 101856 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_322
timestamp 1679581782
transform 1 0 102528 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_329
timestamp 1679581782
transform 1 0 103200 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_336
timestamp 1679581782
transform 1 0 103872 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_343
timestamp 1679581782
transform 1 0 104544 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_350
timestamp 1679581782
transform 1 0 105216 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_357
timestamp 1679581782
transform 1 0 105888 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_364
timestamp 1679581782
transform 1 0 106560 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_371
timestamp 1679581782
transform 1 0 107232 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_378
timestamp 1679581782
transform 1 0 107904 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_385
timestamp 1679581782
transform 1 0 108576 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_392
timestamp 1679581782
transform 1 0 109248 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_399
timestamp 1679581782
transform 1 0 109920 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_406
timestamp 1679581782
transform 1 0 110592 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_413
timestamp 1679581782
transform 1 0 111264 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_420
timestamp 1679581782
transform 1 0 111936 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_427
timestamp 1679581782
transform 1 0 112608 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_434
timestamp 1679581782
transform 1 0 113280 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_441
timestamp 1679581782
transform 1 0 113952 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_448
timestamp 1679581782
transform 1 0 114624 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_455
timestamp 1679581782
transform 1 0 115296 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_462
timestamp 1679581782
transform 1 0 115968 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_469
timestamp 1679581782
transform 1 0 116640 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_476
timestamp 1679581782
transform 1 0 117312 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_483
timestamp 1679581782
transform 1 0 117984 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_490
timestamp 1679581782
transform 1 0 118656 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_497
timestamp 1679581782
transform 1 0 119328 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_504
timestamp 1679581782
transform 1 0 120000 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_511
timestamp 1679581782
transform 1 0 120672 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_518
timestamp 1679581782
transform 1 0 121344 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_525
timestamp 1679581782
transform 1 0 122016 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_532
timestamp 1679581782
transform 1 0 122688 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_539
timestamp 1679581782
transform 1 0 123360 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_546
timestamp 1679581782
transform 1 0 124032 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_553
timestamp 1679581782
transform 1 0 124704 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_560
timestamp 1679581782
transform 1 0 125376 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_567
timestamp 1679581782
transform 1 0 126048 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_574
timestamp 1679581782
transform 1 0 126720 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_581
timestamp 1679581782
transform 1 0 127392 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_588
timestamp 1679581782
transform 1 0 128064 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_595
timestamp 1679581782
transform 1 0 128736 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_602
timestamp 1679581782
transform 1 0 129408 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_609
timestamp 1679581782
transform 1 0 130080 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_616
timestamp 1679581782
transform 1 0 130752 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_623
timestamp 1679581782
transform 1 0 131424 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_630
timestamp 1679581782
transform 1 0 132096 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_637
timestamp 1679581782
transform 1 0 132768 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_644
timestamp 1679581782
transform 1 0 133440 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_651
timestamp 1679581782
transform 1 0 134112 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_658
timestamp 1679581782
transform 1 0 134784 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_665
timestamp 1679581782
transform 1 0 135456 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_672
timestamp 1679581782
transform 1 0 136128 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_679
timestamp 1679581782
transform 1 0 136800 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_686
timestamp 1679581782
transform 1 0 137472 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_693
timestamp 1679581782
transform 1 0 138144 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_700
timestamp 1679581782
transform 1 0 138816 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_707
timestamp 1679581782
transform 1 0 139488 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_714
timestamp 1679581782
transform 1 0 140160 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_721
timestamp 1679581782
transform 1 0 140832 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_728
timestamp 1679581782
transform 1 0 141504 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_735
timestamp 1679581782
transform 1 0 142176 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_742
timestamp 1679581782
transform 1 0 142848 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_749
timestamp 1679581782
transform 1 0 143520 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_756
timestamp 1679581782
transform 1 0 144192 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_763
timestamp 1679581782
transform 1 0 144864 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_770
timestamp 1679581782
transform 1 0 145536 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_777
timestamp 1679581782
transform 1 0 146208 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_784
timestamp 1679581782
transform 1 0 146880 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_791
timestamp 1679581782
transform 1 0 147552 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_798
timestamp 1679581782
transform 1 0 148224 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_805
timestamp 1679581782
transform 1 0 148896 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_812
timestamp 1679581782
transform 1 0 149568 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_819
timestamp 1679581782
transform 1 0 150240 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_826
timestamp 1679581782
transform 1 0 150912 0 1 129276
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_833
timestamp 1679581782
transform 1 0 151584 0 1 129276
box -48 -56 720 834
use sg13g2_fill_1  FILLER_76_840
timestamp 1677579658
transform 1 0 152256 0 1 129276
box -48 -56 144 834
use sg13g2_decap_8  FILLER_77_0
timestamp 1679581782
transform 1 0 71616 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_7
timestamp 1679581782
transform 1 0 72288 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_14
timestamp 1679581782
transform 1 0 72960 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_21
timestamp 1679581782
transform 1 0 73632 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_28
timestamp 1679581782
transform 1 0 74304 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_35
timestamp 1679581782
transform 1 0 74976 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_42
timestamp 1679581782
transform 1 0 75648 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_49
timestamp 1679581782
transform 1 0 76320 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_56
timestamp 1679581782
transform 1 0 76992 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_63
timestamp 1679581782
transform 1 0 77664 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_70
timestamp 1679581782
transform 1 0 78336 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_77
timestamp 1679581782
transform 1 0 79008 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_84
timestamp 1679581782
transform 1 0 79680 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_91
timestamp 1679581782
transform 1 0 80352 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_98
timestamp 1679581782
transform 1 0 81024 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_105
timestamp 1679581782
transform 1 0 81696 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_112
timestamp 1679581782
transform 1 0 82368 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_119
timestamp 1679581782
transform 1 0 83040 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_126
timestamp 1679581782
transform 1 0 83712 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_133
timestamp 1679581782
transform 1 0 84384 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_140
timestamp 1679581782
transform 1 0 85056 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_147
timestamp 1679581782
transform 1 0 85728 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_154
timestamp 1679581782
transform 1 0 86400 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_161
timestamp 1679581782
transform 1 0 87072 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_168
timestamp 1679581782
transform 1 0 87744 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_175
timestamp 1679581782
transform 1 0 88416 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_182
timestamp 1679581782
transform 1 0 89088 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_189
timestamp 1679581782
transform 1 0 89760 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_196
timestamp 1679581782
transform 1 0 90432 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_203
timestamp 1679581782
transform 1 0 91104 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_210
timestamp 1679581782
transform 1 0 91776 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_217
timestamp 1679581782
transform 1 0 92448 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_224
timestamp 1679581782
transform 1 0 93120 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_231
timestamp 1679581782
transform 1 0 93792 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_238
timestamp 1679581782
transform 1 0 94464 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_245
timestamp 1679581782
transform 1 0 95136 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_252
timestamp 1679581782
transform 1 0 95808 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_259
timestamp 1679581782
transform 1 0 96480 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_266
timestamp 1679581782
transform 1 0 97152 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_273
timestamp 1679581782
transform 1 0 97824 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_280
timestamp 1679581782
transform 1 0 98496 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_287
timestamp 1679581782
transform 1 0 99168 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_294
timestamp 1679581782
transform 1 0 99840 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_301
timestamp 1679581782
transform 1 0 100512 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_308
timestamp 1679581782
transform 1 0 101184 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_315
timestamp 1679581782
transform 1 0 101856 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_322
timestamp 1679581782
transform 1 0 102528 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_329
timestamp 1679581782
transform 1 0 103200 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_336
timestamp 1679581782
transform 1 0 103872 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_343
timestamp 1679581782
transform 1 0 104544 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_350
timestamp 1679581782
transform 1 0 105216 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_357
timestamp 1679581782
transform 1 0 105888 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_364
timestamp 1679581782
transform 1 0 106560 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_371
timestamp 1679581782
transform 1 0 107232 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_378
timestamp 1679581782
transform 1 0 107904 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_385
timestamp 1679581782
transform 1 0 108576 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_392
timestamp 1679581782
transform 1 0 109248 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_399
timestamp 1679581782
transform 1 0 109920 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_406
timestamp 1679581782
transform 1 0 110592 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_413
timestamp 1679581782
transform 1 0 111264 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_420
timestamp 1679581782
transform 1 0 111936 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_427
timestamp 1679581782
transform 1 0 112608 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_434
timestamp 1679581782
transform 1 0 113280 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_441
timestamp 1679581782
transform 1 0 113952 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_448
timestamp 1679581782
transform 1 0 114624 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_455
timestamp 1679581782
transform 1 0 115296 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_462
timestamp 1679581782
transform 1 0 115968 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_469
timestamp 1679581782
transform 1 0 116640 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_476
timestamp 1679581782
transform 1 0 117312 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_483
timestamp 1679581782
transform 1 0 117984 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_490
timestamp 1679581782
transform 1 0 118656 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_497
timestamp 1679581782
transform 1 0 119328 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_504
timestamp 1679581782
transform 1 0 120000 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_511
timestamp 1679581782
transform 1 0 120672 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_518
timestamp 1679581782
transform 1 0 121344 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_525
timestamp 1679581782
transform 1 0 122016 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_532
timestamp 1679581782
transform 1 0 122688 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_539
timestamp 1679581782
transform 1 0 123360 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_546
timestamp 1679581782
transform 1 0 124032 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_553
timestamp 1679581782
transform 1 0 124704 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_560
timestamp 1679581782
transform 1 0 125376 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_567
timestamp 1679581782
transform 1 0 126048 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_574
timestamp 1679581782
transform 1 0 126720 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_581
timestamp 1679581782
transform 1 0 127392 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_588
timestamp 1679581782
transform 1 0 128064 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_595
timestamp 1679581782
transform 1 0 128736 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_602
timestamp 1679581782
transform 1 0 129408 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_609
timestamp 1679581782
transform 1 0 130080 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_616
timestamp 1679581782
transform 1 0 130752 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_623
timestamp 1679581782
transform 1 0 131424 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_630
timestamp 1679581782
transform 1 0 132096 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_637
timestamp 1679581782
transform 1 0 132768 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_644
timestamp 1679581782
transform 1 0 133440 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_651
timestamp 1679581782
transform 1 0 134112 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_658
timestamp 1679581782
transform 1 0 134784 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_665
timestamp 1679581782
transform 1 0 135456 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_672
timestamp 1679581782
transform 1 0 136128 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_679
timestamp 1679581782
transform 1 0 136800 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_686
timestamp 1679581782
transform 1 0 137472 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_693
timestamp 1679581782
transform 1 0 138144 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_700
timestamp 1679581782
transform 1 0 138816 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_707
timestamp 1679581782
transform 1 0 139488 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_714
timestamp 1679581782
transform 1 0 140160 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_721
timestamp 1679581782
transform 1 0 140832 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_728
timestamp 1679581782
transform 1 0 141504 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_735
timestamp 1679581782
transform 1 0 142176 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_742
timestamp 1679581782
transform 1 0 142848 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_749
timestamp 1679581782
transform 1 0 143520 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_756
timestamp 1679581782
transform 1 0 144192 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_763
timestamp 1679581782
transform 1 0 144864 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_770
timestamp 1679581782
transform 1 0 145536 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_777
timestamp 1679581782
transform 1 0 146208 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_784
timestamp 1679581782
transform 1 0 146880 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_791
timestamp 1679581782
transform 1 0 147552 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_798
timestamp 1679581782
transform 1 0 148224 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_805
timestamp 1679581782
transform 1 0 148896 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_812
timestamp 1679581782
transform 1 0 149568 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_819
timestamp 1679581782
transform 1 0 150240 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_826
timestamp 1679581782
transform 1 0 150912 0 -1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_833
timestamp 1679581782
transform 1 0 151584 0 -1 130788
box -48 -56 720 834
use sg13g2_fill_1  FILLER_77_840
timestamp 1677579658
transform 1 0 152256 0 -1 130788
box -48 -56 144 834
use sg13g2_decap_8  FILLER_78_0
timestamp 1679581782
transform 1 0 71616 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_7
timestamp 1679581782
transform 1 0 72288 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_14
timestamp 1679581782
transform 1 0 72960 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_21
timestamp 1679581782
transform 1 0 73632 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_28
timestamp 1679581782
transform 1 0 74304 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_35
timestamp 1679581782
transform 1 0 74976 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_42
timestamp 1679581782
transform 1 0 75648 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_49
timestamp 1679581782
transform 1 0 76320 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_56
timestamp 1679581782
transform 1 0 76992 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_63
timestamp 1679581782
transform 1 0 77664 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_70
timestamp 1679581782
transform 1 0 78336 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_77
timestamp 1679581782
transform 1 0 79008 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_84
timestamp 1679581782
transform 1 0 79680 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_91
timestamp 1679581782
transform 1 0 80352 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_98
timestamp 1679581782
transform 1 0 81024 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_105
timestamp 1679581782
transform 1 0 81696 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_112
timestamp 1679581782
transform 1 0 82368 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_119
timestamp 1679581782
transform 1 0 83040 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_126
timestamp 1679581782
transform 1 0 83712 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_133
timestamp 1679581782
transform 1 0 84384 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_140
timestamp 1679581782
transform 1 0 85056 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_147
timestamp 1679581782
transform 1 0 85728 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_154
timestamp 1679581782
transform 1 0 86400 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_161
timestamp 1679581782
transform 1 0 87072 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_168
timestamp 1679581782
transform 1 0 87744 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_175
timestamp 1679581782
transform 1 0 88416 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_182
timestamp 1679581782
transform 1 0 89088 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_189
timestamp 1679581782
transform 1 0 89760 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_196
timestamp 1679581782
transform 1 0 90432 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_203
timestamp 1679581782
transform 1 0 91104 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_210
timestamp 1679581782
transform 1 0 91776 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_217
timestamp 1679581782
transform 1 0 92448 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_224
timestamp 1679581782
transform 1 0 93120 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_231
timestamp 1679581782
transform 1 0 93792 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_238
timestamp 1679581782
transform 1 0 94464 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_245
timestamp 1679581782
transform 1 0 95136 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_252
timestamp 1679581782
transform 1 0 95808 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_259
timestamp 1679581782
transform 1 0 96480 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_266
timestamp 1679581782
transform 1 0 97152 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_273
timestamp 1679581782
transform 1 0 97824 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_280
timestamp 1679581782
transform 1 0 98496 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_287
timestamp 1679581782
transform 1 0 99168 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_294
timestamp 1679581782
transform 1 0 99840 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_301
timestamp 1679581782
transform 1 0 100512 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_308
timestamp 1679581782
transform 1 0 101184 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_315
timestamp 1679581782
transform 1 0 101856 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_322
timestamp 1679581782
transform 1 0 102528 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_329
timestamp 1679581782
transform 1 0 103200 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_336
timestamp 1679581782
transform 1 0 103872 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_343
timestamp 1679581782
transform 1 0 104544 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_350
timestamp 1679581782
transform 1 0 105216 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_357
timestamp 1679581782
transform 1 0 105888 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_364
timestamp 1679581782
transform 1 0 106560 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_371
timestamp 1679581782
transform 1 0 107232 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_378
timestamp 1679581782
transform 1 0 107904 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_385
timestamp 1679581782
transform 1 0 108576 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_392
timestamp 1679581782
transform 1 0 109248 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_399
timestamp 1679581782
transform 1 0 109920 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_406
timestamp 1679581782
transform 1 0 110592 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_413
timestamp 1679581782
transform 1 0 111264 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_420
timestamp 1679581782
transform 1 0 111936 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_427
timestamp 1679581782
transform 1 0 112608 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_434
timestamp 1679581782
transform 1 0 113280 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_441
timestamp 1679581782
transform 1 0 113952 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_448
timestamp 1679581782
transform 1 0 114624 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_455
timestamp 1679581782
transform 1 0 115296 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_462
timestamp 1679581782
transform 1 0 115968 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_469
timestamp 1679581782
transform 1 0 116640 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_476
timestamp 1679581782
transform 1 0 117312 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_483
timestamp 1679581782
transform 1 0 117984 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_490
timestamp 1679581782
transform 1 0 118656 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_497
timestamp 1679581782
transform 1 0 119328 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_504
timestamp 1679581782
transform 1 0 120000 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_511
timestamp 1679581782
transform 1 0 120672 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_518
timestamp 1679581782
transform 1 0 121344 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_525
timestamp 1679581782
transform 1 0 122016 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_532
timestamp 1679581782
transform 1 0 122688 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_539
timestamp 1679581782
transform 1 0 123360 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_546
timestamp 1679581782
transform 1 0 124032 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_553
timestamp 1679581782
transform 1 0 124704 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_560
timestamp 1679581782
transform 1 0 125376 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_567
timestamp 1679581782
transform 1 0 126048 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_574
timestamp 1679581782
transform 1 0 126720 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_581
timestamp 1679581782
transform 1 0 127392 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_588
timestamp 1679581782
transform 1 0 128064 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_595
timestamp 1679581782
transform 1 0 128736 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_602
timestamp 1679581782
transform 1 0 129408 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_609
timestamp 1679581782
transform 1 0 130080 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_616
timestamp 1679581782
transform 1 0 130752 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_623
timestamp 1679581782
transform 1 0 131424 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_630
timestamp 1679581782
transform 1 0 132096 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_637
timestamp 1679581782
transform 1 0 132768 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_644
timestamp 1679581782
transform 1 0 133440 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_651
timestamp 1679581782
transform 1 0 134112 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_658
timestamp 1679581782
transform 1 0 134784 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_665
timestamp 1679581782
transform 1 0 135456 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_672
timestamp 1679581782
transform 1 0 136128 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_679
timestamp 1679581782
transform 1 0 136800 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_686
timestamp 1679581782
transform 1 0 137472 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_693
timestamp 1679581782
transform 1 0 138144 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_700
timestamp 1679581782
transform 1 0 138816 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_707
timestamp 1679581782
transform 1 0 139488 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_714
timestamp 1679581782
transform 1 0 140160 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_721
timestamp 1679581782
transform 1 0 140832 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_728
timestamp 1679581782
transform 1 0 141504 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_735
timestamp 1679581782
transform 1 0 142176 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_742
timestamp 1679581782
transform 1 0 142848 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_749
timestamp 1679581782
transform 1 0 143520 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_756
timestamp 1679581782
transform 1 0 144192 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_763
timestamp 1679581782
transform 1 0 144864 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_770
timestamp 1679581782
transform 1 0 145536 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_777
timestamp 1679581782
transform 1 0 146208 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_784
timestamp 1679581782
transform 1 0 146880 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_791
timestamp 1679581782
transform 1 0 147552 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_798
timestamp 1679581782
transform 1 0 148224 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_805
timestamp 1679581782
transform 1 0 148896 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_812
timestamp 1679581782
transform 1 0 149568 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_819
timestamp 1679581782
transform 1 0 150240 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_826
timestamp 1679581782
transform 1 0 150912 0 1 130788
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_833
timestamp 1679581782
transform 1 0 151584 0 1 130788
box -48 -56 720 834
use sg13g2_fill_1  FILLER_78_840
timestamp 1677579658
transform 1 0 152256 0 1 130788
box -48 -56 144 834
use sg13g2_decap_8  FILLER_79_0
timestamp 1679581782
transform 1 0 71616 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_7
timestamp 1679581782
transform 1 0 72288 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_14
timestamp 1679581782
transform 1 0 72960 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_21
timestamp 1679581782
transform 1 0 73632 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_28
timestamp 1679581782
transform 1 0 74304 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_35
timestamp 1679581782
transform 1 0 74976 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_42
timestamp 1679581782
transform 1 0 75648 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_49
timestamp 1679581782
transform 1 0 76320 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_56
timestamp 1679581782
transform 1 0 76992 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_63
timestamp 1679581782
transform 1 0 77664 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_70
timestamp 1679581782
transform 1 0 78336 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_77
timestamp 1679581782
transform 1 0 79008 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_84
timestamp 1679581782
transform 1 0 79680 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_91
timestamp 1679581782
transform 1 0 80352 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_98
timestamp 1679581782
transform 1 0 81024 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_105
timestamp 1679581782
transform 1 0 81696 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_112
timestamp 1679581782
transform 1 0 82368 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_119
timestamp 1679581782
transform 1 0 83040 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_126
timestamp 1679581782
transform 1 0 83712 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_133
timestamp 1679581782
transform 1 0 84384 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_140
timestamp 1679581782
transform 1 0 85056 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_147
timestamp 1679581782
transform 1 0 85728 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_154
timestamp 1679581782
transform 1 0 86400 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_161
timestamp 1679581782
transform 1 0 87072 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_168
timestamp 1679581782
transform 1 0 87744 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_175
timestamp 1679581782
transform 1 0 88416 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_182
timestamp 1679581782
transform 1 0 89088 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_189
timestamp 1679581782
transform 1 0 89760 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_196
timestamp 1679581782
transform 1 0 90432 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_203
timestamp 1679581782
transform 1 0 91104 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_210
timestamp 1679581782
transform 1 0 91776 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_217
timestamp 1679581782
transform 1 0 92448 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_224
timestamp 1679581782
transform 1 0 93120 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_231
timestamp 1679581782
transform 1 0 93792 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_238
timestamp 1679581782
transform 1 0 94464 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_245
timestamp 1679581782
transform 1 0 95136 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_252
timestamp 1679581782
transform 1 0 95808 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_259
timestamp 1679581782
transform 1 0 96480 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_266
timestamp 1679581782
transform 1 0 97152 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_273
timestamp 1679581782
transform 1 0 97824 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_280
timestamp 1679581782
transform 1 0 98496 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_287
timestamp 1679581782
transform 1 0 99168 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_294
timestamp 1679581782
transform 1 0 99840 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_301
timestamp 1679581782
transform 1 0 100512 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_308
timestamp 1679581782
transform 1 0 101184 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_315
timestamp 1679581782
transform 1 0 101856 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_322
timestamp 1679581782
transform 1 0 102528 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_329
timestamp 1679581782
transform 1 0 103200 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_336
timestamp 1679581782
transform 1 0 103872 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_343
timestamp 1679581782
transform 1 0 104544 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_350
timestamp 1679581782
transform 1 0 105216 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_357
timestamp 1679581782
transform 1 0 105888 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_364
timestamp 1679581782
transform 1 0 106560 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_371
timestamp 1679581782
transform 1 0 107232 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_378
timestamp 1679581782
transform 1 0 107904 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_385
timestamp 1679581782
transform 1 0 108576 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_392
timestamp 1679581782
transform 1 0 109248 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_399
timestamp 1679581782
transform 1 0 109920 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_406
timestamp 1679581782
transform 1 0 110592 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_413
timestamp 1679581782
transform 1 0 111264 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_420
timestamp 1679581782
transform 1 0 111936 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_427
timestamp 1679581782
transform 1 0 112608 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_434
timestamp 1679581782
transform 1 0 113280 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_441
timestamp 1679581782
transform 1 0 113952 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_448
timestamp 1679581782
transform 1 0 114624 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_455
timestamp 1679581782
transform 1 0 115296 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_462
timestamp 1679581782
transform 1 0 115968 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_469
timestamp 1679581782
transform 1 0 116640 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_476
timestamp 1679581782
transform 1 0 117312 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_483
timestamp 1679581782
transform 1 0 117984 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_490
timestamp 1679581782
transform 1 0 118656 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_497
timestamp 1679581782
transform 1 0 119328 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_504
timestamp 1679581782
transform 1 0 120000 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_511
timestamp 1679581782
transform 1 0 120672 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_518
timestamp 1679581782
transform 1 0 121344 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_525
timestamp 1679581782
transform 1 0 122016 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_532
timestamp 1679581782
transform 1 0 122688 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_539
timestamp 1679581782
transform 1 0 123360 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_546
timestamp 1679581782
transform 1 0 124032 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_553
timestamp 1679581782
transform 1 0 124704 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_560
timestamp 1679581782
transform 1 0 125376 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_567
timestamp 1679581782
transform 1 0 126048 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_574
timestamp 1679581782
transform 1 0 126720 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_581
timestamp 1679581782
transform 1 0 127392 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_588
timestamp 1679581782
transform 1 0 128064 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_595
timestamp 1679581782
transform 1 0 128736 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_602
timestamp 1679581782
transform 1 0 129408 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_609
timestamp 1679581782
transform 1 0 130080 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_616
timestamp 1679581782
transform 1 0 130752 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_623
timestamp 1679581782
transform 1 0 131424 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_630
timestamp 1679581782
transform 1 0 132096 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_637
timestamp 1679581782
transform 1 0 132768 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_644
timestamp 1679581782
transform 1 0 133440 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_651
timestamp 1679581782
transform 1 0 134112 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_658
timestamp 1679581782
transform 1 0 134784 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_665
timestamp 1679581782
transform 1 0 135456 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_672
timestamp 1679581782
transform 1 0 136128 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_679
timestamp 1679581782
transform 1 0 136800 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_686
timestamp 1679581782
transform 1 0 137472 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_693
timestamp 1679581782
transform 1 0 138144 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_700
timestamp 1679581782
transform 1 0 138816 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_707
timestamp 1679581782
transform 1 0 139488 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_714
timestamp 1679581782
transform 1 0 140160 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_721
timestamp 1679581782
transform 1 0 140832 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_728
timestamp 1679581782
transform 1 0 141504 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_735
timestamp 1679581782
transform 1 0 142176 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_742
timestamp 1679581782
transform 1 0 142848 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_749
timestamp 1679581782
transform 1 0 143520 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_756
timestamp 1679581782
transform 1 0 144192 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_763
timestamp 1679581782
transform 1 0 144864 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_770
timestamp 1679581782
transform 1 0 145536 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_777
timestamp 1679581782
transform 1 0 146208 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_784
timestamp 1679581782
transform 1 0 146880 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_791
timestamp 1679581782
transform 1 0 147552 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_798
timestamp 1679581782
transform 1 0 148224 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_805
timestamp 1679581782
transform 1 0 148896 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_812
timestamp 1679581782
transform 1 0 149568 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_819
timestamp 1679581782
transform 1 0 150240 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_826
timestamp 1679581782
transform 1 0 150912 0 -1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_833
timestamp 1679581782
transform 1 0 151584 0 -1 132300
box -48 -56 720 834
use sg13g2_fill_1  FILLER_79_840
timestamp 1677579658
transform 1 0 152256 0 -1 132300
box -48 -56 144 834
use sg13g2_decap_8  FILLER_80_0
timestamp 1679581782
transform 1 0 71616 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_7
timestamp 1679581782
transform 1 0 72288 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_14
timestamp 1679581782
transform 1 0 72960 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_21
timestamp 1679581782
transform 1 0 73632 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_28
timestamp 1679581782
transform 1 0 74304 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_35
timestamp 1679581782
transform 1 0 74976 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_42
timestamp 1679581782
transform 1 0 75648 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_49
timestamp 1679581782
transform 1 0 76320 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_56
timestamp 1679581782
transform 1 0 76992 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_63
timestamp 1679581782
transform 1 0 77664 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_70
timestamp 1679581782
transform 1 0 78336 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_77
timestamp 1679581782
transform 1 0 79008 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_84
timestamp 1679581782
transform 1 0 79680 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_91
timestamp 1679581782
transform 1 0 80352 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_98
timestamp 1679581782
transform 1 0 81024 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_105
timestamp 1679581782
transform 1 0 81696 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_112
timestamp 1679581782
transform 1 0 82368 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_119
timestamp 1679581782
transform 1 0 83040 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_126
timestamp 1679581782
transform 1 0 83712 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_133
timestamp 1679581782
transform 1 0 84384 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_140
timestamp 1679581782
transform 1 0 85056 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_147
timestamp 1679581782
transform 1 0 85728 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_154
timestamp 1679581782
transform 1 0 86400 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_161
timestamp 1679581782
transform 1 0 87072 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_168
timestamp 1679581782
transform 1 0 87744 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_175
timestamp 1679581782
transform 1 0 88416 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_182
timestamp 1679581782
transform 1 0 89088 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_189
timestamp 1679581782
transform 1 0 89760 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_196
timestamp 1679581782
transform 1 0 90432 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_203
timestamp 1679581782
transform 1 0 91104 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_210
timestamp 1679581782
transform 1 0 91776 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_217
timestamp 1679581782
transform 1 0 92448 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_224
timestamp 1679581782
transform 1 0 93120 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_231
timestamp 1679581782
transform 1 0 93792 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_238
timestamp 1679581782
transform 1 0 94464 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_245
timestamp 1679581782
transform 1 0 95136 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_252
timestamp 1679581782
transform 1 0 95808 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_259
timestamp 1679581782
transform 1 0 96480 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_266
timestamp 1679581782
transform 1 0 97152 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_273
timestamp 1679581782
transform 1 0 97824 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_280
timestamp 1679581782
transform 1 0 98496 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_287
timestamp 1679581782
transform 1 0 99168 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_294
timestamp 1679581782
transform 1 0 99840 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_301
timestamp 1679581782
transform 1 0 100512 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_308
timestamp 1679581782
transform 1 0 101184 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_315
timestamp 1679581782
transform 1 0 101856 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_322
timestamp 1679581782
transform 1 0 102528 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_329
timestamp 1679581782
transform 1 0 103200 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_336
timestamp 1679581782
transform 1 0 103872 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_343
timestamp 1679581782
transform 1 0 104544 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_350
timestamp 1679581782
transform 1 0 105216 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_357
timestamp 1679581782
transform 1 0 105888 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_364
timestamp 1679581782
transform 1 0 106560 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_371
timestamp 1679581782
transform 1 0 107232 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_378
timestamp 1679581782
transform 1 0 107904 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_385
timestamp 1679581782
transform 1 0 108576 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_392
timestamp 1679581782
transform 1 0 109248 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_399
timestamp 1679581782
transform 1 0 109920 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_406
timestamp 1679581782
transform 1 0 110592 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_413
timestamp 1679581782
transform 1 0 111264 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_420
timestamp 1679581782
transform 1 0 111936 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_427
timestamp 1679581782
transform 1 0 112608 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_434
timestamp 1679581782
transform 1 0 113280 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_441
timestamp 1679581782
transform 1 0 113952 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_448
timestamp 1679581782
transform 1 0 114624 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_455
timestamp 1679581782
transform 1 0 115296 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_462
timestamp 1679581782
transform 1 0 115968 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_469
timestamp 1679581782
transform 1 0 116640 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_476
timestamp 1679581782
transform 1 0 117312 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_483
timestamp 1679581782
transform 1 0 117984 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_490
timestamp 1679581782
transform 1 0 118656 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_497
timestamp 1679581782
transform 1 0 119328 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_504
timestamp 1679581782
transform 1 0 120000 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_511
timestamp 1679581782
transform 1 0 120672 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_518
timestamp 1679581782
transform 1 0 121344 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_525
timestamp 1679581782
transform 1 0 122016 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_532
timestamp 1679581782
transform 1 0 122688 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_539
timestamp 1679581782
transform 1 0 123360 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_546
timestamp 1679581782
transform 1 0 124032 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_553
timestamp 1679581782
transform 1 0 124704 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_560
timestamp 1679581782
transform 1 0 125376 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_567
timestamp 1679581782
transform 1 0 126048 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_574
timestamp 1679581782
transform 1 0 126720 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_581
timestamp 1679581782
transform 1 0 127392 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_588
timestamp 1679581782
transform 1 0 128064 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_595
timestamp 1679581782
transform 1 0 128736 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_602
timestamp 1679581782
transform 1 0 129408 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_609
timestamp 1679581782
transform 1 0 130080 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_616
timestamp 1679581782
transform 1 0 130752 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_623
timestamp 1679581782
transform 1 0 131424 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_630
timestamp 1679581782
transform 1 0 132096 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_637
timestamp 1679581782
transform 1 0 132768 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_644
timestamp 1679581782
transform 1 0 133440 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_651
timestamp 1679581782
transform 1 0 134112 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_658
timestamp 1679581782
transform 1 0 134784 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_665
timestamp 1679581782
transform 1 0 135456 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_672
timestamp 1679581782
transform 1 0 136128 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_679
timestamp 1679581782
transform 1 0 136800 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_686
timestamp 1679581782
transform 1 0 137472 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_693
timestamp 1679581782
transform 1 0 138144 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_700
timestamp 1679581782
transform 1 0 138816 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_707
timestamp 1679581782
transform 1 0 139488 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_714
timestamp 1679581782
transform 1 0 140160 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_721
timestamp 1679581782
transform 1 0 140832 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_728
timestamp 1679581782
transform 1 0 141504 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_735
timestamp 1679581782
transform 1 0 142176 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_742
timestamp 1679581782
transform 1 0 142848 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_749
timestamp 1679581782
transform 1 0 143520 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_756
timestamp 1679581782
transform 1 0 144192 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_763
timestamp 1679581782
transform 1 0 144864 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_770
timestamp 1679581782
transform 1 0 145536 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_777
timestamp 1679581782
transform 1 0 146208 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_784
timestamp 1679581782
transform 1 0 146880 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_791
timestamp 1679581782
transform 1 0 147552 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_798
timestamp 1679581782
transform 1 0 148224 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_805
timestamp 1679581782
transform 1 0 148896 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_812
timestamp 1679581782
transform 1 0 149568 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_819
timestamp 1679581782
transform 1 0 150240 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_826
timestamp 1679581782
transform 1 0 150912 0 1 132300
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_833
timestamp 1679581782
transform 1 0 151584 0 1 132300
box -48 -56 720 834
use sg13g2_fill_1  FILLER_80_840
timestamp 1677579658
transform 1 0 152256 0 1 132300
box -48 -56 144 834
use sg13g2_decap_8  FILLER_81_0
timestamp 1679581782
transform 1 0 71616 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_7
timestamp 1679581782
transform 1 0 72288 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_14
timestamp 1679581782
transform 1 0 72960 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_21
timestamp 1679581782
transform 1 0 73632 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_28
timestamp 1679581782
transform 1 0 74304 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_35
timestamp 1679581782
transform 1 0 74976 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_42
timestamp 1679581782
transform 1 0 75648 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_49
timestamp 1679581782
transform 1 0 76320 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_56
timestamp 1679581782
transform 1 0 76992 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_63
timestamp 1679581782
transform 1 0 77664 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_70
timestamp 1679581782
transform 1 0 78336 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_77
timestamp 1679581782
transform 1 0 79008 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_84
timestamp 1679581782
transform 1 0 79680 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_91
timestamp 1679581782
transform 1 0 80352 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_98
timestamp 1679581782
transform 1 0 81024 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_105
timestamp 1679581782
transform 1 0 81696 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_112
timestamp 1679581782
transform 1 0 82368 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_119
timestamp 1679581782
transform 1 0 83040 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_126
timestamp 1679581782
transform 1 0 83712 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_133
timestamp 1679581782
transform 1 0 84384 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_140
timestamp 1679581782
transform 1 0 85056 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_147
timestamp 1679581782
transform 1 0 85728 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_154
timestamp 1679581782
transform 1 0 86400 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_161
timestamp 1679581782
transform 1 0 87072 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_168
timestamp 1679581782
transform 1 0 87744 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_175
timestamp 1679581782
transform 1 0 88416 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_182
timestamp 1679581782
transform 1 0 89088 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_189
timestamp 1679581782
transform 1 0 89760 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_196
timestamp 1679581782
transform 1 0 90432 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_203
timestamp 1679581782
transform 1 0 91104 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_210
timestamp 1679581782
transform 1 0 91776 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_217
timestamp 1679581782
transform 1 0 92448 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_224
timestamp 1679581782
transform 1 0 93120 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_231
timestamp 1679581782
transform 1 0 93792 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_238
timestamp 1679581782
transform 1 0 94464 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_245
timestamp 1679581782
transform 1 0 95136 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_252
timestamp 1679581782
transform 1 0 95808 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_259
timestamp 1679581782
transform 1 0 96480 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_266
timestamp 1679581782
transform 1 0 97152 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_273
timestamp 1679581782
transform 1 0 97824 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_280
timestamp 1679581782
transform 1 0 98496 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_287
timestamp 1679581782
transform 1 0 99168 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_294
timestamp 1679581782
transform 1 0 99840 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_301
timestamp 1679581782
transform 1 0 100512 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_308
timestamp 1679581782
transform 1 0 101184 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_315
timestamp 1679581782
transform 1 0 101856 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_322
timestamp 1679581782
transform 1 0 102528 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_329
timestamp 1679581782
transform 1 0 103200 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_336
timestamp 1679581782
transform 1 0 103872 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_343
timestamp 1679581782
transform 1 0 104544 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_350
timestamp 1679581782
transform 1 0 105216 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_357
timestamp 1679581782
transform 1 0 105888 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_364
timestamp 1679581782
transform 1 0 106560 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_371
timestamp 1679581782
transform 1 0 107232 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_378
timestamp 1679581782
transform 1 0 107904 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_385
timestamp 1679581782
transform 1 0 108576 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_392
timestamp 1679581782
transform 1 0 109248 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_399
timestamp 1679581782
transform 1 0 109920 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_406
timestamp 1679581782
transform 1 0 110592 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_413
timestamp 1679581782
transform 1 0 111264 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_420
timestamp 1679581782
transform 1 0 111936 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_427
timestamp 1679581782
transform 1 0 112608 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_434
timestamp 1679581782
transform 1 0 113280 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_441
timestamp 1679581782
transform 1 0 113952 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_448
timestamp 1679581782
transform 1 0 114624 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_455
timestamp 1679581782
transform 1 0 115296 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_462
timestamp 1679581782
transform 1 0 115968 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_469
timestamp 1679581782
transform 1 0 116640 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_476
timestamp 1679581782
transform 1 0 117312 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_483
timestamp 1679581782
transform 1 0 117984 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_490
timestamp 1679581782
transform 1 0 118656 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_497
timestamp 1679581782
transform 1 0 119328 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_504
timestamp 1679581782
transform 1 0 120000 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_511
timestamp 1679581782
transform 1 0 120672 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_518
timestamp 1679581782
transform 1 0 121344 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_525
timestamp 1679581782
transform 1 0 122016 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_532
timestamp 1679581782
transform 1 0 122688 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_539
timestamp 1679581782
transform 1 0 123360 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_546
timestamp 1679581782
transform 1 0 124032 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_553
timestamp 1679581782
transform 1 0 124704 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_560
timestamp 1679581782
transform 1 0 125376 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_567
timestamp 1679581782
transform 1 0 126048 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_574
timestamp 1679581782
transform 1 0 126720 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_581
timestamp 1679581782
transform 1 0 127392 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_588
timestamp 1679581782
transform 1 0 128064 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_595
timestamp 1679581782
transform 1 0 128736 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_602
timestamp 1679581782
transform 1 0 129408 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_609
timestamp 1679581782
transform 1 0 130080 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_616
timestamp 1679581782
transform 1 0 130752 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_623
timestamp 1679581782
transform 1 0 131424 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_630
timestamp 1679581782
transform 1 0 132096 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_637
timestamp 1679581782
transform 1 0 132768 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_644
timestamp 1679581782
transform 1 0 133440 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_651
timestamp 1679581782
transform 1 0 134112 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_658
timestamp 1679581782
transform 1 0 134784 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_665
timestamp 1679581782
transform 1 0 135456 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_672
timestamp 1679581782
transform 1 0 136128 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_679
timestamp 1679581782
transform 1 0 136800 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_686
timestamp 1679581782
transform 1 0 137472 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_693
timestamp 1679581782
transform 1 0 138144 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_700
timestamp 1679581782
transform 1 0 138816 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_707
timestamp 1679581782
transform 1 0 139488 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_714
timestamp 1679581782
transform 1 0 140160 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_721
timestamp 1679581782
transform 1 0 140832 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_728
timestamp 1679581782
transform 1 0 141504 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_735
timestamp 1679581782
transform 1 0 142176 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_742
timestamp 1679581782
transform 1 0 142848 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_749
timestamp 1679581782
transform 1 0 143520 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_756
timestamp 1679581782
transform 1 0 144192 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_763
timestamp 1679581782
transform 1 0 144864 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_770
timestamp 1679581782
transform 1 0 145536 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_777
timestamp 1679581782
transform 1 0 146208 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_784
timestamp 1679581782
transform 1 0 146880 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_791
timestamp 1679581782
transform 1 0 147552 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_798
timestamp 1679581782
transform 1 0 148224 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_805
timestamp 1679581782
transform 1 0 148896 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_812
timestamp 1679581782
transform 1 0 149568 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_819
timestamp 1679581782
transform 1 0 150240 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_826
timestamp 1679581782
transform 1 0 150912 0 -1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_833
timestamp 1679581782
transform 1 0 151584 0 -1 133812
box -48 -56 720 834
use sg13g2_fill_1  FILLER_81_840
timestamp 1677579658
transform 1 0 152256 0 -1 133812
box -48 -56 144 834
use sg13g2_decap_8  FILLER_82_0
timestamp 1679581782
transform 1 0 71616 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_7
timestamp 1679581782
transform 1 0 72288 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_14
timestamp 1679581782
transform 1 0 72960 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_21
timestamp 1679581782
transform 1 0 73632 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_28
timestamp 1679581782
transform 1 0 74304 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_35
timestamp 1679581782
transform 1 0 74976 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_42
timestamp 1679581782
transform 1 0 75648 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_49
timestamp 1679581782
transform 1 0 76320 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_56
timestamp 1679581782
transform 1 0 76992 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_63
timestamp 1679581782
transform 1 0 77664 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_70
timestamp 1679581782
transform 1 0 78336 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_77
timestamp 1679581782
transform 1 0 79008 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_84
timestamp 1679581782
transform 1 0 79680 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_91
timestamp 1679581782
transform 1 0 80352 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_98
timestamp 1679581782
transform 1 0 81024 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_105
timestamp 1679581782
transform 1 0 81696 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_112
timestamp 1679581782
transform 1 0 82368 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_119
timestamp 1679581782
transform 1 0 83040 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_126
timestamp 1679581782
transform 1 0 83712 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_133
timestamp 1679581782
transform 1 0 84384 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_140
timestamp 1679581782
transform 1 0 85056 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_147
timestamp 1679581782
transform 1 0 85728 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_154
timestamp 1679581782
transform 1 0 86400 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_161
timestamp 1679581782
transform 1 0 87072 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_168
timestamp 1679581782
transform 1 0 87744 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_175
timestamp 1679581782
transform 1 0 88416 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_182
timestamp 1679581782
transform 1 0 89088 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_189
timestamp 1679581782
transform 1 0 89760 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_196
timestamp 1679581782
transform 1 0 90432 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_203
timestamp 1679581782
transform 1 0 91104 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_210
timestamp 1679581782
transform 1 0 91776 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_217
timestamp 1679581782
transform 1 0 92448 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_224
timestamp 1679581782
transform 1 0 93120 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_231
timestamp 1679581782
transform 1 0 93792 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_238
timestamp 1679581782
transform 1 0 94464 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_245
timestamp 1679581782
transform 1 0 95136 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_252
timestamp 1679581782
transform 1 0 95808 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_259
timestamp 1679581782
transform 1 0 96480 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_266
timestamp 1679581782
transform 1 0 97152 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_273
timestamp 1679581782
transform 1 0 97824 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_280
timestamp 1679581782
transform 1 0 98496 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_287
timestamp 1679581782
transform 1 0 99168 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_294
timestamp 1679581782
transform 1 0 99840 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_301
timestamp 1679581782
transform 1 0 100512 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_308
timestamp 1679581782
transform 1 0 101184 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_315
timestamp 1679581782
transform 1 0 101856 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_322
timestamp 1679581782
transform 1 0 102528 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_329
timestamp 1679581782
transform 1 0 103200 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_336
timestamp 1679581782
transform 1 0 103872 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_343
timestamp 1679581782
transform 1 0 104544 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_350
timestamp 1679581782
transform 1 0 105216 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_357
timestamp 1679581782
transform 1 0 105888 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_364
timestamp 1679581782
transform 1 0 106560 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_371
timestamp 1679581782
transform 1 0 107232 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_378
timestamp 1679581782
transform 1 0 107904 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_385
timestamp 1679581782
transform 1 0 108576 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_392
timestamp 1679581782
transform 1 0 109248 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_399
timestamp 1679581782
transform 1 0 109920 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_406
timestamp 1679581782
transform 1 0 110592 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_413
timestamp 1679581782
transform 1 0 111264 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_420
timestamp 1679581782
transform 1 0 111936 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_427
timestamp 1679581782
transform 1 0 112608 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_434
timestamp 1679581782
transform 1 0 113280 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_441
timestamp 1679581782
transform 1 0 113952 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_448
timestamp 1679581782
transform 1 0 114624 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_455
timestamp 1679581782
transform 1 0 115296 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_462
timestamp 1679581782
transform 1 0 115968 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_469
timestamp 1679581782
transform 1 0 116640 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_476
timestamp 1679581782
transform 1 0 117312 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_483
timestamp 1679581782
transform 1 0 117984 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_490
timestamp 1679581782
transform 1 0 118656 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_497
timestamp 1679581782
transform 1 0 119328 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_504
timestamp 1679581782
transform 1 0 120000 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_511
timestamp 1679581782
transform 1 0 120672 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_518
timestamp 1679581782
transform 1 0 121344 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_525
timestamp 1679581782
transform 1 0 122016 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_532
timestamp 1679581782
transform 1 0 122688 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_539
timestamp 1679581782
transform 1 0 123360 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_546
timestamp 1679581782
transform 1 0 124032 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_553
timestamp 1679581782
transform 1 0 124704 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_560
timestamp 1679581782
transform 1 0 125376 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_567
timestamp 1679581782
transform 1 0 126048 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_574
timestamp 1679581782
transform 1 0 126720 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_581
timestamp 1679581782
transform 1 0 127392 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_588
timestamp 1679581782
transform 1 0 128064 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_595
timestamp 1679581782
transform 1 0 128736 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_602
timestamp 1679581782
transform 1 0 129408 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_609
timestamp 1679581782
transform 1 0 130080 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_616
timestamp 1679581782
transform 1 0 130752 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_623
timestamp 1679581782
transform 1 0 131424 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_630
timestamp 1679581782
transform 1 0 132096 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_637
timestamp 1679581782
transform 1 0 132768 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_644
timestamp 1679581782
transform 1 0 133440 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_651
timestamp 1679581782
transform 1 0 134112 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_658
timestamp 1679581782
transform 1 0 134784 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_665
timestamp 1679581782
transform 1 0 135456 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_672
timestamp 1679581782
transform 1 0 136128 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_679
timestamp 1679581782
transform 1 0 136800 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_686
timestamp 1679581782
transform 1 0 137472 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_693
timestamp 1679581782
transform 1 0 138144 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_700
timestamp 1679581782
transform 1 0 138816 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_707
timestamp 1679581782
transform 1 0 139488 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_714
timestamp 1679581782
transform 1 0 140160 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_721
timestamp 1679581782
transform 1 0 140832 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_728
timestamp 1679581782
transform 1 0 141504 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_735
timestamp 1679581782
transform 1 0 142176 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_742
timestamp 1679581782
transform 1 0 142848 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_749
timestamp 1679581782
transform 1 0 143520 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_756
timestamp 1679581782
transform 1 0 144192 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_763
timestamp 1679581782
transform 1 0 144864 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_770
timestamp 1679581782
transform 1 0 145536 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_777
timestamp 1679581782
transform 1 0 146208 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_784
timestamp 1679581782
transform 1 0 146880 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_791
timestamp 1679581782
transform 1 0 147552 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_798
timestamp 1679581782
transform 1 0 148224 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_805
timestamp 1679581782
transform 1 0 148896 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_812
timestamp 1679581782
transform 1 0 149568 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_819
timestamp 1679581782
transform 1 0 150240 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_826
timestamp 1679581782
transform 1 0 150912 0 1 133812
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_833
timestamp 1679581782
transform 1 0 151584 0 1 133812
box -48 -56 720 834
use sg13g2_fill_1  FILLER_82_840
timestamp 1677579658
transform 1 0 152256 0 1 133812
box -48 -56 144 834
use sg13g2_decap_8  FILLER_83_0
timestamp 1679581782
transform 1 0 71616 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_7
timestamp 1679581782
transform 1 0 72288 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_14
timestamp 1679581782
transform 1 0 72960 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_21
timestamp 1679581782
transform 1 0 73632 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_28
timestamp 1679581782
transform 1 0 74304 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_35
timestamp 1679581782
transform 1 0 74976 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_42
timestamp 1679581782
transform 1 0 75648 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_49
timestamp 1679581782
transform 1 0 76320 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_56
timestamp 1679581782
transform 1 0 76992 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_63
timestamp 1679581782
transform 1 0 77664 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_70
timestamp 1679581782
transform 1 0 78336 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_77
timestamp 1679581782
transform 1 0 79008 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_84
timestamp 1679581782
transform 1 0 79680 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_91
timestamp 1679581782
transform 1 0 80352 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_98
timestamp 1679581782
transform 1 0 81024 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_105
timestamp 1679581782
transform 1 0 81696 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_112
timestamp 1679581782
transform 1 0 82368 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_119
timestamp 1679581782
transform 1 0 83040 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_126
timestamp 1679581782
transform 1 0 83712 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_133
timestamp 1679581782
transform 1 0 84384 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_140
timestamp 1679581782
transform 1 0 85056 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_147
timestamp 1679581782
transform 1 0 85728 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_154
timestamp 1679581782
transform 1 0 86400 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_161
timestamp 1679581782
transform 1 0 87072 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_168
timestamp 1679581782
transform 1 0 87744 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_175
timestamp 1679581782
transform 1 0 88416 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_182
timestamp 1679581782
transform 1 0 89088 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_189
timestamp 1679581782
transform 1 0 89760 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_196
timestamp 1679581782
transform 1 0 90432 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_203
timestamp 1679581782
transform 1 0 91104 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_210
timestamp 1679581782
transform 1 0 91776 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_217
timestamp 1679581782
transform 1 0 92448 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_224
timestamp 1679581782
transform 1 0 93120 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_231
timestamp 1679581782
transform 1 0 93792 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_238
timestamp 1679581782
transform 1 0 94464 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_245
timestamp 1679581782
transform 1 0 95136 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_252
timestamp 1679581782
transform 1 0 95808 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_259
timestamp 1679581782
transform 1 0 96480 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_266
timestamp 1679581782
transform 1 0 97152 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_273
timestamp 1679581782
transform 1 0 97824 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_280
timestamp 1679581782
transform 1 0 98496 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_287
timestamp 1679581782
transform 1 0 99168 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_294
timestamp 1679581782
transform 1 0 99840 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_301
timestamp 1679581782
transform 1 0 100512 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_308
timestamp 1679581782
transform 1 0 101184 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_315
timestamp 1679581782
transform 1 0 101856 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_322
timestamp 1679581782
transform 1 0 102528 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_329
timestamp 1679581782
transform 1 0 103200 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_336
timestamp 1679581782
transform 1 0 103872 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_343
timestamp 1679581782
transform 1 0 104544 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_350
timestamp 1679581782
transform 1 0 105216 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_357
timestamp 1679581782
transform 1 0 105888 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_364
timestamp 1679581782
transform 1 0 106560 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_371
timestamp 1679581782
transform 1 0 107232 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_378
timestamp 1679581782
transform 1 0 107904 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_385
timestamp 1679581782
transform 1 0 108576 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_392
timestamp 1679581782
transform 1 0 109248 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_399
timestamp 1679581782
transform 1 0 109920 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_406
timestamp 1679581782
transform 1 0 110592 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_413
timestamp 1679581782
transform 1 0 111264 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_420
timestamp 1679581782
transform 1 0 111936 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_427
timestamp 1679581782
transform 1 0 112608 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_434
timestamp 1679581782
transform 1 0 113280 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_441
timestamp 1679581782
transform 1 0 113952 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_448
timestamp 1679581782
transform 1 0 114624 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_455
timestamp 1679581782
transform 1 0 115296 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_462
timestamp 1679581782
transform 1 0 115968 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_469
timestamp 1679581782
transform 1 0 116640 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_476
timestamp 1679581782
transform 1 0 117312 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_483
timestamp 1679581782
transform 1 0 117984 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_490
timestamp 1679581782
transform 1 0 118656 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_497
timestamp 1679581782
transform 1 0 119328 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_504
timestamp 1679581782
transform 1 0 120000 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_511
timestamp 1679581782
transform 1 0 120672 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_518
timestamp 1679581782
transform 1 0 121344 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_525
timestamp 1679581782
transform 1 0 122016 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_532
timestamp 1679581782
transform 1 0 122688 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_539
timestamp 1679581782
transform 1 0 123360 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_546
timestamp 1679581782
transform 1 0 124032 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_553
timestamp 1679581782
transform 1 0 124704 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_560
timestamp 1679581782
transform 1 0 125376 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_567
timestamp 1679581782
transform 1 0 126048 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_574
timestamp 1679581782
transform 1 0 126720 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_581
timestamp 1679581782
transform 1 0 127392 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_588
timestamp 1679581782
transform 1 0 128064 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_595
timestamp 1679581782
transform 1 0 128736 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_602
timestamp 1679581782
transform 1 0 129408 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_609
timestamp 1679581782
transform 1 0 130080 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_616
timestamp 1679581782
transform 1 0 130752 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_623
timestamp 1679581782
transform 1 0 131424 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_630
timestamp 1679581782
transform 1 0 132096 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_637
timestamp 1679581782
transform 1 0 132768 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_644
timestamp 1679581782
transform 1 0 133440 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_651
timestamp 1679581782
transform 1 0 134112 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_658
timestamp 1679581782
transform 1 0 134784 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_665
timestamp 1679581782
transform 1 0 135456 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_672
timestamp 1679581782
transform 1 0 136128 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_679
timestamp 1679581782
transform 1 0 136800 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_686
timestamp 1679581782
transform 1 0 137472 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_693
timestamp 1679581782
transform 1 0 138144 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_700
timestamp 1679581782
transform 1 0 138816 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_707
timestamp 1679581782
transform 1 0 139488 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_714
timestamp 1679581782
transform 1 0 140160 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_721
timestamp 1679581782
transform 1 0 140832 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_728
timestamp 1679581782
transform 1 0 141504 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_735
timestamp 1679581782
transform 1 0 142176 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_742
timestamp 1679581782
transform 1 0 142848 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_749
timestamp 1679581782
transform 1 0 143520 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_756
timestamp 1679581782
transform 1 0 144192 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_763
timestamp 1679581782
transform 1 0 144864 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_770
timestamp 1679581782
transform 1 0 145536 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_777
timestamp 1679581782
transform 1 0 146208 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_784
timestamp 1679581782
transform 1 0 146880 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_791
timestamp 1679581782
transform 1 0 147552 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_798
timestamp 1679581782
transform 1 0 148224 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_805
timestamp 1679581782
transform 1 0 148896 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_812
timestamp 1679581782
transform 1 0 149568 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_819
timestamp 1679581782
transform 1 0 150240 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_826
timestamp 1679581782
transform 1 0 150912 0 -1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_833
timestamp 1679581782
transform 1 0 151584 0 -1 135324
box -48 -56 720 834
use sg13g2_fill_1  FILLER_83_840
timestamp 1677579658
transform 1 0 152256 0 -1 135324
box -48 -56 144 834
use sg13g2_decap_8  FILLER_84_0
timestamp 1679581782
transform 1 0 71616 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_7
timestamp 1679581782
transform 1 0 72288 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_14
timestamp 1679581782
transform 1 0 72960 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_21
timestamp 1679581782
transform 1 0 73632 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_28
timestamp 1679581782
transform 1 0 74304 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_35
timestamp 1679581782
transform 1 0 74976 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_42
timestamp 1679581782
transform 1 0 75648 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_49
timestamp 1679581782
transform 1 0 76320 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_56
timestamp 1679581782
transform 1 0 76992 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_63
timestamp 1679581782
transform 1 0 77664 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_70
timestamp 1679581782
transform 1 0 78336 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_77
timestamp 1679581782
transform 1 0 79008 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_84
timestamp 1679581782
transform 1 0 79680 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_91
timestamp 1679581782
transform 1 0 80352 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_98
timestamp 1679581782
transform 1 0 81024 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_105
timestamp 1679581782
transform 1 0 81696 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_112
timestamp 1679581782
transform 1 0 82368 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_119
timestamp 1679581782
transform 1 0 83040 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_126
timestamp 1679581782
transform 1 0 83712 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_133
timestamp 1679581782
transform 1 0 84384 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_140
timestamp 1679581782
transform 1 0 85056 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_147
timestamp 1679581782
transform 1 0 85728 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_154
timestamp 1679581782
transform 1 0 86400 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_161
timestamp 1679581782
transform 1 0 87072 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_168
timestamp 1679581782
transform 1 0 87744 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_175
timestamp 1679581782
transform 1 0 88416 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_182
timestamp 1679581782
transform 1 0 89088 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_189
timestamp 1679581782
transform 1 0 89760 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_196
timestamp 1679581782
transform 1 0 90432 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_203
timestamp 1679581782
transform 1 0 91104 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_210
timestamp 1679581782
transform 1 0 91776 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_217
timestamp 1679581782
transform 1 0 92448 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_224
timestamp 1679581782
transform 1 0 93120 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_231
timestamp 1679581782
transform 1 0 93792 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_238
timestamp 1679581782
transform 1 0 94464 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_245
timestamp 1679581782
transform 1 0 95136 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_252
timestamp 1679581782
transform 1 0 95808 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_259
timestamp 1679581782
transform 1 0 96480 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_266
timestamp 1679581782
transform 1 0 97152 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_273
timestamp 1679581782
transform 1 0 97824 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_280
timestamp 1679581782
transform 1 0 98496 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_287
timestamp 1679581782
transform 1 0 99168 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_294
timestamp 1679581782
transform 1 0 99840 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_301
timestamp 1679581782
transform 1 0 100512 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_308
timestamp 1679581782
transform 1 0 101184 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_315
timestamp 1679581782
transform 1 0 101856 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_322
timestamp 1679581782
transform 1 0 102528 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_329
timestamp 1679581782
transform 1 0 103200 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_336
timestamp 1679581782
transform 1 0 103872 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_343
timestamp 1679581782
transform 1 0 104544 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_350
timestamp 1679581782
transform 1 0 105216 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_357
timestamp 1679581782
transform 1 0 105888 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_364
timestamp 1679581782
transform 1 0 106560 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_371
timestamp 1679581782
transform 1 0 107232 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_378
timestamp 1679581782
transform 1 0 107904 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_385
timestamp 1679581782
transform 1 0 108576 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_392
timestamp 1679581782
transform 1 0 109248 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_399
timestamp 1679581782
transform 1 0 109920 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_406
timestamp 1679581782
transform 1 0 110592 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_413
timestamp 1679581782
transform 1 0 111264 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_420
timestamp 1679581782
transform 1 0 111936 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_427
timestamp 1679581782
transform 1 0 112608 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_434
timestamp 1679581782
transform 1 0 113280 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_441
timestamp 1679581782
transform 1 0 113952 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_448
timestamp 1679581782
transform 1 0 114624 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_455
timestamp 1679581782
transform 1 0 115296 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_462
timestamp 1679581782
transform 1 0 115968 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_469
timestamp 1679581782
transform 1 0 116640 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_476
timestamp 1679581782
transform 1 0 117312 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_483
timestamp 1679581782
transform 1 0 117984 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_490
timestamp 1679581782
transform 1 0 118656 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_497
timestamp 1679581782
transform 1 0 119328 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_504
timestamp 1679581782
transform 1 0 120000 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_511
timestamp 1679581782
transform 1 0 120672 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_518
timestamp 1679581782
transform 1 0 121344 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_525
timestamp 1679581782
transform 1 0 122016 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_532
timestamp 1679581782
transform 1 0 122688 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_539
timestamp 1679581782
transform 1 0 123360 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_546
timestamp 1679581782
transform 1 0 124032 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_553
timestamp 1679581782
transform 1 0 124704 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_560
timestamp 1679581782
transform 1 0 125376 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_567
timestamp 1679581782
transform 1 0 126048 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_574
timestamp 1679581782
transform 1 0 126720 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_581
timestamp 1679581782
transform 1 0 127392 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_588
timestamp 1679581782
transform 1 0 128064 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_595
timestamp 1679581782
transform 1 0 128736 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_602
timestamp 1679581782
transform 1 0 129408 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_609
timestamp 1679581782
transform 1 0 130080 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_616
timestamp 1679581782
transform 1 0 130752 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_623
timestamp 1679581782
transform 1 0 131424 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_630
timestamp 1679581782
transform 1 0 132096 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_637
timestamp 1679581782
transform 1 0 132768 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_644
timestamp 1679581782
transform 1 0 133440 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_651
timestamp 1679581782
transform 1 0 134112 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_658
timestamp 1679581782
transform 1 0 134784 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_665
timestamp 1679581782
transform 1 0 135456 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_672
timestamp 1679581782
transform 1 0 136128 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_679
timestamp 1679581782
transform 1 0 136800 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_686
timestamp 1679581782
transform 1 0 137472 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_693
timestamp 1679581782
transform 1 0 138144 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_700
timestamp 1679581782
transform 1 0 138816 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_707
timestamp 1679581782
transform 1 0 139488 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_714
timestamp 1679581782
transform 1 0 140160 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_721
timestamp 1679581782
transform 1 0 140832 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_728
timestamp 1679581782
transform 1 0 141504 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_735
timestamp 1679581782
transform 1 0 142176 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_742
timestamp 1679581782
transform 1 0 142848 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_749
timestamp 1679581782
transform 1 0 143520 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_756
timestamp 1679581782
transform 1 0 144192 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_763
timestamp 1679581782
transform 1 0 144864 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_770
timestamp 1679581782
transform 1 0 145536 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_777
timestamp 1679581782
transform 1 0 146208 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_784
timestamp 1679581782
transform 1 0 146880 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_791
timestamp 1679581782
transform 1 0 147552 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_798
timestamp 1679581782
transform 1 0 148224 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_805
timestamp 1679581782
transform 1 0 148896 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_812
timestamp 1679581782
transform 1 0 149568 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_819
timestamp 1679581782
transform 1 0 150240 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_826
timestamp 1679581782
transform 1 0 150912 0 1 135324
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_833
timestamp 1679581782
transform 1 0 151584 0 1 135324
box -48 -56 720 834
use sg13g2_fill_1  FILLER_84_840
timestamp 1677579658
transform 1 0 152256 0 1 135324
box -48 -56 144 834
use sg13g2_decap_8  FILLER_85_0
timestamp 1679581782
transform 1 0 71616 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_7
timestamp 1679581782
transform 1 0 72288 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_14
timestamp 1679581782
transform 1 0 72960 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_21
timestamp 1679581782
transform 1 0 73632 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_28
timestamp 1679581782
transform 1 0 74304 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_35
timestamp 1679581782
transform 1 0 74976 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_42
timestamp 1679581782
transform 1 0 75648 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_49
timestamp 1679581782
transform 1 0 76320 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_56
timestamp 1679581782
transform 1 0 76992 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_63
timestamp 1679581782
transform 1 0 77664 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_70
timestamp 1679581782
transform 1 0 78336 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_77
timestamp 1679581782
transform 1 0 79008 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_84
timestamp 1679581782
transform 1 0 79680 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_91
timestamp 1679581782
transform 1 0 80352 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_98
timestamp 1679581782
transform 1 0 81024 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_105
timestamp 1679581782
transform 1 0 81696 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_112
timestamp 1679581782
transform 1 0 82368 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_119
timestamp 1679581782
transform 1 0 83040 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_126
timestamp 1679581782
transform 1 0 83712 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_133
timestamp 1679581782
transform 1 0 84384 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_140
timestamp 1679581782
transform 1 0 85056 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_147
timestamp 1679581782
transform 1 0 85728 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_154
timestamp 1679581782
transform 1 0 86400 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_161
timestamp 1679581782
transform 1 0 87072 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_168
timestamp 1679581782
transform 1 0 87744 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_175
timestamp 1679581782
transform 1 0 88416 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_182
timestamp 1679581782
transform 1 0 89088 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_189
timestamp 1679581782
transform 1 0 89760 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_196
timestamp 1679581782
transform 1 0 90432 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_203
timestamp 1679581782
transform 1 0 91104 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_210
timestamp 1679581782
transform 1 0 91776 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_217
timestamp 1679581782
transform 1 0 92448 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_224
timestamp 1679581782
transform 1 0 93120 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_231
timestamp 1679581782
transform 1 0 93792 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_238
timestamp 1679581782
transform 1 0 94464 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_245
timestamp 1679581782
transform 1 0 95136 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_252
timestamp 1679581782
transform 1 0 95808 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_259
timestamp 1679581782
transform 1 0 96480 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_266
timestamp 1679581782
transform 1 0 97152 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_273
timestamp 1679581782
transform 1 0 97824 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_280
timestamp 1679581782
transform 1 0 98496 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_287
timestamp 1679581782
transform 1 0 99168 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_294
timestamp 1679581782
transform 1 0 99840 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_301
timestamp 1679581782
transform 1 0 100512 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_308
timestamp 1679581782
transform 1 0 101184 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_315
timestamp 1679581782
transform 1 0 101856 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_322
timestamp 1679581782
transform 1 0 102528 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_329
timestamp 1679581782
transform 1 0 103200 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_336
timestamp 1679581782
transform 1 0 103872 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_343
timestamp 1679581782
transform 1 0 104544 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_350
timestamp 1679581782
transform 1 0 105216 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_357
timestamp 1679581782
transform 1 0 105888 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_364
timestamp 1679581782
transform 1 0 106560 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_371
timestamp 1679581782
transform 1 0 107232 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_378
timestamp 1679581782
transform 1 0 107904 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_385
timestamp 1679581782
transform 1 0 108576 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_392
timestamp 1679581782
transform 1 0 109248 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_399
timestamp 1679581782
transform 1 0 109920 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_406
timestamp 1679581782
transform 1 0 110592 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_413
timestamp 1679581782
transform 1 0 111264 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_420
timestamp 1679581782
transform 1 0 111936 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_427
timestamp 1679581782
transform 1 0 112608 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_434
timestamp 1679581782
transform 1 0 113280 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_441
timestamp 1679581782
transform 1 0 113952 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_448
timestamp 1679581782
transform 1 0 114624 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_455
timestamp 1679581782
transform 1 0 115296 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_462
timestamp 1679581782
transform 1 0 115968 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_469
timestamp 1679581782
transform 1 0 116640 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_476
timestamp 1679581782
transform 1 0 117312 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_483
timestamp 1679581782
transform 1 0 117984 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_490
timestamp 1679581782
transform 1 0 118656 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_497
timestamp 1679581782
transform 1 0 119328 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_504
timestamp 1679581782
transform 1 0 120000 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_511
timestamp 1679581782
transform 1 0 120672 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_518
timestamp 1679581782
transform 1 0 121344 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_525
timestamp 1679581782
transform 1 0 122016 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_532
timestamp 1679581782
transform 1 0 122688 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_539
timestamp 1679581782
transform 1 0 123360 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_546
timestamp 1679581782
transform 1 0 124032 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_553
timestamp 1679581782
transform 1 0 124704 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_560
timestamp 1679581782
transform 1 0 125376 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_567
timestamp 1679581782
transform 1 0 126048 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_574
timestamp 1679581782
transform 1 0 126720 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_581
timestamp 1679581782
transform 1 0 127392 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_588
timestamp 1679581782
transform 1 0 128064 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_595
timestamp 1679581782
transform 1 0 128736 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_602
timestamp 1679581782
transform 1 0 129408 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_609
timestamp 1679581782
transform 1 0 130080 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_616
timestamp 1679581782
transform 1 0 130752 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_623
timestamp 1679581782
transform 1 0 131424 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_630
timestamp 1679581782
transform 1 0 132096 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_637
timestamp 1679581782
transform 1 0 132768 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_644
timestamp 1679581782
transform 1 0 133440 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_651
timestamp 1679581782
transform 1 0 134112 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_658
timestamp 1679581782
transform 1 0 134784 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_665
timestamp 1679581782
transform 1 0 135456 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_672
timestamp 1679581782
transform 1 0 136128 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_679
timestamp 1679581782
transform 1 0 136800 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_686
timestamp 1679581782
transform 1 0 137472 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_693
timestamp 1679581782
transform 1 0 138144 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_700
timestamp 1679581782
transform 1 0 138816 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_707
timestamp 1679581782
transform 1 0 139488 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_714
timestamp 1679581782
transform 1 0 140160 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_721
timestamp 1679581782
transform 1 0 140832 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_728
timestamp 1679581782
transform 1 0 141504 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_735
timestamp 1679581782
transform 1 0 142176 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_742
timestamp 1679581782
transform 1 0 142848 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_749
timestamp 1679581782
transform 1 0 143520 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_756
timestamp 1679581782
transform 1 0 144192 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_763
timestamp 1679581782
transform 1 0 144864 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_770
timestamp 1679581782
transform 1 0 145536 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_777
timestamp 1679581782
transform 1 0 146208 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_784
timestamp 1679581782
transform 1 0 146880 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_791
timestamp 1679581782
transform 1 0 147552 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_798
timestamp 1679581782
transform 1 0 148224 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_805
timestamp 1679581782
transform 1 0 148896 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_812
timestamp 1679581782
transform 1 0 149568 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_819
timestamp 1679581782
transform 1 0 150240 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_826
timestamp 1679581782
transform 1 0 150912 0 -1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_833
timestamp 1679581782
transform 1 0 151584 0 -1 136836
box -48 -56 720 834
use sg13g2_fill_1  FILLER_85_840
timestamp 1677579658
transform 1 0 152256 0 -1 136836
box -48 -56 144 834
use sg13g2_decap_8  FILLER_86_0
timestamp 1679581782
transform 1 0 71616 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_7
timestamp 1679581782
transform 1 0 72288 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_14
timestamp 1679581782
transform 1 0 72960 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_21
timestamp 1679581782
transform 1 0 73632 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_28
timestamp 1679581782
transform 1 0 74304 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_35
timestamp 1679581782
transform 1 0 74976 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_42
timestamp 1679581782
transform 1 0 75648 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_49
timestamp 1679581782
transform 1 0 76320 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_56
timestamp 1679581782
transform 1 0 76992 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_63
timestamp 1679581782
transform 1 0 77664 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_70
timestamp 1679581782
transform 1 0 78336 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_77
timestamp 1679581782
transform 1 0 79008 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_84
timestamp 1679581782
transform 1 0 79680 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_91
timestamp 1679581782
transform 1 0 80352 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_98
timestamp 1679581782
transform 1 0 81024 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_105
timestamp 1679581782
transform 1 0 81696 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_112
timestamp 1679581782
transform 1 0 82368 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_119
timestamp 1679581782
transform 1 0 83040 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_126
timestamp 1679581782
transform 1 0 83712 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_133
timestamp 1679581782
transform 1 0 84384 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_140
timestamp 1679581782
transform 1 0 85056 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_147
timestamp 1679581782
transform 1 0 85728 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_154
timestamp 1679581782
transform 1 0 86400 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_161
timestamp 1679581782
transform 1 0 87072 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_168
timestamp 1679581782
transform 1 0 87744 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_175
timestamp 1679581782
transform 1 0 88416 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_182
timestamp 1679581782
transform 1 0 89088 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_189
timestamp 1679581782
transform 1 0 89760 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_196
timestamp 1679581782
transform 1 0 90432 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_203
timestamp 1679581782
transform 1 0 91104 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_210
timestamp 1679581782
transform 1 0 91776 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_217
timestamp 1679581782
transform 1 0 92448 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_224
timestamp 1679581782
transform 1 0 93120 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_231
timestamp 1679581782
transform 1 0 93792 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_238
timestamp 1679581782
transform 1 0 94464 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_245
timestamp 1679581782
transform 1 0 95136 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_252
timestamp 1679581782
transform 1 0 95808 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_259
timestamp 1679581782
transform 1 0 96480 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_266
timestamp 1679581782
transform 1 0 97152 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_273
timestamp 1679581782
transform 1 0 97824 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_280
timestamp 1679581782
transform 1 0 98496 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_287
timestamp 1679581782
transform 1 0 99168 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_294
timestamp 1679581782
transform 1 0 99840 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_301
timestamp 1679581782
transform 1 0 100512 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_308
timestamp 1679581782
transform 1 0 101184 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_315
timestamp 1679581782
transform 1 0 101856 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_322
timestamp 1679581782
transform 1 0 102528 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_329
timestamp 1679581782
transform 1 0 103200 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_336
timestamp 1679581782
transform 1 0 103872 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_343
timestamp 1679581782
transform 1 0 104544 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_350
timestamp 1679581782
transform 1 0 105216 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_357
timestamp 1679581782
transform 1 0 105888 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_364
timestamp 1679581782
transform 1 0 106560 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_371
timestamp 1679581782
transform 1 0 107232 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_378
timestamp 1679581782
transform 1 0 107904 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_385
timestamp 1679581782
transform 1 0 108576 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_392
timestamp 1679581782
transform 1 0 109248 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_399
timestamp 1679581782
transform 1 0 109920 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_406
timestamp 1679581782
transform 1 0 110592 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_413
timestamp 1679581782
transform 1 0 111264 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_420
timestamp 1679581782
transform 1 0 111936 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_427
timestamp 1679581782
transform 1 0 112608 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_434
timestamp 1679581782
transform 1 0 113280 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_441
timestamp 1679581782
transform 1 0 113952 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_448
timestamp 1679581782
transform 1 0 114624 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_455
timestamp 1679581782
transform 1 0 115296 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_462
timestamp 1679581782
transform 1 0 115968 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_469
timestamp 1679581782
transform 1 0 116640 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_476
timestamp 1679581782
transform 1 0 117312 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_483
timestamp 1679581782
transform 1 0 117984 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_490
timestamp 1679581782
transform 1 0 118656 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_497
timestamp 1679581782
transform 1 0 119328 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_504
timestamp 1679581782
transform 1 0 120000 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_511
timestamp 1679581782
transform 1 0 120672 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_518
timestamp 1679581782
transform 1 0 121344 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_525
timestamp 1679581782
transform 1 0 122016 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_532
timestamp 1679581782
transform 1 0 122688 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_539
timestamp 1679581782
transform 1 0 123360 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_546
timestamp 1679581782
transform 1 0 124032 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_553
timestamp 1679581782
transform 1 0 124704 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_560
timestamp 1679581782
transform 1 0 125376 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_567
timestamp 1679581782
transform 1 0 126048 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_574
timestamp 1679581782
transform 1 0 126720 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_581
timestamp 1679581782
transform 1 0 127392 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_588
timestamp 1679581782
transform 1 0 128064 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_595
timestamp 1679581782
transform 1 0 128736 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_602
timestamp 1679581782
transform 1 0 129408 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_609
timestamp 1679581782
transform 1 0 130080 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_616
timestamp 1679581782
transform 1 0 130752 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_623
timestamp 1679581782
transform 1 0 131424 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_630
timestamp 1679581782
transform 1 0 132096 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_637
timestamp 1679581782
transform 1 0 132768 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_644
timestamp 1679581782
transform 1 0 133440 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_651
timestamp 1679581782
transform 1 0 134112 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_658
timestamp 1679581782
transform 1 0 134784 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_665
timestamp 1679581782
transform 1 0 135456 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_672
timestamp 1679581782
transform 1 0 136128 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_679
timestamp 1679581782
transform 1 0 136800 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_686
timestamp 1679581782
transform 1 0 137472 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_693
timestamp 1679581782
transform 1 0 138144 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_700
timestamp 1679581782
transform 1 0 138816 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_707
timestamp 1679581782
transform 1 0 139488 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_714
timestamp 1679581782
transform 1 0 140160 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_721
timestamp 1679581782
transform 1 0 140832 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_728
timestamp 1679581782
transform 1 0 141504 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_735
timestamp 1679581782
transform 1 0 142176 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_742
timestamp 1679581782
transform 1 0 142848 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_749
timestamp 1679581782
transform 1 0 143520 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_756
timestamp 1679581782
transform 1 0 144192 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_763
timestamp 1679581782
transform 1 0 144864 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_770
timestamp 1679581782
transform 1 0 145536 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_777
timestamp 1679581782
transform 1 0 146208 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_784
timestamp 1679581782
transform 1 0 146880 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_791
timestamp 1679581782
transform 1 0 147552 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_798
timestamp 1679581782
transform 1 0 148224 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_805
timestamp 1679581782
transform 1 0 148896 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_812
timestamp 1679581782
transform 1 0 149568 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_819
timestamp 1679581782
transform 1 0 150240 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_826
timestamp 1679581782
transform 1 0 150912 0 1 136836
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_833
timestamp 1679581782
transform 1 0 151584 0 1 136836
box -48 -56 720 834
use sg13g2_fill_1  FILLER_86_840
timestamp 1677579658
transform 1 0 152256 0 1 136836
box -48 -56 144 834
use sg13g2_decap_8  FILLER_87_0
timestamp 1679581782
transform 1 0 71616 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_7
timestamp 1679581782
transform 1 0 72288 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_14
timestamp 1679581782
transform 1 0 72960 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_21
timestamp 1679581782
transform 1 0 73632 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_28
timestamp 1679581782
transform 1 0 74304 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_35
timestamp 1679581782
transform 1 0 74976 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_42
timestamp 1679581782
transform 1 0 75648 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_49
timestamp 1679581782
transform 1 0 76320 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_56
timestamp 1679581782
transform 1 0 76992 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_63
timestamp 1679581782
transform 1 0 77664 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_70
timestamp 1679581782
transform 1 0 78336 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_77
timestamp 1679581782
transform 1 0 79008 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_84
timestamp 1679581782
transform 1 0 79680 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_91
timestamp 1679581782
transform 1 0 80352 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_98
timestamp 1679581782
transform 1 0 81024 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_105
timestamp 1679581782
transform 1 0 81696 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_112
timestamp 1679581782
transform 1 0 82368 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_119
timestamp 1679581782
transform 1 0 83040 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_126
timestamp 1679581782
transform 1 0 83712 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_133
timestamp 1679581782
transform 1 0 84384 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_140
timestamp 1679581782
transform 1 0 85056 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_147
timestamp 1679581782
transform 1 0 85728 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_154
timestamp 1679581782
transform 1 0 86400 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_161
timestamp 1679581782
transform 1 0 87072 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_168
timestamp 1679581782
transform 1 0 87744 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_175
timestamp 1679581782
transform 1 0 88416 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_182
timestamp 1679581782
transform 1 0 89088 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_189
timestamp 1679581782
transform 1 0 89760 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_196
timestamp 1679581782
transform 1 0 90432 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_203
timestamp 1679581782
transform 1 0 91104 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_210
timestamp 1679581782
transform 1 0 91776 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_217
timestamp 1679581782
transform 1 0 92448 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_224
timestamp 1679581782
transform 1 0 93120 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_231
timestamp 1679581782
transform 1 0 93792 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_238
timestamp 1679581782
transform 1 0 94464 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_245
timestamp 1679581782
transform 1 0 95136 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_252
timestamp 1679581782
transform 1 0 95808 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_259
timestamp 1679581782
transform 1 0 96480 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_266
timestamp 1679581782
transform 1 0 97152 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_273
timestamp 1679581782
transform 1 0 97824 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_280
timestamp 1679581782
transform 1 0 98496 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_287
timestamp 1679581782
transform 1 0 99168 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_294
timestamp 1679581782
transform 1 0 99840 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_301
timestamp 1679581782
transform 1 0 100512 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_308
timestamp 1679581782
transform 1 0 101184 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_315
timestamp 1679581782
transform 1 0 101856 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_322
timestamp 1679581782
transform 1 0 102528 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_329
timestamp 1679581782
transform 1 0 103200 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_336
timestamp 1679581782
transform 1 0 103872 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_343
timestamp 1679581782
transform 1 0 104544 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_350
timestamp 1679581782
transform 1 0 105216 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_357
timestamp 1679581782
transform 1 0 105888 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_364
timestamp 1679581782
transform 1 0 106560 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_371
timestamp 1679581782
transform 1 0 107232 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_378
timestamp 1679581782
transform 1 0 107904 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_385
timestamp 1679581782
transform 1 0 108576 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_392
timestamp 1679581782
transform 1 0 109248 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_399
timestamp 1679581782
transform 1 0 109920 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_406
timestamp 1679581782
transform 1 0 110592 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_413
timestamp 1679581782
transform 1 0 111264 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_420
timestamp 1679581782
transform 1 0 111936 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_427
timestamp 1679581782
transform 1 0 112608 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_434
timestamp 1679581782
transform 1 0 113280 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_441
timestamp 1679581782
transform 1 0 113952 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_448
timestamp 1679581782
transform 1 0 114624 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_455
timestamp 1679581782
transform 1 0 115296 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_462
timestamp 1679581782
transform 1 0 115968 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_469
timestamp 1679581782
transform 1 0 116640 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_476
timestamp 1679581782
transform 1 0 117312 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_483
timestamp 1679581782
transform 1 0 117984 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_490
timestamp 1679581782
transform 1 0 118656 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_497
timestamp 1679581782
transform 1 0 119328 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_504
timestamp 1679581782
transform 1 0 120000 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_511
timestamp 1679581782
transform 1 0 120672 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_518
timestamp 1679581782
transform 1 0 121344 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_525
timestamp 1679581782
transform 1 0 122016 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_532
timestamp 1679581782
transform 1 0 122688 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_539
timestamp 1679581782
transform 1 0 123360 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_546
timestamp 1679581782
transform 1 0 124032 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_553
timestamp 1679581782
transform 1 0 124704 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_560
timestamp 1679581782
transform 1 0 125376 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_567
timestamp 1679581782
transform 1 0 126048 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_574
timestamp 1679581782
transform 1 0 126720 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_581
timestamp 1679581782
transform 1 0 127392 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_588
timestamp 1679581782
transform 1 0 128064 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_595
timestamp 1679581782
transform 1 0 128736 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_602
timestamp 1679581782
transform 1 0 129408 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_609
timestamp 1679581782
transform 1 0 130080 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_616
timestamp 1679581782
transform 1 0 130752 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_623
timestamp 1679581782
transform 1 0 131424 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_630
timestamp 1679581782
transform 1 0 132096 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_637
timestamp 1679581782
transform 1 0 132768 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_644
timestamp 1679581782
transform 1 0 133440 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_651
timestamp 1679581782
transform 1 0 134112 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_658
timestamp 1679581782
transform 1 0 134784 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_665
timestamp 1679581782
transform 1 0 135456 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_672
timestamp 1679581782
transform 1 0 136128 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_679
timestamp 1679581782
transform 1 0 136800 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_686
timestamp 1679581782
transform 1 0 137472 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_693
timestamp 1679581782
transform 1 0 138144 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_700
timestamp 1679581782
transform 1 0 138816 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_707
timestamp 1679581782
transform 1 0 139488 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_714
timestamp 1679581782
transform 1 0 140160 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_721
timestamp 1679581782
transform 1 0 140832 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_728
timestamp 1679581782
transform 1 0 141504 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_735
timestamp 1679581782
transform 1 0 142176 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_742
timestamp 1679581782
transform 1 0 142848 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_749
timestamp 1679581782
transform 1 0 143520 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_756
timestamp 1679581782
transform 1 0 144192 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_763
timestamp 1679581782
transform 1 0 144864 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_770
timestamp 1679581782
transform 1 0 145536 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_777
timestamp 1679581782
transform 1 0 146208 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_784
timestamp 1679581782
transform 1 0 146880 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_791
timestamp 1679581782
transform 1 0 147552 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_798
timestamp 1679581782
transform 1 0 148224 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_805
timestamp 1679581782
transform 1 0 148896 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_812
timestamp 1679581782
transform 1 0 149568 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_819
timestamp 1679581782
transform 1 0 150240 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_826
timestamp 1679581782
transform 1 0 150912 0 -1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_833
timestamp 1679581782
transform 1 0 151584 0 -1 138348
box -48 -56 720 834
use sg13g2_fill_1  FILLER_87_840
timestamp 1677579658
transform 1 0 152256 0 -1 138348
box -48 -56 144 834
use sg13g2_decap_8  FILLER_88_0
timestamp 1679581782
transform 1 0 71616 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_7
timestamp 1679581782
transform 1 0 72288 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_14
timestamp 1679581782
transform 1 0 72960 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_21
timestamp 1679581782
transform 1 0 73632 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_28
timestamp 1679581782
transform 1 0 74304 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_35
timestamp 1679581782
transform 1 0 74976 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_42
timestamp 1679581782
transform 1 0 75648 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_49
timestamp 1679581782
transform 1 0 76320 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_56
timestamp 1679581782
transform 1 0 76992 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_63
timestamp 1679581782
transform 1 0 77664 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_70
timestamp 1679581782
transform 1 0 78336 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_77
timestamp 1679581782
transform 1 0 79008 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_84
timestamp 1679581782
transform 1 0 79680 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_91
timestamp 1679581782
transform 1 0 80352 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_98
timestamp 1679581782
transform 1 0 81024 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_105
timestamp 1679581782
transform 1 0 81696 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_112
timestamp 1679581782
transform 1 0 82368 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_119
timestamp 1679581782
transform 1 0 83040 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_126
timestamp 1679581782
transform 1 0 83712 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_133
timestamp 1679581782
transform 1 0 84384 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_140
timestamp 1679581782
transform 1 0 85056 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_147
timestamp 1679581782
transform 1 0 85728 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_154
timestamp 1679581782
transform 1 0 86400 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_161
timestamp 1679581782
transform 1 0 87072 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_168
timestamp 1679581782
transform 1 0 87744 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_175
timestamp 1679581782
transform 1 0 88416 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_182
timestamp 1679581782
transform 1 0 89088 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_189
timestamp 1679581782
transform 1 0 89760 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_196
timestamp 1679581782
transform 1 0 90432 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_203
timestamp 1679581782
transform 1 0 91104 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_210
timestamp 1679581782
transform 1 0 91776 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_217
timestamp 1679581782
transform 1 0 92448 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_224
timestamp 1679581782
transform 1 0 93120 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_231
timestamp 1679581782
transform 1 0 93792 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_238
timestamp 1679581782
transform 1 0 94464 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_245
timestamp 1679581782
transform 1 0 95136 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_252
timestamp 1679581782
transform 1 0 95808 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_259
timestamp 1679581782
transform 1 0 96480 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_266
timestamp 1679581782
transform 1 0 97152 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_273
timestamp 1679581782
transform 1 0 97824 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_280
timestamp 1679581782
transform 1 0 98496 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_287
timestamp 1679581782
transform 1 0 99168 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_294
timestamp 1679581782
transform 1 0 99840 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_301
timestamp 1679581782
transform 1 0 100512 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_308
timestamp 1679581782
transform 1 0 101184 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_315
timestamp 1679581782
transform 1 0 101856 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_322
timestamp 1679581782
transform 1 0 102528 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_329
timestamp 1679581782
transform 1 0 103200 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_336
timestamp 1679581782
transform 1 0 103872 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_343
timestamp 1679581782
transform 1 0 104544 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_350
timestamp 1679581782
transform 1 0 105216 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_357
timestamp 1679581782
transform 1 0 105888 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_364
timestamp 1679581782
transform 1 0 106560 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_371
timestamp 1679581782
transform 1 0 107232 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_378
timestamp 1679581782
transform 1 0 107904 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_385
timestamp 1679581782
transform 1 0 108576 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_392
timestamp 1679581782
transform 1 0 109248 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_399
timestamp 1679581782
transform 1 0 109920 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_406
timestamp 1679581782
transform 1 0 110592 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_413
timestamp 1679581782
transform 1 0 111264 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_420
timestamp 1679581782
transform 1 0 111936 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_427
timestamp 1679581782
transform 1 0 112608 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_434
timestamp 1679581782
transform 1 0 113280 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_441
timestamp 1679581782
transform 1 0 113952 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_448
timestamp 1679581782
transform 1 0 114624 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_455
timestamp 1679581782
transform 1 0 115296 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_462
timestamp 1679581782
transform 1 0 115968 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_469
timestamp 1679581782
transform 1 0 116640 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_476
timestamp 1679581782
transform 1 0 117312 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_483
timestamp 1679581782
transform 1 0 117984 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_490
timestamp 1679581782
transform 1 0 118656 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_497
timestamp 1679581782
transform 1 0 119328 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_504
timestamp 1679581782
transform 1 0 120000 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_511
timestamp 1679581782
transform 1 0 120672 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_518
timestamp 1679581782
transform 1 0 121344 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_525
timestamp 1679581782
transform 1 0 122016 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_532
timestamp 1679581782
transform 1 0 122688 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_539
timestamp 1679581782
transform 1 0 123360 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_546
timestamp 1679581782
transform 1 0 124032 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_553
timestamp 1679581782
transform 1 0 124704 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_560
timestamp 1679581782
transform 1 0 125376 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_567
timestamp 1679581782
transform 1 0 126048 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_574
timestamp 1679581782
transform 1 0 126720 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_581
timestamp 1679581782
transform 1 0 127392 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_588
timestamp 1679581782
transform 1 0 128064 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_595
timestamp 1679581782
transform 1 0 128736 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_602
timestamp 1679581782
transform 1 0 129408 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_609
timestamp 1679581782
transform 1 0 130080 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_616
timestamp 1679581782
transform 1 0 130752 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_623
timestamp 1679581782
transform 1 0 131424 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_630
timestamp 1679581782
transform 1 0 132096 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_637
timestamp 1679581782
transform 1 0 132768 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_644
timestamp 1679581782
transform 1 0 133440 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_651
timestamp 1679581782
transform 1 0 134112 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_658
timestamp 1679581782
transform 1 0 134784 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_665
timestamp 1679581782
transform 1 0 135456 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_672
timestamp 1679581782
transform 1 0 136128 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_679
timestamp 1679581782
transform 1 0 136800 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_686
timestamp 1679581782
transform 1 0 137472 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_693
timestamp 1679581782
transform 1 0 138144 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_700
timestamp 1679581782
transform 1 0 138816 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_707
timestamp 1679581782
transform 1 0 139488 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_714
timestamp 1679581782
transform 1 0 140160 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_721
timestamp 1679581782
transform 1 0 140832 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_728
timestamp 1679581782
transform 1 0 141504 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_735
timestamp 1679581782
transform 1 0 142176 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_742
timestamp 1679581782
transform 1 0 142848 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_749
timestamp 1679581782
transform 1 0 143520 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_756
timestamp 1679581782
transform 1 0 144192 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_763
timestamp 1679581782
transform 1 0 144864 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_770
timestamp 1679581782
transform 1 0 145536 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_777
timestamp 1679581782
transform 1 0 146208 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_784
timestamp 1679581782
transform 1 0 146880 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_791
timestamp 1679581782
transform 1 0 147552 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_798
timestamp 1679581782
transform 1 0 148224 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_805
timestamp 1679581782
transform 1 0 148896 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_812
timestamp 1679581782
transform 1 0 149568 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_819
timestamp 1679581782
transform 1 0 150240 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_826
timestamp 1679581782
transform 1 0 150912 0 1 138348
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_833
timestamp 1679581782
transform 1 0 151584 0 1 138348
box -48 -56 720 834
use sg13g2_fill_1  FILLER_88_840
timestamp 1677579658
transform 1 0 152256 0 1 138348
box -48 -56 144 834
use sg13g2_decap_8  FILLER_89_0
timestamp 1679581782
transform 1 0 71616 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_7
timestamp 1679581782
transform 1 0 72288 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_14
timestamp 1679581782
transform 1 0 72960 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_21
timestamp 1679581782
transform 1 0 73632 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_28
timestamp 1679581782
transform 1 0 74304 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_35
timestamp 1679581782
transform 1 0 74976 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_42
timestamp 1679581782
transform 1 0 75648 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_49
timestamp 1679581782
transform 1 0 76320 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_56
timestamp 1679581782
transform 1 0 76992 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_63
timestamp 1679581782
transform 1 0 77664 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_70
timestamp 1679581782
transform 1 0 78336 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_77
timestamp 1679581782
transform 1 0 79008 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_84
timestamp 1679581782
transform 1 0 79680 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_91
timestamp 1679581782
transform 1 0 80352 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_98
timestamp 1679581782
transform 1 0 81024 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_105
timestamp 1679581782
transform 1 0 81696 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_112
timestamp 1679581782
transform 1 0 82368 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_119
timestamp 1679581782
transform 1 0 83040 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_126
timestamp 1679581782
transform 1 0 83712 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_133
timestamp 1679581782
transform 1 0 84384 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_140
timestamp 1679581782
transform 1 0 85056 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_147
timestamp 1679581782
transform 1 0 85728 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_154
timestamp 1679581782
transform 1 0 86400 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_161
timestamp 1679581782
transform 1 0 87072 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_168
timestamp 1679581782
transform 1 0 87744 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_175
timestamp 1679581782
transform 1 0 88416 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_182
timestamp 1679581782
transform 1 0 89088 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_189
timestamp 1679581782
transform 1 0 89760 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_196
timestamp 1679581782
transform 1 0 90432 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_203
timestamp 1679581782
transform 1 0 91104 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_210
timestamp 1679581782
transform 1 0 91776 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_217
timestamp 1679581782
transform 1 0 92448 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_224
timestamp 1679581782
transform 1 0 93120 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_231
timestamp 1679581782
transform 1 0 93792 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_238
timestamp 1679581782
transform 1 0 94464 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_245
timestamp 1679581782
transform 1 0 95136 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_252
timestamp 1679581782
transform 1 0 95808 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_259
timestamp 1679581782
transform 1 0 96480 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_266
timestamp 1679581782
transform 1 0 97152 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_273
timestamp 1679581782
transform 1 0 97824 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_280
timestamp 1679581782
transform 1 0 98496 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_287
timestamp 1679581782
transform 1 0 99168 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_294
timestamp 1679581782
transform 1 0 99840 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_301
timestamp 1679581782
transform 1 0 100512 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_308
timestamp 1679581782
transform 1 0 101184 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_315
timestamp 1679581782
transform 1 0 101856 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_322
timestamp 1679581782
transform 1 0 102528 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_329
timestamp 1679581782
transform 1 0 103200 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_336
timestamp 1679581782
transform 1 0 103872 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_343
timestamp 1679581782
transform 1 0 104544 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_350
timestamp 1679581782
transform 1 0 105216 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_357
timestamp 1679581782
transform 1 0 105888 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_364
timestamp 1679581782
transform 1 0 106560 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_371
timestamp 1679581782
transform 1 0 107232 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_378
timestamp 1679581782
transform 1 0 107904 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_385
timestamp 1679581782
transform 1 0 108576 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_392
timestamp 1679581782
transform 1 0 109248 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_399
timestamp 1679581782
transform 1 0 109920 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_406
timestamp 1679581782
transform 1 0 110592 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_413
timestamp 1679581782
transform 1 0 111264 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_420
timestamp 1679581782
transform 1 0 111936 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_427
timestamp 1679581782
transform 1 0 112608 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_434
timestamp 1679581782
transform 1 0 113280 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_441
timestamp 1679581782
transform 1 0 113952 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_448
timestamp 1679581782
transform 1 0 114624 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_455
timestamp 1679581782
transform 1 0 115296 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_462
timestamp 1679581782
transform 1 0 115968 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_469
timestamp 1679581782
transform 1 0 116640 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_476
timestamp 1679581782
transform 1 0 117312 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_483
timestamp 1679581782
transform 1 0 117984 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_490
timestamp 1679581782
transform 1 0 118656 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_497
timestamp 1679581782
transform 1 0 119328 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_504
timestamp 1679581782
transform 1 0 120000 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_511
timestamp 1679581782
transform 1 0 120672 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_518
timestamp 1679581782
transform 1 0 121344 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_525
timestamp 1679581782
transform 1 0 122016 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_532
timestamp 1679581782
transform 1 0 122688 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_539
timestamp 1679581782
transform 1 0 123360 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_546
timestamp 1679581782
transform 1 0 124032 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_553
timestamp 1679581782
transform 1 0 124704 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_560
timestamp 1679581782
transform 1 0 125376 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_567
timestamp 1679581782
transform 1 0 126048 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_574
timestamp 1679581782
transform 1 0 126720 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_581
timestamp 1679581782
transform 1 0 127392 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_588
timestamp 1679581782
transform 1 0 128064 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_595
timestamp 1679581782
transform 1 0 128736 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_602
timestamp 1679581782
transform 1 0 129408 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_609
timestamp 1679581782
transform 1 0 130080 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_616
timestamp 1679581782
transform 1 0 130752 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_623
timestamp 1679581782
transform 1 0 131424 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_630
timestamp 1679581782
transform 1 0 132096 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_637
timestamp 1679581782
transform 1 0 132768 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_644
timestamp 1679581782
transform 1 0 133440 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_651
timestamp 1679581782
transform 1 0 134112 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_658
timestamp 1679581782
transform 1 0 134784 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_665
timestamp 1679581782
transform 1 0 135456 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_672
timestamp 1679581782
transform 1 0 136128 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_679
timestamp 1679581782
transform 1 0 136800 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_686
timestamp 1679581782
transform 1 0 137472 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_693
timestamp 1679581782
transform 1 0 138144 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_700
timestamp 1679581782
transform 1 0 138816 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_707
timestamp 1679581782
transform 1 0 139488 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_714
timestamp 1679581782
transform 1 0 140160 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_721
timestamp 1679581782
transform 1 0 140832 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_728
timestamp 1679581782
transform 1 0 141504 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_735
timestamp 1679581782
transform 1 0 142176 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_742
timestamp 1679581782
transform 1 0 142848 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_749
timestamp 1679581782
transform 1 0 143520 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_756
timestamp 1679581782
transform 1 0 144192 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_763
timestamp 1679581782
transform 1 0 144864 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_770
timestamp 1679581782
transform 1 0 145536 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_777
timestamp 1679581782
transform 1 0 146208 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_784
timestamp 1679581782
transform 1 0 146880 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_791
timestamp 1679581782
transform 1 0 147552 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_798
timestamp 1679581782
transform 1 0 148224 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_805
timestamp 1679581782
transform 1 0 148896 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_812
timestamp 1679581782
transform 1 0 149568 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_819
timestamp 1679581782
transform 1 0 150240 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_826
timestamp 1679581782
transform 1 0 150912 0 -1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_833
timestamp 1679581782
transform 1 0 151584 0 -1 139860
box -48 -56 720 834
use sg13g2_fill_1  FILLER_89_840
timestamp 1677579658
transform 1 0 152256 0 -1 139860
box -48 -56 144 834
use sg13g2_decap_8  FILLER_90_0
timestamp 1679581782
transform 1 0 71616 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_7
timestamp 1679581782
transform 1 0 72288 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_14
timestamp 1679581782
transform 1 0 72960 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_21
timestamp 1679581782
transform 1 0 73632 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_28
timestamp 1679581782
transform 1 0 74304 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_35
timestamp 1679581782
transform 1 0 74976 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_42
timestamp 1679581782
transform 1 0 75648 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_49
timestamp 1679581782
transform 1 0 76320 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_56
timestamp 1679581782
transform 1 0 76992 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_63
timestamp 1679581782
transform 1 0 77664 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_70
timestamp 1679581782
transform 1 0 78336 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_77
timestamp 1679581782
transform 1 0 79008 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_84
timestamp 1679581782
transform 1 0 79680 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_91
timestamp 1679581782
transform 1 0 80352 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_98
timestamp 1679581782
transform 1 0 81024 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_105
timestamp 1679581782
transform 1 0 81696 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_112
timestamp 1679581782
transform 1 0 82368 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_119
timestamp 1679581782
transform 1 0 83040 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_126
timestamp 1679581782
transform 1 0 83712 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_133
timestamp 1679581782
transform 1 0 84384 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_140
timestamp 1679581782
transform 1 0 85056 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_147
timestamp 1679581782
transform 1 0 85728 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_154
timestamp 1679581782
transform 1 0 86400 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_161
timestamp 1679581782
transform 1 0 87072 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_168
timestamp 1679581782
transform 1 0 87744 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_175
timestamp 1679581782
transform 1 0 88416 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_182
timestamp 1679581782
transform 1 0 89088 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_189
timestamp 1679581782
transform 1 0 89760 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_196
timestamp 1679581782
transform 1 0 90432 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_203
timestamp 1679581782
transform 1 0 91104 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_210
timestamp 1679581782
transform 1 0 91776 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_217
timestamp 1679581782
transform 1 0 92448 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_224
timestamp 1679581782
transform 1 0 93120 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_231
timestamp 1679581782
transform 1 0 93792 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_238
timestamp 1679581782
transform 1 0 94464 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_245
timestamp 1679581782
transform 1 0 95136 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_252
timestamp 1679581782
transform 1 0 95808 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_259
timestamp 1679581782
transform 1 0 96480 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_266
timestamp 1679581782
transform 1 0 97152 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_273
timestamp 1679581782
transform 1 0 97824 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_280
timestamp 1679581782
transform 1 0 98496 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_287
timestamp 1679581782
transform 1 0 99168 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_294
timestamp 1679581782
transform 1 0 99840 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_301
timestamp 1679581782
transform 1 0 100512 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_308
timestamp 1679581782
transform 1 0 101184 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_315
timestamp 1679581782
transform 1 0 101856 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_322
timestamp 1679581782
transform 1 0 102528 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_329
timestamp 1679581782
transform 1 0 103200 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_336
timestamp 1679581782
transform 1 0 103872 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_343
timestamp 1679581782
transform 1 0 104544 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_350
timestamp 1679581782
transform 1 0 105216 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_357
timestamp 1679581782
transform 1 0 105888 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_364
timestamp 1679581782
transform 1 0 106560 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_371
timestamp 1679581782
transform 1 0 107232 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_378
timestamp 1679581782
transform 1 0 107904 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_385
timestamp 1679581782
transform 1 0 108576 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_392
timestamp 1679581782
transform 1 0 109248 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_399
timestamp 1679581782
transform 1 0 109920 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_406
timestamp 1679581782
transform 1 0 110592 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_413
timestamp 1679581782
transform 1 0 111264 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_420
timestamp 1679581782
transform 1 0 111936 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_427
timestamp 1679581782
transform 1 0 112608 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_434
timestamp 1679581782
transform 1 0 113280 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_441
timestamp 1679581782
transform 1 0 113952 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_448
timestamp 1679581782
transform 1 0 114624 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_455
timestamp 1679581782
transform 1 0 115296 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_462
timestamp 1679581782
transform 1 0 115968 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_469
timestamp 1679581782
transform 1 0 116640 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_476
timestamp 1679581782
transform 1 0 117312 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_483
timestamp 1679581782
transform 1 0 117984 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_490
timestamp 1679581782
transform 1 0 118656 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_497
timestamp 1679581782
transform 1 0 119328 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_504
timestamp 1679581782
transform 1 0 120000 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_511
timestamp 1679581782
transform 1 0 120672 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_518
timestamp 1679581782
transform 1 0 121344 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_525
timestamp 1679581782
transform 1 0 122016 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_532
timestamp 1679581782
transform 1 0 122688 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_539
timestamp 1679581782
transform 1 0 123360 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_546
timestamp 1679581782
transform 1 0 124032 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_553
timestamp 1679581782
transform 1 0 124704 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_560
timestamp 1679581782
transform 1 0 125376 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_567
timestamp 1679581782
transform 1 0 126048 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_574
timestamp 1679581782
transform 1 0 126720 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_581
timestamp 1679581782
transform 1 0 127392 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_588
timestamp 1679581782
transform 1 0 128064 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_595
timestamp 1679581782
transform 1 0 128736 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_602
timestamp 1679581782
transform 1 0 129408 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_609
timestamp 1679581782
transform 1 0 130080 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_616
timestamp 1679581782
transform 1 0 130752 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_623
timestamp 1679581782
transform 1 0 131424 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_630
timestamp 1679581782
transform 1 0 132096 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_637
timestamp 1679581782
transform 1 0 132768 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_644
timestamp 1679581782
transform 1 0 133440 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_651
timestamp 1679581782
transform 1 0 134112 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_658
timestamp 1679581782
transform 1 0 134784 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_665
timestamp 1679581782
transform 1 0 135456 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_672
timestamp 1679581782
transform 1 0 136128 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_679
timestamp 1679581782
transform 1 0 136800 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_686
timestamp 1679581782
transform 1 0 137472 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_693
timestamp 1679581782
transform 1 0 138144 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_700
timestamp 1679581782
transform 1 0 138816 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_707
timestamp 1679581782
transform 1 0 139488 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_714
timestamp 1679581782
transform 1 0 140160 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_721
timestamp 1679581782
transform 1 0 140832 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_728
timestamp 1679581782
transform 1 0 141504 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_735
timestamp 1679581782
transform 1 0 142176 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_742
timestamp 1679581782
transform 1 0 142848 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_749
timestamp 1679581782
transform 1 0 143520 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_756
timestamp 1679581782
transform 1 0 144192 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_763
timestamp 1679581782
transform 1 0 144864 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_770
timestamp 1679581782
transform 1 0 145536 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_777
timestamp 1679581782
transform 1 0 146208 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_784
timestamp 1679581782
transform 1 0 146880 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_791
timestamp 1679581782
transform 1 0 147552 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_798
timestamp 1679581782
transform 1 0 148224 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_805
timestamp 1679581782
transform 1 0 148896 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_812
timestamp 1679581782
transform 1 0 149568 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_819
timestamp 1679581782
transform 1 0 150240 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_826
timestamp 1679581782
transform 1 0 150912 0 1 139860
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_833
timestamp 1679581782
transform 1 0 151584 0 1 139860
box -48 -56 720 834
use sg13g2_fill_1  FILLER_90_840
timestamp 1677579658
transform 1 0 152256 0 1 139860
box -48 -56 144 834
use sg13g2_decap_8  FILLER_91_0
timestamp 1679581782
transform 1 0 71616 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_7
timestamp 1679581782
transform 1 0 72288 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_14
timestamp 1679581782
transform 1 0 72960 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_21
timestamp 1679581782
transform 1 0 73632 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_28
timestamp 1679581782
transform 1 0 74304 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_35
timestamp 1679581782
transform 1 0 74976 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_42
timestamp 1679581782
transform 1 0 75648 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_49
timestamp 1679581782
transform 1 0 76320 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_56
timestamp 1679581782
transform 1 0 76992 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_63
timestamp 1679581782
transform 1 0 77664 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_70
timestamp 1679581782
transform 1 0 78336 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_77
timestamp 1679581782
transform 1 0 79008 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_84
timestamp 1679581782
transform 1 0 79680 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_91
timestamp 1679581782
transform 1 0 80352 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_98
timestamp 1679581782
transform 1 0 81024 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_105
timestamp 1679581782
transform 1 0 81696 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_112
timestamp 1679581782
transform 1 0 82368 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_119
timestamp 1679581782
transform 1 0 83040 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_126
timestamp 1679581782
transform 1 0 83712 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_133
timestamp 1679581782
transform 1 0 84384 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_140
timestamp 1679581782
transform 1 0 85056 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_147
timestamp 1679581782
transform 1 0 85728 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_154
timestamp 1679581782
transform 1 0 86400 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_161
timestamp 1679581782
transform 1 0 87072 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_168
timestamp 1679581782
transform 1 0 87744 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_175
timestamp 1679581782
transform 1 0 88416 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_182
timestamp 1679581782
transform 1 0 89088 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_189
timestamp 1679581782
transform 1 0 89760 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_196
timestamp 1679581782
transform 1 0 90432 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_203
timestamp 1679581782
transform 1 0 91104 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_210
timestamp 1679581782
transform 1 0 91776 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_217
timestamp 1679581782
transform 1 0 92448 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_224
timestamp 1679581782
transform 1 0 93120 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_231
timestamp 1679581782
transform 1 0 93792 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_238
timestamp 1679581782
transform 1 0 94464 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_245
timestamp 1679581782
transform 1 0 95136 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_252
timestamp 1679581782
transform 1 0 95808 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_259
timestamp 1679581782
transform 1 0 96480 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_266
timestamp 1679581782
transform 1 0 97152 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_273
timestamp 1679581782
transform 1 0 97824 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_280
timestamp 1679581782
transform 1 0 98496 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_287
timestamp 1679581782
transform 1 0 99168 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_294
timestamp 1679581782
transform 1 0 99840 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_301
timestamp 1679581782
transform 1 0 100512 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_308
timestamp 1679581782
transform 1 0 101184 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_315
timestamp 1679581782
transform 1 0 101856 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_322
timestamp 1679581782
transform 1 0 102528 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_329
timestamp 1679581782
transform 1 0 103200 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_336
timestamp 1679581782
transform 1 0 103872 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_343
timestamp 1679581782
transform 1 0 104544 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_350
timestamp 1679581782
transform 1 0 105216 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_357
timestamp 1679581782
transform 1 0 105888 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_364
timestamp 1679581782
transform 1 0 106560 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_371
timestamp 1679581782
transform 1 0 107232 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_378
timestamp 1679581782
transform 1 0 107904 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_385
timestamp 1679581782
transform 1 0 108576 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_392
timestamp 1679581782
transform 1 0 109248 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_399
timestamp 1679581782
transform 1 0 109920 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_406
timestamp 1679581782
transform 1 0 110592 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_413
timestamp 1679581782
transform 1 0 111264 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_420
timestamp 1679581782
transform 1 0 111936 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_427
timestamp 1679581782
transform 1 0 112608 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_434
timestamp 1679581782
transform 1 0 113280 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_441
timestamp 1679581782
transform 1 0 113952 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_448
timestamp 1679581782
transform 1 0 114624 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_455
timestamp 1679581782
transform 1 0 115296 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_462
timestamp 1679581782
transform 1 0 115968 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_469
timestamp 1679581782
transform 1 0 116640 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_476
timestamp 1679581782
transform 1 0 117312 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_483
timestamp 1679581782
transform 1 0 117984 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_490
timestamp 1679581782
transform 1 0 118656 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_497
timestamp 1679581782
transform 1 0 119328 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_504
timestamp 1679581782
transform 1 0 120000 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_511
timestamp 1679581782
transform 1 0 120672 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_518
timestamp 1679581782
transform 1 0 121344 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_525
timestamp 1679581782
transform 1 0 122016 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_532
timestamp 1679581782
transform 1 0 122688 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_539
timestamp 1679581782
transform 1 0 123360 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_546
timestamp 1679581782
transform 1 0 124032 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_553
timestamp 1679581782
transform 1 0 124704 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_560
timestamp 1679581782
transform 1 0 125376 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_567
timestamp 1679581782
transform 1 0 126048 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_574
timestamp 1679581782
transform 1 0 126720 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_581
timestamp 1679581782
transform 1 0 127392 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_588
timestamp 1679581782
transform 1 0 128064 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_595
timestamp 1679581782
transform 1 0 128736 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_602
timestamp 1679581782
transform 1 0 129408 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_609
timestamp 1679581782
transform 1 0 130080 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_616
timestamp 1679581782
transform 1 0 130752 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_623
timestamp 1679581782
transform 1 0 131424 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_630
timestamp 1679581782
transform 1 0 132096 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_637
timestamp 1679581782
transform 1 0 132768 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_644
timestamp 1679581782
transform 1 0 133440 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_651
timestamp 1679581782
transform 1 0 134112 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_658
timestamp 1679581782
transform 1 0 134784 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_665
timestamp 1679581782
transform 1 0 135456 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_672
timestamp 1679581782
transform 1 0 136128 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_679
timestamp 1679581782
transform 1 0 136800 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_686
timestamp 1679581782
transform 1 0 137472 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_693
timestamp 1679581782
transform 1 0 138144 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_700
timestamp 1679581782
transform 1 0 138816 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_707
timestamp 1679581782
transform 1 0 139488 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_714
timestamp 1679581782
transform 1 0 140160 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_721
timestamp 1679581782
transform 1 0 140832 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_728
timestamp 1679581782
transform 1 0 141504 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_735
timestamp 1679581782
transform 1 0 142176 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_742
timestamp 1679581782
transform 1 0 142848 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_749
timestamp 1679581782
transform 1 0 143520 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_756
timestamp 1679581782
transform 1 0 144192 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_763
timestamp 1679581782
transform 1 0 144864 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_770
timestamp 1679581782
transform 1 0 145536 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_777
timestamp 1679581782
transform 1 0 146208 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_784
timestamp 1679581782
transform 1 0 146880 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_791
timestamp 1679581782
transform 1 0 147552 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_798
timestamp 1679581782
transform 1 0 148224 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_805
timestamp 1679581782
transform 1 0 148896 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_812
timestamp 1679581782
transform 1 0 149568 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_819
timestamp 1679581782
transform 1 0 150240 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_826
timestamp 1679581782
transform 1 0 150912 0 -1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_833
timestamp 1679581782
transform 1 0 151584 0 -1 141372
box -48 -56 720 834
use sg13g2_fill_1  FILLER_91_840
timestamp 1677579658
transform 1 0 152256 0 -1 141372
box -48 -56 144 834
use sg13g2_decap_8  FILLER_92_0
timestamp 1679581782
transform 1 0 71616 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_7
timestamp 1679581782
transform 1 0 72288 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_14
timestamp 1679581782
transform 1 0 72960 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_21
timestamp 1679581782
transform 1 0 73632 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_28
timestamp 1679581782
transform 1 0 74304 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_35
timestamp 1679581782
transform 1 0 74976 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_42
timestamp 1679581782
transform 1 0 75648 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_49
timestamp 1679581782
transform 1 0 76320 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_56
timestamp 1679581782
transform 1 0 76992 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_63
timestamp 1679581782
transform 1 0 77664 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_70
timestamp 1679581782
transform 1 0 78336 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_77
timestamp 1679581782
transform 1 0 79008 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_84
timestamp 1679581782
transform 1 0 79680 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_91
timestamp 1679581782
transform 1 0 80352 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_98
timestamp 1679581782
transform 1 0 81024 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_105
timestamp 1679581782
transform 1 0 81696 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_112
timestamp 1679581782
transform 1 0 82368 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_119
timestamp 1679581782
transform 1 0 83040 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_126
timestamp 1679581782
transform 1 0 83712 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_133
timestamp 1679581782
transform 1 0 84384 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_140
timestamp 1679581782
transform 1 0 85056 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_147
timestamp 1679581782
transform 1 0 85728 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_154
timestamp 1679581782
transform 1 0 86400 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_161
timestamp 1679581782
transform 1 0 87072 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_168
timestamp 1679581782
transform 1 0 87744 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_175
timestamp 1679581782
transform 1 0 88416 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_182
timestamp 1679581782
transform 1 0 89088 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_189
timestamp 1679581782
transform 1 0 89760 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_196
timestamp 1679581782
transform 1 0 90432 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_203
timestamp 1679581782
transform 1 0 91104 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_210
timestamp 1679581782
transform 1 0 91776 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_217
timestamp 1679581782
transform 1 0 92448 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_224
timestamp 1679581782
transform 1 0 93120 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_231
timestamp 1679581782
transform 1 0 93792 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_238
timestamp 1679581782
transform 1 0 94464 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_245
timestamp 1679581782
transform 1 0 95136 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_252
timestamp 1679581782
transform 1 0 95808 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_259
timestamp 1679581782
transform 1 0 96480 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_266
timestamp 1679581782
transform 1 0 97152 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_273
timestamp 1679581782
transform 1 0 97824 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_280
timestamp 1679581782
transform 1 0 98496 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_287
timestamp 1679581782
transform 1 0 99168 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_294
timestamp 1679581782
transform 1 0 99840 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_301
timestamp 1679581782
transform 1 0 100512 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_308
timestamp 1679581782
transform 1 0 101184 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_315
timestamp 1679581782
transform 1 0 101856 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_322
timestamp 1679581782
transform 1 0 102528 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_329
timestamp 1679581782
transform 1 0 103200 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_336
timestamp 1679581782
transform 1 0 103872 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_343
timestamp 1679581782
transform 1 0 104544 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_350
timestamp 1679581782
transform 1 0 105216 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_357
timestamp 1679581782
transform 1 0 105888 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_364
timestamp 1679581782
transform 1 0 106560 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_371
timestamp 1679581782
transform 1 0 107232 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_378
timestamp 1679581782
transform 1 0 107904 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_385
timestamp 1679581782
transform 1 0 108576 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_392
timestamp 1679581782
transform 1 0 109248 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_399
timestamp 1679581782
transform 1 0 109920 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_406
timestamp 1679581782
transform 1 0 110592 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_413
timestamp 1679581782
transform 1 0 111264 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_420
timestamp 1679581782
transform 1 0 111936 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_427
timestamp 1679581782
transform 1 0 112608 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_434
timestamp 1679581782
transform 1 0 113280 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_441
timestamp 1679581782
transform 1 0 113952 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_448
timestamp 1679581782
transform 1 0 114624 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_455
timestamp 1679581782
transform 1 0 115296 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_462
timestamp 1679581782
transform 1 0 115968 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_469
timestamp 1679581782
transform 1 0 116640 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_476
timestamp 1679581782
transform 1 0 117312 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_483
timestamp 1679581782
transform 1 0 117984 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_490
timestamp 1679581782
transform 1 0 118656 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_497
timestamp 1679581782
transform 1 0 119328 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_504
timestamp 1679581782
transform 1 0 120000 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_511
timestamp 1679581782
transform 1 0 120672 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_518
timestamp 1679581782
transform 1 0 121344 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_525
timestamp 1679581782
transform 1 0 122016 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_532
timestamp 1679581782
transform 1 0 122688 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_539
timestamp 1679581782
transform 1 0 123360 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_546
timestamp 1679581782
transform 1 0 124032 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_553
timestamp 1679581782
transform 1 0 124704 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_560
timestamp 1679581782
transform 1 0 125376 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_567
timestamp 1679581782
transform 1 0 126048 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_574
timestamp 1679581782
transform 1 0 126720 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_581
timestamp 1679581782
transform 1 0 127392 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_588
timestamp 1679581782
transform 1 0 128064 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_595
timestamp 1679581782
transform 1 0 128736 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_602
timestamp 1679581782
transform 1 0 129408 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_609
timestamp 1679581782
transform 1 0 130080 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_616
timestamp 1679581782
transform 1 0 130752 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_623
timestamp 1679581782
transform 1 0 131424 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_630
timestamp 1679581782
transform 1 0 132096 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_637
timestamp 1679581782
transform 1 0 132768 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_644
timestamp 1679581782
transform 1 0 133440 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_651
timestamp 1679581782
transform 1 0 134112 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_658
timestamp 1679581782
transform 1 0 134784 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_665
timestamp 1679581782
transform 1 0 135456 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_672
timestamp 1679581782
transform 1 0 136128 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_679
timestamp 1679581782
transform 1 0 136800 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_686
timestamp 1679581782
transform 1 0 137472 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_693
timestamp 1679581782
transform 1 0 138144 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_700
timestamp 1679581782
transform 1 0 138816 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_707
timestamp 1679581782
transform 1 0 139488 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_714
timestamp 1679581782
transform 1 0 140160 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_721
timestamp 1679581782
transform 1 0 140832 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_728
timestamp 1679581782
transform 1 0 141504 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_735
timestamp 1679581782
transform 1 0 142176 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_742
timestamp 1679581782
transform 1 0 142848 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_749
timestamp 1679581782
transform 1 0 143520 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_756
timestamp 1679581782
transform 1 0 144192 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_763
timestamp 1679581782
transform 1 0 144864 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_770
timestamp 1679581782
transform 1 0 145536 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_777
timestamp 1679581782
transform 1 0 146208 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_784
timestamp 1679581782
transform 1 0 146880 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_791
timestamp 1679581782
transform 1 0 147552 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_798
timestamp 1679581782
transform 1 0 148224 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_805
timestamp 1679581782
transform 1 0 148896 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_812
timestamp 1679581782
transform 1 0 149568 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_819
timestamp 1679581782
transform 1 0 150240 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_826
timestamp 1679581782
transform 1 0 150912 0 1 141372
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_833
timestamp 1679581782
transform 1 0 151584 0 1 141372
box -48 -56 720 834
use sg13g2_fill_1  FILLER_92_840
timestamp 1677579658
transform 1 0 152256 0 1 141372
box -48 -56 144 834
use sg13g2_decap_8  FILLER_93_0
timestamp 1679581782
transform 1 0 71616 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_7
timestamp 1679581782
transform 1 0 72288 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_14
timestamp 1679581782
transform 1 0 72960 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_21
timestamp 1679581782
transform 1 0 73632 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_28
timestamp 1679581782
transform 1 0 74304 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_35
timestamp 1679581782
transform 1 0 74976 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_42
timestamp 1679581782
transform 1 0 75648 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_49
timestamp 1679581782
transform 1 0 76320 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_56
timestamp 1679581782
transform 1 0 76992 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_63
timestamp 1679581782
transform 1 0 77664 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_70
timestamp 1679581782
transform 1 0 78336 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_77
timestamp 1679581782
transform 1 0 79008 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_84
timestamp 1679581782
transform 1 0 79680 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_91
timestamp 1679581782
transform 1 0 80352 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_98
timestamp 1679581782
transform 1 0 81024 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_105
timestamp 1679581782
transform 1 0 81696 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_112
timestamp 1679581782
transform 1 0 82368 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_119
timestamp 1679581782
transform 1 0 83040 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_126
timestamp 1679581782
transform 1 0 83712 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_133
timestamp 1679581782
transform 1 0 84384 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_140
timestamp 1679581782
transform 1 0 85056 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_147
timestamp 1679581782
transform 1 0 85728 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_154
timestamp 1679581782
transform 1 0 86400 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_161
timestamp 1679581782
transform 1 0 87072 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_168
timestamp 1679581782
transform 1 0 87744 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_175
timestamp 1679581782
transform 1 0 88416 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_182
timestamp 1679581782
transform 1 0 89088 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_189
timestamp 1679581782
transform 1 0 89760 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_196
timestamp 1679581782
transform 1 0 90432 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_203
timestamp 1679581782
transform 1 0 91104 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_210
timestamp 1679581782
transform 1 0 91776 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_217
timestamp 1679581782
transform 1 0 92448 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_224
timestamp 1679581782
transform 1 0 93120 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_231
timestamp 1679581782
transform 1 0 93792 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_238
timestamp 1679581782
transform 1 0 94464 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_245
timestamp 1679581782
transform 1 0 95136 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_252
timestamp 1679581782
transform 1 0 95808 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_259
timestamp 1679581782
transform 1 0 96480 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_266
timestamp 1679581782
transform 1 0 97152 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_273
timestamp 1679581782
transform 1 0 97824 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_280
timestamp 1679581782
transform 1 0 98496 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_287
timestamp 1679581782
transform 1 0 99168 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_294
timestamp 1679581782
transform 1 0 99840 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_301
timestamp 1679581782
transform 1 0 100512 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_308
timestamp 1679581782
transform 1 0 101184 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_315
timestamp 1679581782
transform 1 0 101856 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_322
timestamp 1679581782
transform 1 0 102528 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_329
timestamp 1679581782
transform 1 0 103200 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_336
timestamp 1679581782
transform 1 0 103872 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_343
timestamp 1679581782
transform 1 0 104544 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_350
timestamp 1679581782
transform 1 0 105216 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_357
timestamp 1679581782
transform 1 0 105888 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_364
timestamp 1679581782
transform 1 0 106560 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_371
timestamp 1679581782
transform 1 0 107232 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_378
timestamp 1679581782
transform 1 0 107904 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_385
timestamp 1679581782
transform 1 0 108576 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_392
timestamp 1679581782
transform 1 0 109248 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_399
timestamp 1679581782
transform 1 0 109920 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_406
timestamp 1679581782
transform 1 0 110592 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_413
timestamp 1679581782
transform 1 0 111264 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_420
timestamp 1679581782
transform 1 0 111936 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_427
timestamp 1679581782
transform 1 0 112608 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_434
timestamp 1679581782
transform 1 0 113280 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_441
timestamp 1679581782
transform 1 0 113952 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_448
timestamp 1679581782
transform 1 0 114624 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_455
timestamp 1679581782
transform 1 0 115296 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_462
timestamp 1679581782
transform 1 0 115968 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_469
timestamp 1679581782
transform 1 0 116640 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_476
timestamp 1679581782
transform 1 0 117312 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_483
timestamp 1679581782
transform 1 0 117984 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_490
timestamp 1679581782
transform 1 0 118656 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_497
timestamp 1679581782
transform 1 0 119328 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_504
timestamp 1679581782
transform 1 0 120000 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_511
timestamp 1679581782
transform 1 0 120672 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_518
timestamp 1679581782
transform 1 0 121344 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_525
timestamp 1679581782
transform 1 0 122016 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_532
timestamp 1679581782
transform 1 0 122688 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_539
timestamp 1679581782
transform 1 0 123360 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_546
timestamp 1679581782
transform 1 0 124032 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_553
timestamp 1679581782
transform 1 0 124704 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_560
timestamp 1679581782
transform 1 0 125376 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_567
timestamp 1679581782
transform 1 0 126048 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_574
timestamp 1679581782
transform 1 0 126720 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_581
timestamp 1679581782
transform 1 0 127392 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_588
timestamp 1679581782
transform 1 0 128064 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_595
timestamp 1679581782
transform 1 0 128736 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_602
timestamp 1679581782
transform 1 0 129408 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_609
timestamp 1679581782
transform 1 0 130080 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_616
timestamp 1679581782
transform 1 0 130752 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_623
timestamp 1679581782
transform 1 0 131424 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_630
timestamp 1679581782
transform 1 0 132096 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_637
timestamp 1679581782
transform 1 0 132768 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_644
timestamp 1679581782
transform 1 0 133440 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_651
timestamp 1679581782
transform 1 0 134112 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_658
timestamp 1679581782
transform 1 0 134784 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_665
timestamp 1679581782
transform 1 0 135456 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_672
timestamp 1679581782
transform 1 0 136128 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_679
timestamp 1679581782
transform 1 0 136800 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_686
timestamp 1679581782
transform 1 0 137472 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_693
timestamp 1679581782
transform 1 0 138144 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_700
timestamp 1679581782
transform 1 0 138816 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_707
timestamp 1679581782
transform 1 0 139488 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_714
timestamp 1679581782
transform 1 0 140160 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_721
timestamp 1679581782
transform 1 0 140832 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_728
timestamp 1679581782
transform 1 0 141504 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_735
timestamp 1679581782
transform 1 0 142176 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_742
timestamp 1679581782
transform 1 0 142848 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_749
timestamp 1679581782
transform 1 0 143520 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_756
timestamp 1679581782
transform 1 0 144192 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_763
timestamp 1679581782
transform 1 0 144864 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_770
timestamp 1679581782
transform 1 0 145536 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_777
timestamp 1679581782
transform 1 0 146208 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_784
timestamp 1679581782
transform 1 0 146880 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_791
timestamp 1679581782
transform 1 0 147552 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_798
timestamp 1679581782
transform 1 0 148224 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_805
timestamp 1679581782
transform 1 0 148896 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_812
timestamp 1679581782
transform 1 0 149568 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_819
timestamp 1679581782
transform 1 0 150240 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_826
timestamp 1679581782
transform 1 0 150912 0 -1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_833
timestamp 1679581782
transform 1 0 151584 0 -1 142884
box -48 -56 720 834
use sg13g2_fill_1  FILLER_93_840
timestamp 1677579658
transform 1 0 152256 0 -1 142884
box -48 -56 144 834
use sg13g2_decap_8  FILLER_94_0
timestamp 1679581782
transform 1 0 71616 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_7
timestamp 1679581782
transform 1 0 72288 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_14
timestamp 1679581782
transform 1 0 72960 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_21
timestamp 1679581782
transform 1 0 73632 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_28
timestamp 1679581782
transform 1 0 74304 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_35
timestamp 1679581782
transform 1 0 74976 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_42
timestamp 1679581782
transform 1 0 75648 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_49
timestamp 1679581782
transform 1 0 76320 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_56
timestamp 1679581782
transform 1 0 76992 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_63
timestamp 1679581782
transform 1 0 77664 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_70
timestamp 1679581782
transform 1 0 78336 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_77
timestamp 1679581782
transform 1 0 79008 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_84
timestamp 1679581782
transform 1 0 79680 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_91
timestamp 1679581782
transform 1 0 80352 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_98
timestamp 1679581782
transform 1 0 81024 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_105
timestamp 1679581782
transform 1 0 81696 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_112
timestamp 1679581782
transform 1 0 82368 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_119
timestamp 1679581782
transform 1 0 83040 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_126
timestamp 1679581782
transform 1 0 83712 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_133
timestamp 1679581782
transform 1 0 84384 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_140
timestamp 1679581782
transform 1 0 85056 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_147
timestamp 1679581782
transform 1 0 85728 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_154
timestamp 1679581782
transform 1 0 86400 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_161
timestamp 1679581782
transform 1 0 87072 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_168
timestamp 1679581782
transform 1 0 87744 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_175
timestamp 1679581782
transform 1 0 88416 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_182
timestamp 1679581782
transform 1 0 89088 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_189
timestamp 1679581782
transform 1 0 89760 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_196
timestamp 1679581782
transform 1 0 90432 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_203
timestamp 1679581782
transform 1 0 91104 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_210
timestamp 1679581782
transform 1 0 91776 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_217
timestamp 1679581782
transform 1 0 92448 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_224
timestamp 1679581782
transform 1 0 93120 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_231
timestamp 1679581782
transform 1 0 93792 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_238
timestamp 1679581782
transform 1 0 94464 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_245
timestamp 1679581782
transform 1 0 95136 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_252
timestamp 1679581782
transform 1 0 95808 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_259
timestamp 1679581782
transform 1 0 96480 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_266
timestamp 1679581782
transform 1 0 97152 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_273
timestamp 1679581782
transform 1 0 97824 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_280
timestamp 1679581782
transform 1 0 98496 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_287
timestamp 1679581782
transform 1 0 99168 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_294
timestamp 1679581782
transform 1 0 99840 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_301
timestamp 1679581782
transform 1 0 100512 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_308
timestamp 1679581782
transform 1 0 101184 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_315
timestamp 1679581782
transform 1 0 101856 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_322
timestamp 1679581782
transform 1 0 102528 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_329
timestamp 1679581782
transform 1 0 103200 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_336
timestamp 1679581782
transform 1 0 103872 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_343
timestamp 1679581782
transform 1 0 104544 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_350
timestamp 1679581782
transform 1 0 105216 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_357
timestamp 1679581782
transform 1 0 105888 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_364
timestamp 1679581782
transform 1 0 106560 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_371
timestamp 1679581782
transform 1 0 107232 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_378
timestamp 1679581782
transform 1 0 107904 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_385
timestamp 1679581782
transform 1 0 108576 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_392
timestamp 1679581782
transform 1 0 109248 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_399
timestamp 1679581782
transform 1 0 109920 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_406
timestamp 1679581782
transform 1 0 110592 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_413
timestamp 1679581782
transform 1 0 111264 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_420
timestamp 1679581782
transform 1 0 111936 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_427
timestamp 1679581782
transform 1 0 112608 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_434
timestamp 1679581782
transform 1 0 113280 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_441
timestamp 1679581782
transform 1 0 113952 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_448
timestamp 1679581782
transform 1 0 114624 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_455
timestamp 1679581782
transform 1 0 115296 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_462
timestamp 1679581782
transform 1 0 115968 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_469
timestamp 1679581782
transform 1 0 116640 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_476
timestamp 1679581782
transform 1 0 117312 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_483
timestamp 1679581782
transform 1 0 117984 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_490
timestamp 1679581782
transform 1 0 118656 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_497
timestamp 1679581782
transform 1 0 119328 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_504
timestamp 1679581782
transform 1 0 120000 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_511
timestamp 1679581782
transform 1 0 120672 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_518
timestamp 1679581782
transform 1 0 121344 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_525
timestamp 1679581782
transform 1 0 122016 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_532
timestamp 1679581782
transform 1 0 122688 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_539
timestamp 1679581782
transform 1 0 123360 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_546
timestamp 1679581782
transform 1 0 124032 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_553
timestamp 1679581782
transform 1 0 124704 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_560
timestamp 1679581782
transform 1 0 125376 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_567
timestamp 1679581782
transform 1 0 126048 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_574
timestamp 1679581782
transform 1 0 126720 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_581
timestamp 1679581782
transform 1 0 127392 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_588
timestamp 1679581782
transform 1 0 128064 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_595
timestamp 1679581782
transform 1 0 128736 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_602
timestamp 1679581782
transform 1 0 129408 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_609
timestamp 1679581782
transform 1 0 130080 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_616
timestamp 1679581782
transform 1 0 130752 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_623
timestamp 1679581782
transform 1 0 131424 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_630
timestamp 1679581782
transform 1 0 132096 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_637
timestamp 1679581782
transform 1 0 132768 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_644
timestamp 1679581782
transform 1 0 133440 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_651
timestamp 1679581782
transform 1 0 134112 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_658
timestamp 1679581782
transform 1 0 134784 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_665
timestamp 1679581782
transform 1 0 135456 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_672
timestamp 1679581782
transform 1 0 136128 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_679
timestamp 1679581782
transform 1 0 136800 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_686
timestamp 1679581782
transform 1 0 137472 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_693
timestamp 1679581782
transform 1 0 138144 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_700
timestamp 1679581782
transform 1 0 138816 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_707
timestamp 1679581782
transform 1 0 139488 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_714
timestamp 1679581782
transform 1 0 140160 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_721
timestamp 1679581782
transform 1 0 140832 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_728
timestamp 1679581782
transform 1 0 141504 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_735
timestamp 1679581782
transform 1 0 142176 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_742
timestamp 1679581782
transform 1 0 142848 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_749
timestamp 1679581782
transform 1 0 143520 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_756
timestamp 1679581782
transform 1 0 144192 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_763
timestamp 1679581782
transform 1 0 144864 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_770
timestamp 1679581782
transform 1 0 145536 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_777
timestamp 1679581782
transform 1 0 146208 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_784
timestamp 1679581782
transform 1 0 146880 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_791
timestamp 1679581782
transform 1 0 147552 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_798
timestamp 1679581782
transform 1 0 148224 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_805
timestamp 1679581782
transform 1 0 148896 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_812
timestamp 1679581782
transform 1 0 149568 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_819
timestamp 1679581782
transform 1 0 150240 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_826
timestamp 1679581782
transform 1 0 150912 0 1 142884
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_833
timestamp 1679581782
transform 1 0 151584 0 1 142884
box -48 -56 720 834
use sg13g2_fill_1  FILLER_94_840
timestamp 1677579658
transform 1 0 152256 0 1 142884
box -48 -56 144 834
use sg13g2_decap_8  FILLER_95_0
timestamp 1679581782
transform 1 0 71616 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_7
timestamp 1679581782
transform 1 0 72288 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_14
timestamp 1679581782
transform 1 0 72960 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_21
timestamp 1679581782
transform 1 0 73632 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_28
timestamp 1679581782
transform 1 0 74304 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_35
timestamp 1679581782
transform 1 0 74976 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_42
timestamp 1679581782
transform 1 0 75648 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_49
timestamp 1679581782
transform 1 0 76320 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_56
timestamp 1679581782
transform 1 0 76992 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_63
timestamp 1679581782
transform 1 0 77664 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_70
timestamp 1679581782
transform 1 0 78336 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_77
timestamp 1679581782
transform 1 0 79008 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_84
timestamp 1679581782
transform 1 0 79680 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_91
timestamp 1679581782
transform 1 0 80352 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_98
timestamp 1679581782
transform 1 0 81024 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_105
timestamp 1679581782
transform 1 0 81696 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_112
timestamp 1679581782
transform 1 0 82368 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_119
timestamp 1679581782
transform 1 0 83040 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_126
timestamp 1679581782
transform 1 0 83712 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_133
timestamp 1679581782
transform 1 0 84384 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_140
timestamp 1679581782
transform 1 0 85056 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_147
timestamp 1679581782
transform 1 0 85728 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_154
timestamp 1679581782
transform 1 0 86400 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_161
timestamp 1679581782
transform 1 0 87072 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_168
timestamp 1679581782
transform 1 0 87744 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_175
timestamp 1679581782
transform 1 0 88416 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_182
timestamp 1679581782
transform 1 0 89088 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_189
timestamp 1679581782
transform 1 0 89760 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_196
timestamp 1679581782
transform 1 0 90432 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_203
timestamp 1679581782
transform 1 0 91104 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_210
timestamp 1679581782
transform 1 0 91776 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_217
timestamp 1679581782
transform 1 0 92448 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_224
timestamp 1679581782
transform 1 0 93120 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_231
timestamp 1679581782
transform 1 0 93792 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_238
timestamp 1679581782
transform 1 0 94464 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_245
timestamp 1679581782
transform 1 0 95136 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_252
timestamp 1679581782
transform 1 0 95808 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_259
timestamp 1679581782
transform 1 0 96480 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_266
timestamp 1679581782
transform 1 0 97152 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_273
timestamp 1679581782
transform 1 0 97824 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_280
timestamp 1679581782
transform 1 0 98496 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_287
timestamp 1679581782
transform 1 0 99168 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_294
timestamp 1679581782
transform 1 0 99840 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_301
timestamp 1679581782
transform 1 0 100512 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_308
timestamp 1679581782
transform 1 0 101184 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_315
timestamp 1679581782
transform 1 0 101856 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_322
timestamp 1679581782
transform 1 0 102528 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_329
timestamp 1679581782
transform 1 0 103200 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_336
timestamp 1679581782
transform 1 0 103872 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_343
timestamp 1679581782
transform 1 0 104544 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_350
timestamp 1679581782
transform 1 0 105216 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_357
timestamp 1679581782
transform 1 0 105888 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_364
timestamp 1679581782
transform 1 0 106560 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_371
timestamp 1679581782
transform 1 0 107232 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_378
timestamp 1679581782
transform 1 0 107904 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_385
timestamp 1679581782
transform 1 0 108576 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_392
timestamp 1679581782
transform 1 0 109248 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_399
timestamp 1679581782
transform 1 0 109920 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_406
timestamp 1679581782
transform 1 0 110592 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_413
timestamp 1679581782
transform 1 0 111264 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_420
timestamp 1679581782
transform 1 0 111936 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_427
timestamp 1679581782
transform 1 0 112608 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_434
timestamp 1679581782
transform 1 0 113280 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_441
timestamp 1679581782
transform 1 0 113952 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_448
timestamp 1679581782
transform 1 0 114624 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_455
timestamp 1679581782
transform 1 0 115296 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_462
timestamp 1679581782
transform 1 0 115968 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_469
timestamp 1679581782
transform 1 0 116640 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_476
timestamp 1679581782
transform 1 0 117312 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_483
timestamp 1679581782
transform 1 0 117984 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_490
timestamp 1679581782
transform 1 0 118656 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_497
timestamp 1679581782
transform 1 0 119328 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_504
timestamp 1679581782
transform 1 0 120000 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_511
timestamp 1679581782
transform 1 0 120672 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_518
timestamp 1679581782
transform 1 0 121344 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_525
timestamp 1679581782
transform 1 0 122016 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_532
timestamp 1679581782
transform 1 0 122688 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_539
timestamp 1679581782
transform 1 0 123360 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_546
timestamp 1679581782
transform 1 0 124032 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_553
timestamp 1679581782
transform 1 0 124704 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_560
timestamp 1679581782
transform 1 0 125376 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_567
timestamp 1679581782
transform 1 0 126048 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_574
timestamp 1679581782
transform 1 0 126720 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_581
timestamp 1679581782
transform 1 0 127392 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_588
timestamp 1679581782
transform 1 0 128064 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_595
timestamp 1679581782
transform 1 0 128736 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_602
timestamp 1679581782
transform 1 0 129408 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_609
timestamp 1679581782
transform 1 0 130080 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_616
timestamp 1679581782
transform 1 0 130752 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_623
timestamp 1679581782
transform 1 0 131424 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_630
timestamp 1679581782
transform 1 0 132096 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_637
timestamp 1679581782
transform 1 0 132768 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_644
timestamp 1679581782
transform 1 0 133440 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_651
timestamp 1679581782
transform 1 0 134112 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_658
timestamp 1679581782
transform 1 0 134784 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_665
timestamp 1679581782
transform 1 0 135456 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_672
timestamp 1679581782
transform 1 0 136128 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_679
timestamp 1679581782
transform 1 0 136800 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_686
timestamp 1679581782
transform 1 0 137472 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_693
timestamp 1679581782
transform 1 0 138144 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_700
timestamp 1679581782
transform 1 0 138816 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_707
timestamp 1679581782
transform 1 0 139488 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_714
timestamp 1679581782
transform 1 0 140160 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_721
timestamp 1679581782
transform 1 0 140832 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_728
timestamp 1679581782
transform 1 0 141504 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_735
timestamp 1679581782
transform 1 0 142176 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_742
timestamp 1679581782
transform 1 0 142848 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_749
timestamp 1679581782
transform 1 0 143520 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_756
timestamp 1679581782
transform 1 0 144192 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_763
timestamp 1679581782
transform 1 0 144864 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_770
timestamp 1679581782
transform 1 0 145536 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_777
timestamp 1679581782
transform 1 0 146208 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_784
timestamp 1679581782
transform 1 0 146880 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_791
timestamp 1679581782
transform 1 0 147552 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_798
timestamp 1679581782
transform 1 0 148224 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_805
timestamp 1679581782
transform 1 0 148896 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_812
timestamp 1679581782
transform 1 0 149568 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_819
timestamp 1679581782
transform 1 0 150240 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_826
timestamp 1679581782
transform 1 0 150912 0 -1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_833
timestamp 1679581782
transform 1 0 151584 0 -1 144396
box -48 -56 720 834
use sg13g2_fill_1  FILLER_95_840
timestamp 1677579658
transform 1 0 152256 0 -1 144396
box -48 -56 144 834
use sg13g2_decap_8  FILLER_96_0
timestamp 1679581782
transform 1 0 71616 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_7
timestamp 1679581782
transform 1 0 72288 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_14
timestamp 1679581782
transform 1 0 72960 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_21
timestamp 1679581782
transform 1 0 73632 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_28
timestamp 1679581782
transform 1 0 74304 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_35
timestamp 1679581782
transform 1 0 74976 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_42
timestamp 1679581782
transform 1 0 75648 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_49
timestamp 1679581782
transform 1 0 76320 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_56
timestamp 1679581782
transform 1 0 76992 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_63
timestamp 1679581782
transform 1 0 77664 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_70
timestamp 1679581782
transform 1 0 78336 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_77
timestamp 1679581782
transform 1 0 79008 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_84
timestamp 1679581782
transform 1 0 79680 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_91
timestamp 1679581782
transform 1 0 80352 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_98
timestamp 1679581782
transform 1 0 81024 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_105
timestamp 1679581782
transform 1 0 81696 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_112
timestamp 1679581782
transform 1 0 82368 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_119
timestamp 1679581782
transform 1 0 83040 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_126
timestamp 1679581782
transform 1 0 83712 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_133
timestamp 1679581782
transform 1 0 84384 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_140
timestamp 1679581782
transform 1 0 85056 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_147
timestamp 1679581782
transform 1 0 85728 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_154
timestamp 1679581782
transform 1 0 86400 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_161
timestamp 1679581782
transform 1 0 87072 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_168
timestamp 1679581782
transform 1 0 87744 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_175
timestamp 1679581782
transform 1 0 88416 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_182
timestamp 1679581782
transform 1 0 89088 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_189
timestamp 1679581782
transform 1 0 89760 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_196
timestamp 1679581782
transform 1 0 90432 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_203
timestamp 1679581782
transform 1 0 91104 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_210
timestamp 1679581782
transform 1 0 91776 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_217
timestamp 1679581782
transform 1 0 92448 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_224
timestamp 1679581782
transform 1 0 93120 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_231
timestamp 1679581782
transform 1 0 93792 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_238
timestamp 1679581782
transform 1 0 94464 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_245
timestamp 1679581782
transform 1 0 95136 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_252
timestamp 1679581782
transform 1 0 95808 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_259
timestamp 1679581782
transform 1 0 96480 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_266
timestamp 1679581782
transform 1 0 97152 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_273
timestamp 1679581782
transform 1 0 97824 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_280
timestamp 1679581782
transform 1 0 98496 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_287
timestamp 1679581782
transform 1 0 99168 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_294
timestamp 1679581782
transform 1 0 99840 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_301
timestamp 1679581782
transform 1 0 100512 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_308
timestamp 1679581782
transform 1 0 101184 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_315
timestamp 1679581782
transform 1 0 101856 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_322
timestamp 1679581782
transform 1 0 102528 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_329
timestamp 1679581782
transform 1 0 103200 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_336
timestamp 1679581782
transform 1 0 103872 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_343
timestamp 1679581782
transform 1 0 104544 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_350
timestamp 1679581782
transform 1 0 105216 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_357
timestamp 1679581782
transform 1 0 105888 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_364
timestamp 1679581782
transform 1 0 106560 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_371
timestamp 1679581782
transform 1 0 107232 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_378
timestamp 1679581782
transform 1 0 107904 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_385
timestamp 1679581782
transform 1 0 108576 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_392
timestamp 1679581782
transform 1 0 109248 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_399
timestamp 1679581782
transform 1 0 109920 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_406
timestamp 1679581782
transform 1 0 110592 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_413
timestamp 1679581782
transform 1 0 111264 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_420
timestamp 1679581782
transform 1 0 111936 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_427
timestamp 1679581782
transform 1 0 112608 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_434
timestamp 1679581782
transform 1 0 113280 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_441
timestamp 1679581782
transform 1 0 113952 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_448
timestamp 1679581782
transform 1 0 114624 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_455
timestamp 1679581782
transform 1 0 115296 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_462
timestamp 1679581782
transform 1 0 115968 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_469
timestamp 1679581782
transform 1 0 116640 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_476
timestamp 1679581782
transform 1 0 117312 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_483
timestamp 1679581782
transform 1 0 117984 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_490
timestamp 1679581782
transform 1 0 118656 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_497
timestamp 1679581782
transform 1 0 119328 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_504
timestamp 1679581782
transform 1 0 120000 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_511
timestamp 1679581782
transform 1 0 120672 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_518
timestamp 1679581782
transform 1 0 121344 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_525
timestamp 1679581782
transform 1 0 122016 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_532
timestamp 1679581782
transform 1 0 122688 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_539
timestamp 1679581782
transform 1 0 123360 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_546
timestamp 1679581782
transform 1 0 124032 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_553
timestamp 1679581782
transform 1 0 124704 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_560
timestamp 1679581782
transform 1 0 125376 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_567
timestamp 1679581782
transform 1 0 126048 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_574
timestamp 1679581782
transform 1 0 126720 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_581
timestamp 1679581782
transform 1 0 127392 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_588
timestamp 1679581782
transform 1 0 128064 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_595
timestamp 1679581782
transform 1 0 128736 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_602
timestamp 1679581782
transform 1 0 129408 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_609
timestamp 1679581782
transform 1 0 130080 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_616
timestamp 1679581782
transform 1 0 130752 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_623
timestamp 1679581782
transform 1 0 131424 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_630
timestamp 1679581782
transform 1 0 132096 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_637
timestamp 1679581782
transform 1 0 132768 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_644
timestamp 1679581782
transform 1 0 133440 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_651
timestamp 1679581782
transform 1 0 134112 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_658
timestamp 1679581782
transform 1 0 134784 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_665
timestamp 1679581782
transform 1 0 135456 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_672
timestamp 1679581782
transform 1 0 136128 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_679
timestamp 1679581782
transform 1 0 136800 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_686
timestamp 1679581782
transform 1 0 137472 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_693
timestamp 1679581782
transform 1 0 138144 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_700
timestamp 1679581782
transform 1 0 138816 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_707
timestamp 1679581782
transform 1 0 139488 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_714
timestamp 1679581782
transform 1 0 140160 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_721
timestamp 1679581782
transform 1 0 140832 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_728
timestamp 1679581782
transform 1 0 141504 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_735
timestamp 1679581782
transform 1 0 142176 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_742
timestamp 1679581782
transform 1 0 142848 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_749
timestamp 1679581782
transform 1 0 143520 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_756
timestamp 1679581782
transform 1 0 144192 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_763
timestamp 1679581782
transform 1 0 144864 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_770
timestamp 1679581782
transform 1 0 145536 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_777
timestamp 1679581782
transform 1 0 146208 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_784
timestamp 1679581782
transform 1 0 146880 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_791
timestamp 1679581782
transform 1 0 147552 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_798
timestamp 1679581782
transform 1 0 148224 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_805
timestamp 1679581782
transform 1 0 148896 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_812
timestamp 1679581782
transform 1 0 149568 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_819
timestamp 1679581782
transform 1 0 150240 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_826
timestamp 1679581782
transform 1 0 150912 0 1 144396
box -48 -56 720 834
use sg13g2_decap_8  FILLER_96_833
timestamp 1679581782
transform 1 0 151584 0 1 144396
box -48 -56 720 834
use sg13g2_fill_1  FILLER_96_840
timestamp 1677579658
transform 1 0 152256 0 1 144396
box -48 -56 144 834
use sg13g2_decap_8  FILLER_97_0
timestamp 1679581782
transform 1 0 71616 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_7
timestamp 1679581782
transform 1 0 72288 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_14
timestamp 1679581782
transform 1 0 72960 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_21
timestamp 1679581782
transform 1 0 73632 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_28
timestamp 1679581782
transform 1 0 74304 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_35
timestamp 1679581782
transform 1 0 74976 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_42
timestamp 1679581782
transform 1 0 75648 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_49
timestamp 1679581782
transform 1 0 76320 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_56
timestamp 1679581782
transform 1 0 76992 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_63
timestamp 1679581782
transform 1 0 77664 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_70
timestamp 1679581782
transform 1 0 78336 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_77
timestamp 1679581782
transform 1 0 79008 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_84
timestamp 1679581782
transform 1 0 79680 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_91
timestamp 1679581782
transform 1 0 80352 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_98
timestamp 1679581782
transform 1 0 81024 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_105
timestamp 1679581782
transform 1 0 81696 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_112
timestamp 1679581782
transform 1 0 82368 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_119
timestamp 1679581782
transform 1 0 83040 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_126
timestamp 1679581782
transform 1 0 83712 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_133
timestamp 1679581782
transform 1 0 84384 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_140
timestamp 1679581782
transform 1 0 85056 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_147
timestamp 1679581782
transform 1 0 85728 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_154
timestamp 1679581782
transform 1 0 86400 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_161
timestamp 1679581782
transform 1 0 87072 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_168
timestamp 1679581782
transform 1 0 87744 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_175
timestamp 1679581782
transform 1 0 88416 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_182
timestamp 1679581782
transform 1 0 89088 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_189
timestamp 1679581782
transform 1 0 89760 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_196
timestamp 1679581782
transform 1 0 90432 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_203
timestamp 1679581782
transform 1 0 91104 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_210
timestamp 1679581782
transform 1 0 91776 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_217
timestamp 1679581782
transform 1 0 92448 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_224
timestamp 1679581782
transform 1 0 93120 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_231
timestamp 1679581782
transform 1 0 93792 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_238
timestamp 1679581782
transform 1 0 94464 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_245
timestamp 1679581782
transform 1 0 95136 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_252
timestamp 1679581782
transform 1 0 95808 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_259
timestamp 1679581782
transform 1 0 96480 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_266
timestamp 1679581782
transform 1 0 97152 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_273
timestamp 1679581782
transform 1 0 97824 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_280
timestamp 1679581782
transform 1 0 98496 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_287
timestamp 1679581782
transform 1 0 99168 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_294
timestamp 1679581782
transform 1 0 99840 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_301
timestamp 1679581782
transform 1 0 100512 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_308
timestamp 1679581782
transform 1 0 101184 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_315
timestamp 1679581782
transform 1 0 101856 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_322
timestamp 1679581782
transform 1 0 102528 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_329
timestamp 1679581782
transform 1 0 103200 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_336
timestamp 1679581782
transform 1 0 103872 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_343
timestamp 1679581782
transform 1 0 104544 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_350
timestamp 1679581782
transform 1 0 105216 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_357
timestamp 1679581782
transform 1 0 105888 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_364
timestamp 1679581782
transform 1 0 106560 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_371
timestamp 1679581782
transform 1 0 107232 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_378
timestamp 1679581782
transform 1 0 107904 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_385
timestamp 1679581782
transform 1 0 108576 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_392
timestamp 1679581782
transform 1 0 109248 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_399
timestamp 1679581782
transform 1 0 109920 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_406
timestamp 1679581782
transform 1 0 110592 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_413
timestamp 1679581782
transform 1 0 111264 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_420
timestamp 1679581782
transform 1 0 111936 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_427
timestamp 1679581782
transform 1 0 112608 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_434
timestamp 1679581782
transform 1 0 113280 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_441
timestamp 1679581782
transform 1 0 113952 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_448
timestamp 1679581782
transform 1 0 114624 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_455
timestamp 1679581782
transform 1 0 115296 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_462
timestamp 1679581782
transform 1 0 115968 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_469
timestamp 1679581782
transform 1 0 116640 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_476
timestamp 1679581782
transform 1 0 117312 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_483
timestamp 1679581782
transform 1 0 117984 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_490
timestamp 1679581782
transform 1 0 118656 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_497
timestamp 1679581782
transform 1 0 119328 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_504
timestamp 1679581782
transform 1 0 120000 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_511
timestamp 1679581782
transform 1 0 120672 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_518
timestamp 1679581782
transform 1 0 121344 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_525
timestamp 1679581782
transform 1 0 122016 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_532
timestamp 1679581782
transform 1 0 122688 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_539
timestamp 1679581782
transform 1 0 123360 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_546
timestamp 1679581782
transform 1 0 124032 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_553
timestamp 1679581782
transform 1 0 124704 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_560
timestamp 1679581782
transform 1 0 125376 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_567
timestamp 1679581782
transform 1 0 126048 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_574
timestamp 1679581782
transform 1 0 126720 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_581
timestamp 1679581782
transform 1 0 127392 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_588
timestamp 1679581782
transform 1 0 128064 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_595
timestamp 1679581782
transform 1 0 128736 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_602
timestamp 1679581782
transform 1 0 129408 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_609
timestamp 1679581782
transform 1 0 130080 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_616
timestamp 1679581782
transform 1 0 130752 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_623
timestamp 1679581782
transform 1 0 131424 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_630
timestamp 1679581782
transform 1 0 132096 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_637
timestamp 1679581782
transform 1 0 132768 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_644
timestamp 1679581782
transform 1 0 133440 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_651
timestamp 1679581782
transform 1 0 134112 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_658
timestamp 1679581782
transform 1 0 134784 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_665
timestamp 1679581782
transform 1 0 135456 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_672
timestamp 1679581782
transform 1 0 136128 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_679
timestamp 1679581782
transform 1 0 136800 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_686
timestamp 1679581782
transform 1 0 137472 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_693
timestamp 1679581782
transform 1 0 138144 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_700
timestamp 1679581782
transform 1 0 138816 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_707
timestamp 1679581782
transform 1 0 139488 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_714
timestamp 1679581782
transform 1 0 140160 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_721
timestamp 1679581782
transform 1 0 140832 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_728
timestamp 1679581782
transform 1 0 141504 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_735
timestamp 1679581782
transform 1 0 142176 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_742
timestamp 1679581782
transform 1 0 142848 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_749
timestamp 1679581782
transform 1 0 143520 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_756
timestamp 1679581782
transform 1 0 144192 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_763
timestamp 1679581782
transform 1 0 144864 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_770
timestamp 1679581782
transform 1 0 145536 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_777
timestamp 1679581782
transform 1 0 146208 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_784
timestamp 1679581782
transform 1 0 146880 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_791
timestamp 1679581782
transform 1 0 147552 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_798
timestamp 1679581782
transform 1 0 148224 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_805
timestamp 1679581782
transform 1 0 148896 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_812
timestamp 1679581782
transform 1 0 149568 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_819
timestamp 1679581782
transform 1 0 150240 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_826
timestamp 1679581782
transform 1 0 150912 0 -1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_833
timestamp 1679581782
transform 1 0 151584 0 -1 145908
box -48 -56 720 834
use sg13g2_fill_1  FILLER_97_840
timestamp 1677579658
transform 1 0 152256 0 -1 145908
box -48 -56 144 834
use sg13g2_decap_8  FILLER_98_0
timestamp 1679581782
transform 1 0 71616 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_7
timestamp 1679581782
transform 1 0 72288 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_14
timestamp 1679581782
transform 1 0 72960 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_21
timestamp 1679581782
transform 1 0 73632 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_28
timestamp 1679581782
transform 1 0 74304 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_35
timestamp 1679581782
transform 1 0 74976 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_42
timestamp 1679581782
transform 1 0 75648 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_49
timestamp 1679581782
transform 1 0 76320 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_56
timestamp 1679581782
transform 1 0 76992 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_63
timestamp 1679581782
transform 1 0 77664 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_70
timestamp 1679581782
transform 1 0 78336 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_77
timestamp 1679581782
transform 1 0 79008 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_84
timestamp 1679581782
transform 1 0 79680 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_91
timestamp 1679581782
transform 1 0 80352 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_98
timestamp 1679581782
transform 1 0 81024 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_105
timestamp 1679581782
transform 1 0 81696 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_112
timestamp 1679581782
transform 1 0 82368 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_119
timestamp 1679581782
transform 1 0 83040 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_126
timestamp 1679581782
transform 1 0 83712 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_133
timestamp 1679581782
transform 1 0 84384 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_140
timestamp 1679581782
transform 1 0 85056 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_147
timestamp 1679581782
transform 1 0 85728 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_154
timestamp 1679581782
transform 1 0 86400 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_161
timestamp 1679581782
transform 1 0 87072 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_168
timestamp 1679581782
transform 1 0 87744 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_175
timestamp 1679581782
transform 1 0 88416 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_182
timestamp 1679581782
transform 1 0 89088 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_189
timestamp 1679581782
transform 1 0 89760 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_196
timestamp 1679581782
transform 1 0 90432 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_203
timestamp 1679581782
transform 1 0 91104 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_210
timestamp 1679581782
transform 1 0 91776 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_217
timestamp 1679581782
transform 1 0 92448 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_224
timestamp 1679581782
transform 1 0 93120 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_231
timestamp 1679581782
transform 1 0 93792 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_238
timestamp 1679581782
transform 1 0 94464 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_245
timestamp 1679581782
transform 1 0 95136 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_252
timestamp 1679581782
transform 1 0 95808 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_259
timestamp 1679581782
transform 1 0 96480 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_266
timestamp 1679581782
transform 1 0 97152 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_273
timestamp 1679581782
transform 1 0 97824 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_280
timestamp 1679581782
transform 1 0 98496 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_287
timestamp 1679581782
transform 1 0 99168 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_294
timestamp 1679581782
transform 1 0 99840 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_301
timestamp 1679581782
transform 1 0 100512 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_308
timestamp 1679581782
transform 1 0 101184 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_315
timestamp 1679581782
transform 1 0 101856 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_322
timestamp 1679581782
transform 1 0 102528 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_329
timestamp 1679581782
transform 1 0 103200 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_336
timestamp 1679581782
transform 1 0 103872 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_343
timestamp 1679581782
transform 1 0 104544 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_350
timestamp 1679581782
transform 1 0 105216 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_357
timestamp 1679581782
transform 1 0 105888 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_364
timestamp 1679581782
transform 1 0 106560 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_371
timestamp 1679581782
transform 1 0 107232 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_378
timestamp 1679581782
transform 1 0 107904 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_385
timestamp 1679581782
transform 1 0 108576 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_392
timestamp 1679581782
transform 1 0 109248 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_399
timestamp 1679581782
transform 1 0 109920 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_406
timestamp 1679581782
transform 1 0 110592 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_413
timestamp 1679581782
transform 1 0 111264 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_420
timestamp 1679581782
transform 1 0 111936 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_427
timestamp 1679581782
transform 1 0 112608 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_434
timestamp 1679581782
transform 1 0 113280 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_441
timestamp 1679581782
transform 1 0 113952 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_448
timestamp 1679581782
transform 1 0 114624 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_455
timestamp 1679581782
transform 1 0 115296 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_462
timestamp 1679581782
transform 1 0 115968 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_469
timestamp 1679581782
transform 1 0 116640 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_476
timestamp 1679581782
transform 1 0 117312 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_483
timestamp 1679581782
transform 1 0 117984 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_490
timestamp 1679581782
transform 1 0 118656 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_497
timestamp 1679581782
transform 1 0 119328 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_504
timestamp 1679581782
transform 1 0 120000 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_511
timestamp 1679581782
transform 1 0 120672 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_518
timestamp 1679581782
transform 1 0 121344 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_525
timestamp 1679581782
transform 1 0 122016 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_532
timestamp 1679581782
transform 1 0 122688 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_539
timestamp 1679581782
transform 1 0 123360 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_546
timestamp 1679581782
transform 1 0 124032 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_553
timestamp 1679581782
transform 1 0 124704 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_560
timestamp 1679581782
transform 1 0 125376 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_567
timestamp 1679581782
transform 1 0 126048 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_574
timestamp 1679581782
transform 1 0 126720 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_581
timestamp 1679581782
transform 1 0 127392 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_588
timestamp 1679581782
transform 1 0 128064 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_595
timestamp 1679581782
transform 1 0 128736 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_602
timestamp 1679581782
transform 1 0 129408 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_609
timestamp 1679581782
transform 1 0 130080 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_616
timestamp 1679581782
transform 1 0 130752 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_623
timestamp 1679581782
transform 1 0 131424 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_630
timestamp 1679581782
transform 1 0 132096 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_637
timestamp 1679581782
transform 1 0 132768 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_644
timestamp 1679581782
transform 1 0 133440 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_651
timestamp 1679581782
transform 1 0 134112 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_658
timestamp 1679581782
transform 1 0 134784 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_665
timestamp 1679581782
transform 1 0 135456 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_672
timestamp 1679581782
transform 1 0 136128 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_679
timestamp 1679581782
transform 1 0 136800 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_686
timestamp 1679581782
transform 1 0 137472 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_693
timestamp 1679581782
transform 1 0 138144 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_700
timestamp 1679581782
transform 1 0 138816 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_707
timestamp 1679581782
transform 1 0 139488 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_714
timestamp 1679581782
transform 1 0 140160 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_721
timestamp 1679581782
transform 1 0 140832 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_728
timestamp 1679581782
transform 1 0 141504 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_735
timestamp 1679581782
transform 1 0 142176 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_742
timestamp 1679581782
transform 1 0 142848 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_749
timestamp 1679581782
transform 1 0 143520 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_756
timestamp 1679581782
transform 1 0 144192 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_763
timestamp 1679581782
transform 1 0 144864 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_770
timestamp 1679581782
transform 1 0 145536 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_777
timestamp 1679581782
transform 1 0 146208 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_784
timestamp 1679581782
transform 1 0 146880 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_791
timestamp 1679581782
transform 1 0 147552 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_798
timestamp 1679581782
transform 1 0 148224 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_805
timestamp 1679581782
transform 1 0 148896 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_812
timestamp 1679581782
transform 1 0 149568 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_819
timestamp 1679581782
transform 1 0 150240 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_826
timestamp 1679581782
transform 1 0 150912 0 1 145908
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_833
timestamp 1679581782
transform 1 0 151584 0 1 145908
box -48 -56 720 834
use sg13g2_fill_1  FILLER_98_840
timestamp 1677579658
transform 1 0 152256 0 1 145908
box -48 -56 144 834
use sg13g2_decap_8  FILLER_99_0
timestamp 1679581782
transform 1 0 71616 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_7
timestamp 1679581782
transform 1 0 72288 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_14
timestamp 1679581782
transform 1 0 72960 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_21
timestamp 1679581782
transform 1 0 73632 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_28
timestamp 1679581782
transform 1 0 74304 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_35
timestamp 1679581782
transform 1 0 74976 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_42
timestamp 1679581782
transform 1 0 75648 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_49
timestamp 1679581782
transform 1 0 76320 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_56
timestamp 1679581782
transform 1 0 76992 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_63
timestamp 1679581782
transform 1 0 77664 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_70
timestamp 1679581782
transform 1 0 78336 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_77
timestamp 1679581782
transform 1 0 79008 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_84
timestamp 1679581782
transform 1 0 79680 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_91
timestamp 1679581782
transform 1 0 80352 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_98
timestamp 1679581782
transform 1 0 81024 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_105
timestamp 1679581782
transform 1 0 81696 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_112
timestamp 1679581782
transform 1 0 82368 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_119
timestamp 1679581782
transform 1 0 83040 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_126
timestamp 1679581782
transform 1 0 83712 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_133
timestamp 1679581782
transform 1 0 84384 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_140
timestamp 1679581782
transform 1 0 85056 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_147
timestamp 1679581782
transform 1 0 85728 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_154
timestamp 1679581782
transform 1 0 86400 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_161
timestamp 1679581782
transform 1 0 87072 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_168
timestamp 1679581782
transform 1 0 87744 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_175
timestamp 1679581782
transform 1 0 88416 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_182
timestamp 1679581782
transform 1 0 89088 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_189
timestamp 1679581782
transform 1 0 89760 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_196
timestamp 1679581782
transform 1 0 90432 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_203
timestamp 1679581782
transform 1 0 91104 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_210
timestamp 1679581782
transform 1 0 91776 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_217
timestamp 1679581782
transform 1 0 92448 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_224
timestamp 1679581782
transform 1 0 93120 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_231
timestamp 1679581782
transform 1 0 93792 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_238
timestamp 1679581782
transform 1 0 94464 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_245
timestamp 1679581782
transform 1 0 95136 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_252
timestamp 1679581782
transform 1 0 95808 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_259
timestamp 1679581782
transform 1 0 96480 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_266
timestamp 1679581782
transform 1 0 97152 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_273
timestamp 1679581782
transform 1 0 97824 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_280
timestamp 1679581782
transform 1 0 98496 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_287
timestamp 1679581782
transform 1 0 99168 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_294
timestamp 1679581782
transform 1 0 99840 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_301
timestamp 1679581782
transform 1 0 100512 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_308
timestamp 1679581782
transform 1 0 101184 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_315
timestamp 1679581782
transform 1 0 101856 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_322
timestamp 1679581782
transform 1 0 102528 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_329
timestamp 1679581782
transform 1 0 103200 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_336
timestamp 1679581782
transform 1 0 103872 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_343
timestamp 1679581782
transform 1 0 104544 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_350
timestamp 1679581782
transform 1 0 105216 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_357
timestamp 1679581782
transform 1 0 105888 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_364
timestamp 1679581782
transform 1 0 106560 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_371
timestamp 1679581782
transform 1 0 107232 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_378
timestamp 1679581782
transform 1 0 107904 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_385
timestamp 1679581782
transform 1 0 108576 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_392
timestamp 1679581782
transform 1 0 109248 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_399
timestamp 1679581782
transform 1 0 109920 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_406
timestamp 1679581782
transform 1 0 110592 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_413
timestamp 1679581782
transform 1 0 111264 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_420
timestamp 1679581782
transform 1 0 111936 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_427
timestamp 1679581782
transform 1 0 112608 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_434
timestamp 1679581782
transform 1 0 113280 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_441
timestamp 1679581782
transform 1 0 113952 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_448
timestamp 1679581782
transform 1 0 114624 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_455
timestamp 1679581782
transform 1 0 115296 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_462
timestamp 1679581782
transform 1 0 115968 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_469
timestamp 1679581782
transform 1 0 116640 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_476
timestamp 1679581782
transform 1 0 117312 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_483
timestamp 1679581782
transform 1 0 117984 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_490
timestamp 1679581782
transform 1 0 118656 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_497
timestamp 1679581782
transform 1 0 119328 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_504
timestamp 1679581782
transform 1 0 120000 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_511
timestamp 1679581782
transform 1 0 120672 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_518
timestamp 1679581782
transform 1 0 121344 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_525
timestamp 1679581782
transform 1 0 122016 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_532
timestamp 1679581782
transform 1 0 122688 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_539
timestamp 1679581782
transform 1 0 123360 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_546
timestamp 1679581782
transform 1 0 124032 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_553
timestamp 1679581782
transform 1 0 124704 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_560
timestamp 1679581782
transform 1 0 125376 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_567
timestamp 1679581782
transform 1 0 126048 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_574
timestamp 1679581782
transform 1 0 126720 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_581
timestamp 1679581782
transform 1 0 127392 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_588
timestamp 1679581782
transform 1 0 128064 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_595
timestamp 1679581782
transform 1 0 128736 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_602
timestamp 1679581782
transform 1 0 129408 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_609
timestamp 1679581782
transform 1 0 130080 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_616
timestamp 1679581782
transform 1 0 130752 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_623
timestamp 1679581782
transform 1 0 131424 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_630
timestamp 1679581782
transform 1 0 132096 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_637
timestamp 1679581782
transform 1 0 132768 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_644
timestamp 1679581782
transform 1 0 133440 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_651
timestamp 1679581782
transform 1 0 134112 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_658
timestamp 1679581782
transform 1 0 134784 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_665
timestamp 1679581782
transform 1 0 135456 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_672
timestamp 1679581782
transform 1 0 136128 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_679
timestamp 1679581782
transform 1 0 136800 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_686
timestamp 1679581782
transform 1 0 137472 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_693
timestamp 1679581782
transform 1 0 138144 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_700
timestamp 1679581782
transform 1 0 138816 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_707
timestamp 1679581782
transform 1 0 139488 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_714
timestamp 1679581782
transform 1 0 140160 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_721
timestamp 1679581782
transform 1 0 140832 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_728
timestamp 1679581782
transform 1 0 141504 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_735
timestamp 1679581782
transform 1 0 142176 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_742
timestamp 1679581782
transform 1 0 142848 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_749
timestamp 1679581782
transform 1 0 143520 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_756
timestamp 1679581782
transform 1 0 144192 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_763
timestamp 1679581782
transform 1 0 144864 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_770
timestamp 1679581782
transform 1 0 145536 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_777
timestamp 1679581782
transform 1 0 146208 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_784
timestamp 1679581782
transform 1 0 146880 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_791
timestamp 1679581782
transform 1 0 147552 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_798
timestamp 1679581782
transform 1 0 148224 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_805
timestamp 1679581782
transform 1 0 148896 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_812
timestamp 1679581782
transform 1 0 149568 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_819
timestamp 1679581782
transform 1 0 150240 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_826
timestamp 1679581782
transform 1 0 150912 0 -1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_833
timestamp 1679581782
transform 1 0 151584 0 -1 147420
box -48 -56 720 834
use sg13g2_fill_1  FILLER_99_840
timestamp 1677579658
transform 1 0 152256 0 -1 147420
box -48 -56 144 834
use sg13g2_decap_8  FILLER_100_0
timestamp 1679581782
transform 1 0 71616 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_7
timestamp 1679581782
transform 1 0 72288 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_14
timestamp 1679581782
transform 1 0 72960 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_21
timestamp 1679581782
transform 1 0 73632 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_28
timestamp 1679581782
transform 1 0 74304 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_35
timestamp 1679581782
transform 1 0 74976 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_42
timestamp 1679581782
transform 1 0 75648 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_49
timestamp 1679581782
transform 1 0 76320 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_56
timestamp 1679581782
transform 1 0 76992 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_63
timestamp 1679581782
transform 1 0 77664 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_70
timestamp 1679581782
transform 1 0 78336 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_77
timestamp 1679581782
transform 1 0 79008 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_84
timestamp 1679581782
transform 1 0 79680 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_91
timestamp 1679581782
transform 1 0 80352 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_98
timestamp 1679581782
transform 1 0 81024 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_105
timestamp 1679581782
transform 1 0 81696 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_112
timestamp 1679581782
transform 1 0 82368 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_119
timestamp 1679581782
transform 1 0 83040 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_126
timestamp 1679581782
transform 1 0 83712 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_133
timestamp 1679581782
transform 1 0 84384 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_140
timestamp 1679581782
transform 1 0 85056 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_147
timestamp 1679581782
transform 1 0 85728 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_154
timestamp 1679581782
transform 1 0 86400 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_161
timestamp 1679581782
transform 1 0 87072 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_168
timestamp 1679581782
transform 1 0 87744 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_175
timestamp 1679581782
transform 1 0 88416 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_182
timestamp 1679581782
transform 1 0 89088 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_189
timestamp 1679581782
transform 1 0 89760 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_196
timestamp 1679581782
transform 1 0 90432 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_203
timestamp 1679581782
transform 1 0 91104 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_210
timestamp 1679581782
transform 1 0 91776 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_217
timestamp 1679581782
transform 1 0 92448 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_224
timestamp 1679581782
transform 1 0 93120 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_231
timestamp 1679581782
transform 1 0 93792 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_238
timestamp 1679581782
transform 1 0 94464 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_245
timestamp 1679581782
transform 1 0 95136 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_252
timestamp 1679581782
transform 1 0 95808 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_259
timestamp 1679581782
transform 1 0 96480 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_266
timestamp 1679581782
transform 1 0 97152 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_273
timestamp 1679581782
transform 1 0 97824 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_280
timestamp 1679581782
transform 1 0 98496 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_287
timestamp 1679581782
transform 1 0 99168 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_294
timestamp 1679581782
transform 1 0 99840 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_301
timestamp 1679581782
transform 1 0 100512 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_308
timestamp 1679581782
transform 1 0 101184 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_315
timestamp 1679581782
transform 1 0 101856 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_322
timestamp 1679581782
transform 1 0 102528 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_329
timestamp 1679581782
transform 1 0 103200 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_336
timestamp 1679581782
transform 1 0 103872 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_343
timestamp 1679581782
transform 1 0 104544 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_350
timestamp 1679581782
transform 1 0 105216 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_357
timestamp 1679581782
transform 1 0 105888 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_364
timestamp 1679581782
transform 1 0 106560 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_371
timestamp 1679581782
transform 1 0 107232 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_378
timestamp 1679581782
transform 1 0 107904 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_385
timestamp 1679581782
transform 1 0 108576 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_392
timestamp 1679581782
transform 1 0 109248 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_399
timestamp 1679581782
transform 1 0 109920 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_406
timestamp 1679581782
transform 1 0 110592 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_413
timestamp 1679581782
transform 1 0 111264 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_420
timestamp 1679581782
transform 1 0 111936 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_427
timestamp 1679581782
transform 1 0 112608 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_434
timestamp 1679581782
transform 1 0 113280 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_441
timestamp 1679581782
transform 1 0 113952 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_448
timestamp 1679581782
transform 1 0 114624 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_455
timestamp 1679581782
transform 1 0 115296 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_462
timestamp 1679581782
transform 1 0 115968 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_469
timestamp 1679581782
transform 1 0 116640 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_476
timestamp 1679581782
transform 1 0 117312 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_483
timestamp 1679581782
transform 1 0 117984 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_490
timestamp 1679581782
transform 1 0 118656 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_497
timestamp 1679581782
transform 1 0 119328 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_504
timestamp 1679581782
transform 1 0 120000 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_511
timestamp 1679581782
transform 1 0 120672 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_518
timestamp 1679581782
transform 1 0 121344 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_525
timestamp 1679581782
transform 1 0 122016 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_532
timestamp 1679581782
transform 1 0 122688 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_539
timestamp 1679581782
transform 1 0 123360 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_546
timestamp 1679581782
transform 1 0 124032 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_553
timestamp 1679581782
transform 1 0 124704 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_560
timestamp 1679581782
transform 1 0 125376 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_567
timestamp 1679581782
transform 1 0 126048 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_574
timestamp 1679581782
transform 1 0 126720 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_581
timestamp 1679581782
transform 1 0 127392 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_588
timestamp 1679581782
transform 1 0 128064 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_595
timestamp 1679581782
transform 1 0 128736 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_602
timestamp 1679581782
transform 1 0 129408 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_609
timestamp 1679581782
transform 1 0 130080 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_616
timestamp 1679581782
transform 1 0 130752 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_623
timestamp 1679581782
transform 1 0 131424 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_630
timestamp 1679581782
transform 1 0 132096 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_637
timestamp 1679581782
transform 1 0 132768 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_644
timestamp 1679581782
transform 1 0 133440 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_651
timestamp 1679581782
transform 1 0 134112 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_658
timestamp 1679581782
transform 1 0 134784 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_665
timestamp 1679581782
transform 1 0 135456 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_672
timestamp 1679581782
transform 1 0 136128 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_679
timestamp 1679581782
transform 1 0 136800 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_686
timestamp 1679581782
transform 1 0 137472 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_693
timestamp 1679581782
transform 1 0 138144 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_700
timestamp 1679581782
transform 1 0 138816 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_707
timestamp 1679581782
transform 1 0 139488 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_714
timestamp 1679581782
transform 1 0 140160 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_721
timestamp 1679581782
transform 1 0 140832 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_728
timestamp 1679581782
transform 1 0 141504 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_735
timestamp 1679581782
transform 1 0 142176 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_742
timestamp 1679581782
transform 1 0 142848 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_749
timestamp 1679581782
transform 1 0 143520 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_756
timestamp 1679581782
transform 1 0 144192 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_763
timestamp 1679581782
transform 1 0 144864 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_770
timestamp 1679581782
transform 1 0 145536 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_777
timestamp 1679581782
transform 1 0 146208 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_784
timestamp 1679581782
transform 1 0 146880 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_791
timestamp 1679581782
transform 1 0 147552 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_798
timestamp 1679581782
transform 1 0 148224 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_805
timestamp 1679581782
transform 1 0 148896 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_812
timestamp 1679581782
transform 1 0 149568 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_819
timestamp 1679581782
transform 1 0 150240 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_826
timestamp 1679581782
transform 1 0 150912 0 1 147420
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_833
timestamp 1679581782
transform 1 0 151584 0 1 147420
box -48 -56 720 834
use sg13g2_fill_1  FILLER_100_840
timestamp 1677579658
transform 1 0 152256 0 1 147420
box -48 -56 144 834
use sg13g2_decap_8  FILLER_101_0
timestamp 1679581782
transform 1 0 71616 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_7
timestamp 1679581782
transform 1 0 72288 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_14
timestamp 1679581782
transform 1 0 72960 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_21
timestamp 1679581782
transform 1 0 73632 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_28
timestamp 1679581782
transform 1 0 74304 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_35
timestamp 1679581782
transform 1 0 74976 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_42
timestamp 1679581782
transform 1 0 75648 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_49
timestamp 1679581782
transform 1 0 76320 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_56
timestamp 1679581782
transform 1 0 76992 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_63
timestamp 1679581782
transform 1 0 77664 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_70
timestamp 1679581782
transform 1 0 78336 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_77
timestamp 1679581782
transform 1 0 79008 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_84
timestamp 1679581782
transform 1 0 79680 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_91
timestamp 1679581782
transform 1 0 80352 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_98
timestamp 1679581782
transform 1 0 81024 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_105
timestamp 1679581782
transform 1 0 81696 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_112
timestamp 1679581782
transform 1 0 82368 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_119
timestamp 1679581782
transform 1 0 83040 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_126
timestamp 1679581782
transform 1 0 83712 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_133
timestamp 1679581782
transform 1 0 84384 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_140
timestamp 1679581782
transform 1 0 85056 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_147
timestamp 1679581782
transform 1 0 85728 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_154
timestamp 1679581782
transform 1 0 86400 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_161
timestamp 1679581782
transform 1 0 87072 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_168
timestamp 1679581782
transform 1 0 87744 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_175
timestamp 1679581782
transform 1 0 88416 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_182
timestamp 1679581782
transform 1 0 89088 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_189
timestamp 1679581782
transform 1 0 89760 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_196
timestamp 1679581782
transform 1 0 90432 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_203
timestamp 1679581782
transform 1 0 91104 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_210
timestamp 1679581782
transform 1 0 91776 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_217
timestamp 1679581782
transform 1 0 92448 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_224
timestamp 1679581782
transform 1 0 93120 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_231
timestamp 1679581782
transform 1 0 93792 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_238
timestamp 1679581782
transform 1 0 94464 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_245
timestamp 1679581782
transform 1 0 95136 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_252
timestamp 1679581782
transform 1 0 95808 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_259
timestamp 1679581782
transform 1 0 96480 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_266
timestamp 1679581782
transform 1 0 97152 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_273
timestamp 1679581782
transform 1 0 97824 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_280
timestamp 1679581782
transform 1 0 98496 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_287
timestamp 1679581782
transform 1 0 99168 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_294
timestamp 1679581782
transform 1 0 99840 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_301
timestamp 1679581782
transform 1 0 100512 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_308
timestamp 1679581782
transform 1 0 101184 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_315
timestamp 1679581782
transform 1 0 101856 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_322
timestamp 1679581782
transform 1 0 102528 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_329
timestamp 1679581782
transform 1 0 103200 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_336
timestamp 1679581782
transform 1 0 103872 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_343
timestamp 1679581782
transform 1 0 104544 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_350
timestamp 1679581782
transform 1 0 105216 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_357
timestamp 1679581782
transform 1 0 105888 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_364
timestamp 1679581782
transform 1 0 106560 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_371
timestamp 1679581782
transform 1 0 107232 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_378
timestamp 1679581782
transform 1 0 107904 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_385
timestamp 1679581782
transform 1 0 108576 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_392
timestamp 1679581782
transform 1 0 109248 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_399
timestamp 1679581782
transform 1 0 109920 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_406
timestamp 1679581782
transform 1 0 110592 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_413
timestamp 1679581782
transform 1 0 111264 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_420
timestamp 1679581782
transform 1 0 111936 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_427
timestamp 1679581782
transform 1 0 112608 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_434
timestamp 1679581782
transform 1 0 113280 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_441
timestamp 1679581782
transform 1 0 113952 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_448
timestamp 1679581782
transform 1 0 114624 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_455
timestamp 1679581782
transform 1 0 115296 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_462
timestamp 1679581782
transform 1 0 115968 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_469
timestamp 1679581782
transform 1 0 116640 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_476
timestamp 1679581782
transform 1 0 117312 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_483
timestamp 1679581782
transform 1 0 117984 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_490
timestamp 1679581782
transform 1 0 118656 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_497
timestamp 1679581782
transform 1 0 119328 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_504
timestamp 1679581782
transform 1 0 120000 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_511
timestamp 1679581782
transform 1 0 120672 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_518
timestamp 1679581782
transform 1 0 121344 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_525
timestamp 1679581782
transform 1 0 122016 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_532
timestamp 1679581782
transform 1 0 122688 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_539
timestamp 1679581782
transform 1 0 123360 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_546
timestamp 1679581782
transform 1 0 124032 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_553
timestamp 1679581782
transform 1 0 124704 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_560
timestamp 1679581782
transform 1 0 125376 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_567
timestamp 1679581782
transform 1 0 126048 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_574
timestamp 1679581782
transform 1 0 126720 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_581
timestamp 1679581782
transform 1 0 127392 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_588
timestamp 1679581782
transform 1 0 128064 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_595
timestamp 1679581782
transform 1 0 128736 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_602
timestamp 1679581782
transform 1 0 129408 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_609
timestamp 1679581782
transform 1 0 130080 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_616
timestamp 1679581782
transform 1 0 130752 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_623
timestamp 1679581782
transform 1 0 131424 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_630
timestamp 1679581782
transform 1 0 132096 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_637
timestamp 1679581782
transform 1 0 132768 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_644
timestamp 1679581782
transform 1 0 133440 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_651
timestamp 1679581782
transform 1 0 134112 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_658
timestamp 1679581782
transform 1 0 134784 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_665
timestamp 1679581782
transform 1 0 135456 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_672
timestamp 1679581782
transform 1 0 136128 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_679
timestamp 1679581782
transform 1 0 136800 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_686
timestamp 1679581782
transform 1 0 137472 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_693
timestamp 1679581782
transform 1 0 138144 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_700
timestamp 1679581782
transform 1 0 138816 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_707
timestamp 1679581782
transform 1 0 139488 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_714
timestamp 1679581782
transform 1 0 140160 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_721
timestamp 1679581782
transform 1 0 140832 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_728
timestamp 1679581782
transform 1 0 141504 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_735
timestamp 1679581782
transform 1 0 142176 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_742
timestamp 1679581782
transform 1 0 142848 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_749
timestamp 1679581782
transform 1 0 143520 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_756
timestamp 1679581782
transform 1 0 144192 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_763
timestamp 1679581782
transform 1 0 144864 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_770
timestamp 1679581782
transform 1 0 145536 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_777
timestamp 1679581782
transform 1 0 146208 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_784
timestamp 1679581782
transform 1 0 146880 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_791
timestamp 1679581782
transform 1 0 147552 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_798
timestamp 1679581782
transform 1 0 148224 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_805
timestamp 1679581782
transform 1 0 148896 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_812
timestamp 1679581782
transform 1 0 149568 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_819
timestamp 1679581782
transform 1 0 150240 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_826
timestamp 1679581782
transform 1 0 150912 0 -1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_101_833
timestamp 1679581782
transform 1 0 151584 0 -1 148932
box -48 -56 720 834
use sg13g2_fill_1  FILLER_101_840
timestamp 1677579658
transform 1 0 152256 0 -1 148932
box -48 -56 144 834
use sg13g2_decap_8  FILLER_102_0
timestamp 1679581782
transform 1 0 71616 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_7
timestamp 1679581782
transform 1 0 72288 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_14
timestamp 1679581782
transform 1 0 72960 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_21
timestamp 1679581782
transform 1 0 73632 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_28
timestamp 1679581782
transform 1 0 74304 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_35
timestamp 1679581782
transform 1 0 74976 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_42
timestamp 1679581782
transform 1 0 75648 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_49
timestamp 1679581782
transform 1 0 76320 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_56
timestamp 1679581782
transform 1 0 76992 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_63
timestamp 1679581782
transform 1 0 77664 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_70
timestamp 1679581782
transform 1 0 78336 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_77
timestamp 1679581782
transform 1 0 79008 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_84
timestamp 1679581782
transform 1 0 79680 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_91
timestamp 1679581782
transform 1 0 80352 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_98
timestamp 1679581782
transform 1 0 81024 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_105
timestamp 1679581782
transform 1 0 81696 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_112
timestamp 1679581782
transform 1 0 82368 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_119
timestamp 1679581782
transform 1 0 83040 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_126
timestamp 1679581782
transform 1 0 83712 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_133
timestamp 1679581782
transform 1 0 84384 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_140
timestamp 1679581782
transform 1 0 85056 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_147
timestamp 1679581782
transform 1 0 85728 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_154
timestamp 1679581782
transform 1 0 86400 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_161
timestamp 1679581782
transform 1 0 87072 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_168
timestamp 1679581782
transform 1 0 87744 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_175
timestamp 1679581782
transform 1 0 88416 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_182
timestamp 1679581782
transform 1 0 89088 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_189
timestamp 1679581782
transform 1 0 89760 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_196
timestamp 1679581782
transform 1 0 90432 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_203
timestamp 1679581782
transform 1 0 91104 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_210
timestamp 1679581782
transform 1 0 91776 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_217
timestamp 1679581782
transform 1 0 92448 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_224
timestamp 1679581782
transform 1 0 93120 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_231
timestamp 1679581782
transform 1 0 93792 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_238
timestamp 1679581782
transform 1 0 94464 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_245
timestamp 1679581782
transform 1 0 95136 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_252
timestamp 1679581782
transform 1 0 95808 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_259
timestamp 1679581782
transform 1 0 96480 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_266
timestamp 1679581782
transform 1 0 97152 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_273
timestamp 1679581782
transform 1 0 97824 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_280
timestamp 1679581782
transform 1 0 98496 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_287
timestamp 1679581782
transform 1 0 99168 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_294
timestamp 1679581782
transform 1 0 99840 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_301
timestamp 1679581782
transform 1 0 100512 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_308
timestamp 1679581782
transform 1 0 101184 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_315
timestamp 1679581782
transform 1 0 101856 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_322
timestamp 1679581782
transform 1 0 102528 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_329
timestamp 1679581782
transform 1 0 103200 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_336
timestamp 1679581782
transform 1 0 103872 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_343
timestamp 1679581782
transform 1 0 104544 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_350
timestamp 1679581782
transform 1 0 105216 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_357
timestamp 1679581782
transform 1 0 105888 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_364
timestamp 1679581782
transform 1 0 106560 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_371
timestamp 1679581782
transform 1 0 107232 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_378
timestamp 1679581782
transform 1 0 107904 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_385
timestamp 1679581782
transform 1 0 108576 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_392
timestamp 1679581782
transform 1 0 109248 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_399
timestamp 1679581782
transform 1 0 109920 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_406
timestamp 1679581782
transform 1 0 110592 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_413
timestamp 1679581782
transform 1 0 111264 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_420
timestamp 1679581782
transform 1 0 111936 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_427
timestamp 1679581782
transform 1 0 112608 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_434
timestamp 1679581782
transform 1 0 113280 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_441
timestamp 1679581782
transform 1 0 113952 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_448
timestamp 1679581782
transform 1 0 114624 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_455
timestamp 1679581782
transform 1 0 115296 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_462
timestamp 1679581782
transform 1 0 115968 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_469
timestamp 1679581782
transform 1 0 116640 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_476
timestamp 1679581782
transform 1 0 117312 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_483
timestamp 1679581782
transform 1 0 117984 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_490
timestamp 1679581782
transform 1 0 118656 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_497
timestamp 1679581782
transform 1 0 119328 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_504
timestamp 1679581782
transform 1 0 120000 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_511
timestamp 1679581782
transform 1 0 120672 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_518
timestamp 1679581782
transform 1 0 121344 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_525
timestamp 1679581782
transform 1 0 122016 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_532
timestamp 1679581782
transform 1 0 122688 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_539
timestamp 1679581782
transform 1 0 123360 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_546
timestamp 1679581782
transform 1 0 124032 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_553
timestamp 1679581782
transform 1 0 124704 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_560
timestamp 1679581782
transform 1 0 125376 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_567
timestamp 1679581782
transform 1 0 126048 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_574
timestamp 1679581782
transform 1 0 126720 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_581
timestamp 1679581782
transform 1 0 127392 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_588
timestamp 1679581782
transform 1 0 128064 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_595
timestamp 1679581782
transform 1 0 128736 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_602
timestamp 1679581782
transform 1 0 129408 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_609
timestamp 1679581782
transform 1 0 130080 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_616
timestamp 1679581782
transform 1 0 130752 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_623
timestamp 1679581782
transform 1 0 131424 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_630
timestamp 1679581782
transform 1 0 132096 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_637
timestamp 1679581782
transform 1 0 132768 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_644
timestamp 1679581782
transform 1 0 133440 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_651
timestamp 1679581782
transform 1 0 134112 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_658
timestamp 1679581782
transform 1 0 134784 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_665
timestamp 1679581782
transform 1 0 135456 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_672
timestamp 1679581782
transform 1 0 136128 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_679
timestamp 1679581782
transform 1 0 136800 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_686
timestamp 1679581782
transform 1 0 137472 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_693
timestamp 1679581782
transform 1 0 138144 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_700
timestamp 1679581782
transform 1 0 138816 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_707
timestamp 1679581782
transform 1 0 139488 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_714
timestamp 1679581782
transform 1 0 140160 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_721
timestamp 1679581782
transform 1 0 140832 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_728
timestamp 1679581782
transform 1 0 141504 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_735
timestamp 1679581782
transform 1 0 142176 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_742
timestamp 1679581782
transform 1 0 142848 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_749
timestamp 1679581782
transform 1 0 143520 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_756
timestamp 1679581782
transform 1 0 144192 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_763
timestamp 1679581782
transform 1 0 144864 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_770
timestamp 1679581782
transform 1 0 145536 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_777
timestamp 1679581782
transform 1 0 146208 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_784
timestamp 1679581782
transform 1 0 146880 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_791
timestamp 1679581782
transform 1 0 147552 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_798
timestamp 1679581782
transform 1 0 148224 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_805
timestamp 1679581782
transform 1 0 148896 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_812
timestamp 1679581782
transform 1 0 149568 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_819
timestamp 1679581782
transform 1 0 150240 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_826
timestamp 1679581782
transform 1 0 150912 0 1 148932
box -48 -56 720 834
use sg13g2_decap_8  FILLER_102_833
timestamp 1679581782
transform 1 0 151584 0 1 148932
box -48 -56 720 834
use sg13g2_fill_1  FILLER_102_840
timestamp 1677579658
transform 1 0 152256 0 1 148932
box -48 -56 144 834
use sg13g2_decap_8  FILLER_103_0
timestamp 1679581782
transform 1 0 71616 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_7
timestamp 1679581782
transform 1 0 72288 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_14
timestamp 1679581782
transform 1 0 72960 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_21
timestamp 1679581782
transform 1 0 73632 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_28
timestamp 1679581782
transform 1 0 74304 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_35
timestamp 1679581782
transform 1 0 74976 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_42
timestamp 1679581782
transform 1 0 75648 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_49
timestamp 1679581782
transform 1 0 76320 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_56
timestamp 1679581782
transform 1 0 76992 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_63
timestamp 1679581782
transform 1 0 77664 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_70
timestamp 1679581782
transform 1 0 78336 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_77
timestamp 1679581782
transform 1 0 79008 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_84
timestamp 1679581782
transform 1 0 79680 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_91
timestamp 1679581782
transform 1 0 80352 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_98
timestamp 1679581782
transform 1 0 81024 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_105
timestamp 1679581782
transform 1 0 81696 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_112
timestamp 1679581782
transform 1 0 82368 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_119
timestamp 1679581782
transform 1 0 83040 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_126
timestamp 1679581782
transform 1 0 83712 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_133
timestamp 1679581782
transform 1 0 84384 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_140
timestamp 1679581782
transform 1 0 85056 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_147
timestamp 1679581782
transform 1 0 85728 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_154
timestamp 1679581782
transform 1 0 86400 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_161
timestamp 1679581782
transform 1 0 87072 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_168
timestamp 1679581782
transform 1 0 87744 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_175
timestamp 1679581782
transform 1 0 88416 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_182
timestamp 1679581782
transform 1 0 89088 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_189
timestamp 1679581782
transform 1 0 89760 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_196
timestamp 1679581782
transform 1 0 90432 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_203
timestamp 1679581782
transform 1 0 91104 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_210
timestamp 1679581782
transform 1 0 91776 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_217
timestamp 1679581782
transform 1 0 92448 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_224
timestamp 1679581782
transform 1 0 93120 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_231
timestamp 1679581782
transform 1 0 93792 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_238
timestamp 1679581782
transform 1 0 94464 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_245
timestamp 1679581782
transform 1 0 95136 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_252
timestamp 1679581782
transform 1 0 95808 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_259
timestamp 1679581782
transform 1 0 96480 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_266
timestamp 1679581782
transform 1 0 97152 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_273
timestamp 1679581782
transform 1 0 97824 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_280
timestamp 1679581782
transform 1 0 98496 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_287
timestamp 1679581782
transform 1 0 99168 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_294
timestamp 1679581782
transform 1 0 99840 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_301
timestamp 1679581782
transform 1 0 100512 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_308
timestamp 1679581782
transform 1 0 101184 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_315
timestamp 1679581782
transform 1 0 101856 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_322
timestamp 1679581782
transform 1 0 102528 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_329
timestamp 1679581782
transform 1 0 103200 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_336
timestamp 1679581782
transform 1 0 103872 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_343
timestamp 1679581782
transform 1 0 104544 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_350
timestamp 1679581782
transform 1 0 105216 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_357
timestamp 1679581782
transform 1 0 105888 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_364
timestamp 1679581782
transform 1 0 106560 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_371
timestamp 1679581782
transform 1 0 107232 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_378
timestamp 1679581782
transform 1 0 107904 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_385
timestamp 1679581782
transform 1 0 108576 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_392
timestamp 1679581782
transform 1 0 109248 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_399
timestamp 1679581782
transform 1 0 109920 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_406
timestamp 1679581782
transform 1 0 110592 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_413
timestamp 1679581782
transform 1 0 111264 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_420
timestamp 1679581782
transform 1 0 111936 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_427
timestamp 1679581782
transform 1 0 112608 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_434
timestamp 1679581782
transform 1 0 113280 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_441
timestamp 1679581782
transform 1 0 113952 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_448
timestamp 1679581782
transform 1 0 114624 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_455
timestamp 1679581782
transform 1 0 115296 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_462
timestamp 1679581782
transform 1 0 115968 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_469
timestamp 1679581782
transform 1 0 116640 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_476
timestamp 1679581782
transform 1 0 117312 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_483
timestamp 1679581782
transform 1 0 117984 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_490
timestamp 1679581782
transform 1 0 118656 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_497
timestamp 1679581782
transform 1 0 119328 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_504
timestamp 1679581782
transform 1 0 120000 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_511
timestamp 1679581782
transform 1 0 120672 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_518
timestamp 1679581782
transform 1 0 121344 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_525
timestamp 1679581782
transform 1 0 122016 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_532
timestamp 1679581782
transform 1 0 122688 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_539
timestamp 1679581782
transform 1 0 123360 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_546
timestamp 1679581782
transform 1 0 124032 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_553
timestamp 1679581782
transform 1 0 124704 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_560
timestamp 1679581782
transform 1 0 125376 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_567
timestamp 1679581782
transform 1 0 126048 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_574
timestamp 1679581782
transform 1 0 126720 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_581
timestamp 1679581782
transform 1 0 127392 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_588
timestamp 1679581782
transform 1 0 128064 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_595
timestamp 1679581782
transform 1 0 128736 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_602
timestamp 1679581782
transform 1 0 129408 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_609
timestamp 1679581782
transform 1 0 130080 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_616
timestamp 1679581782
transform 1 0 130752 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_623
timestamp 1679581782
transform 1 0 131424 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_630
timestamp 1679581782
transform 1 0 132096 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_637
timestamp 1679581782
transform 1 0 132768 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_644
timestamp 1679581782
transform 1 0 133440 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_651
timestamp 1679581782
transform 1 0 134112 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_658
timestamp 1679581782
transform 1 0 134784 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_665
timestamp 1679581782
transform 1 0 135456 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_672
timestamp 1679581782
transform 1 0 136128 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_679
timestamp 1679581782
transform 1 0 136800 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_686
timestamp 1679581782
transform 1 0 137472 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_693
timestamp 1679581782
transform 1 0 138144 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_700
timestamp 1679581782
transform 1 0 138816 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_707
timestamp 1679581782
transform 1 0 139488 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_714
timestamp 1679581782
transform 1 0 140160 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_721
timestamp 1679581782
transform 1 0 140832 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_728
timestamp 1679581782
transform 1 0 141504 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_735
timestamp 1679581782
transform 1 0 142176 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_742
timestamp 1679581782
transform 1 0 142848 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_749
timestamp 1679581782
transform 1 0 143520 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_756
timestamp 1679581782
transform 1 0 144192 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_763
timestamp 1679581782
transform 1 0 144864 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_770
timestamp 1679581782
transform 1 0 145536 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_777
timestamp 1679581782
transform 1 0 146208 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_784
timestamp 1679581782
transform 1 0 146880 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_791
timestamp 1679581782
transform 1 0 147552 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_798
timestamp 1679581782
transform 1 0 148224 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_805
timestamp 1679581782
transform 1 0 148896 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_812
timestamp 1679581782
transform 1 0 149568 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_819
timestamp 1679581782
transform 1 0 150240 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_826
timestamp 1679581782
transform 1 0 150912 0 -1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_103_833
timestamp 1679581782
transform 1 0 151584 0 -1 150444
box -48 -56 720 834
use sg13g2_fill_1  FILLER_103_840
timestamp 1677579658
transform 1 0 152256 0 -1 150444
box -48 -56 144 834
use sg13g2_decap_8  FILLER_104_0
timestamp 1679581782
transform 1 0 71616 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_7
timestamp 1679581782
transform 1 0 72288 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_14
timestamp 1679581782
transform 1 0 72960 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_21
timestamp 1679581782
transform 1 0 73632 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_28
timestamp 1679581782
transform 1 0 74304 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_35
timestamp 1679581782
transform 1 0 74976 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_42
timestamp 1679581782
transform 1 0 75648 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_49
timestamp 1679581782
transform 1 0 76320 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_56
timestamp 1679581782
transform 1 0 76992 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_63
timestamp 1679581782
transform 1 0 77664 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_70
timestamp 1679581782
transform 1 0 78336 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_77
timestamp 1679581782
transform 1 0 79008 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_84
timestamp 1679581782
transform 1 0 79680 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_91
timestamp 1679581782
transform 1 0 80352 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_98
timestamp 1679581782
transform 1 0 81024 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_105
timestamp 1679581782
transform 1 0 81696 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_112
timestamp 1679581782
transform 1 0 82368 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_119
timestamp 1679581782
transform 1 0 83040 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_126
timestamp 1679581782
transform 1 0 83712 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_133
timestamp 1679581782
transform 1 0 84384 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_140
timestamp 1679581782
transform 1 0 85056 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_147
timestamp 1679581782
transform 1 0 85728 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_154
timestamp 1679581782
transform 1 0 86400 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_161
timestamp 1679581782
transform 1 0 87072 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_168
timestamp 1679581782
transform 1 0 87744 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_175
timestamp 1679581782
transform 1 0 88416 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_182
timestamp 1679581782
transform 1 0 89088 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_189
timestamp 1679581782
transform 1 0 89760 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_196
timestamp 1679581782
transform 1 0 90432 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_203
timestamp 1679581782
transform 1 0 91104 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_210
timestamp 1679581782
transform 1 0 91776 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_217
timestamp 1679581782
transform 1 0 92448 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_224
timestamp 1679581782
transform 1 0 93120 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_231
timestamp 1679581782
transform 1 0 93792 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_238
timestamp 1679581782
transform 1 0 94464 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_245
timestamp 1679581782
transform 1 0 95136 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_252
timestamp 1679581782
transform 1 0 95808 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_259
timestamp 1679581782
transform 1 0 96480 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_266
timestamp 1679581782
transform 1 0 97152 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_273
timestamp 1679581782
transform 1 0 97824 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_280
timestamp 1679581782
transform 1 0 98496 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_287
timestamp 1679581782
transform 1 0 99168 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_294
timestamp 1679581782
transform 1 0 99840 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_301
timestamp 1679581782
transform 1 0 100512 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_308
timestamp 1679581782
transform 1 0 101184 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_315
timestamp 1679581782
transform 1 0 101856 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_322
timestamp 1679581782
transform 1 0 102528 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_329
timestamp 1679581782
transform 1 0 103200 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_336
timestamp 1679581782
transform 1 0 103872 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_343
timestamp 1679581782
transform 1 0 104544 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_350
timestamp 1679581782
transform 1 0 105216 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_357
timestamp 1679581782
transform 1 0 105888 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_364
timestamp 1679581782
transform 1 0 106560 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_371
timestamp 1679581782
transform 1 0 107232 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_378
timestamp 1679581782
transform 1 0 107904 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_385
timestamp 1679581782
transform 1 0 108576 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_392
timestamp 1679581782
transform 1 0 109248 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_399
timestamp 1679581782
transform 1 0 109920 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_406
timestamp 1679581782
transform 1 0 110592 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_413
timestamp 1679581782
transform 1 0 111264 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_420
timestamp 1679581782
transform 1 0 111936 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_427
timestamp 1679581782
transform 1 0 112608 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_434
timestamp 1679581782
transform 1 0 113280 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_441
timestamp 1679581782
transform 1 0 113952 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_448
timestamp 1679581782
transform 1 0 114624 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_455
timestamp 1679581782
transform 1 0 115296 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_462
timestamp 1679581782
transform 1 0 115968 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_469
timestamp 1679581782
transform 1 0 116640 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_476
timestamp 1679581782
transform 1 0 117312 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_483
timestamp 1679581782
transform 1 0 117984 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_490
timestamp 1679581782
transform 1 0 118656 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_497
timestamp 1679581782
transform 1 0 119328 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_504
timestamp 1679581782
transform 1 0 120000 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_511
timestamp 1679581782
transform 1 0 120672 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_518
timestamp 1679581782
transform 1 0 121344 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_525
timestamp 1679581782
transform 1 0 122016 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_532
timestamp 1679581782
transform 1 0 122688 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_539
timestamp 1679581782
transform 1 0 123360 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_546
timestamp 1679581782
transform 1 0 124032 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_553
timestamp 1679581782
transform 1 0 124704 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_560
timestamp 1679581782
transform 1 0 125376 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_567
timestamp 1679581782
transform 1 0 126048 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_574
timestamp 1679581782
transform 1 0 126720 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_581
timestamp 1679581782
transform 1 0 127392 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_588
timestamp 1679581782
transform 1 0 128064 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_595
timestamp 1679581782
transform 1 0 128736 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_602
timestamp 1679581782
transform 1 0 129408 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_609
timestamp 1679581782
transform 1 0 130080 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_616
timestamp 1679581782
transform 1 0 130752 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_623
timestamp 1679581782
transform 1 0 131424 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_630
timestamp 1679581782
transform 1 0 132096 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_637
timestamp 1679581782
transform 1 0 132768 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_644
timestamp 1679581782
transform 1 0 133440 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_651
timestamp 1679581782
transform 1 0 134112 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_658
timestamp 1679581782
transform 1 0 134784 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_665
timestamp 1679581782
transform 1 0 135456 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_672
timestamp 1679581782
transform 1 0 136128 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_679
timestamp 1679581782
transform 1 0 136800 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_686
timestamp 1679581782
transform 1 0 137472 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_693
timestamp 1679581782
transform 1 0 138144 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_700
timestamp 1679581782
transform 1 0 138816 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_707
timestamp 1679581782
transform 1 0 139488 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_714
timestamp 1679581782
transform 1 0 140160 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_721
timestamp 1679581782
transform 1 0 140832 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_728
timestamp 1679581782
transform 1 0 141504 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_735
timestamp 1679581782
transform 1 0 142176 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_742
timestamp 1679581782
transform 1 0 142848 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_749
timestamp 1679581782
transform 1 0 143520 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_756
timestamp 1679581782
transform 1 0 144192 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_763
timestamp 1679581782
transform 1 0 144864 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_770
timestamp 1679581782
transform 1 0 145536 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_777
timestamp 1679581782
transform 1 0 146208 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_784
timestamp 1679581782
transform 1 0 146880 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_791
timestamp 1679581782
transform 1 0 147552 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_798
timestamp 1679581782
transform 1 0 148224 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_805
timestamp 1679581782
transform 1 0 148896 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_812
timestamp 1679581782
transform 1 0 149568 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_819
timestamp 1679581782
transform 1 0 150240 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_826
timestamp 1679581782
transform 1 0 150912 0 1 150444
box -48 -56 720 834
use sg13g2_decap_8  FILLER_104_833
timestamp 1679581782
transform 1 0 151584 0 1 150444
box -48 -56 720 834
use sg13g2_fill_1  FILLER_104_840
timestamp 1677579658
transform 1 0 152256 0 1 150444
box -48 -56 144 834
use sg13g2_decap_8  FILLER_105_0
timestamp 1679581782
transform 1 0 71616 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_7
timestamp 1679581782
transform 1 0 72288 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_14
timestamp 1679581782
transform 1 0 72960 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_21
timestamp 1679581782
transform 1 0 73632 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_28
timestamp 1679581782
transform 1 0 74304 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_35
timestamp 1679581782
transform 1 0 74976 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_42
timestamp 1679581782
transform 1 0 75648 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_49
timestamp 1679581782
transform 1 0 76320 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_56
timestamp 1679581782
transform 1 0 76992 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_63
timestamp 1679581782
transform 1 0 77664 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_70
timestamp 1679581782
transform 1 0 78336 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_77
timestamp 1679581782
transform 1 0 79008 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_84
timestamp 1679581782
transform 1 0 79680 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_91
timestamp 1679581782
transform 1 0 80352 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_98
timestamp 1679581782
transform 1 0 81024 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_105
timestamp 1679581782
transform 1 0 81696 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_112
timestamp 1679581782
transform 1 0 82368 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_119
timestamp 1679581782
transform 1 0 83040 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_126
timestamp 1679581782
transform 1 0 83712 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_133
timestamp 1679581782
transform 1 0 84384 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_140
timestamp 1679581782
transform 1 0 85056 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_147
timestamp 1679581782
transform 1 0 85728 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_154
timestamp 1679581782
transform 1 0 86400 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_161
timestamp 1679581782
transform 1 0 87072 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_168
timestamp 1679581782
transform 1 0 87744 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_175
timestamp 1679581782
transform 1 0 88416 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_182
timestamp 1679581782
transform 1 0 89088 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_189
timestamp 1679581782
transform 1 0 89760 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_196
timestamp 1679581782
transform 1 0 90432 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_203
timestamp 1679581782
transform 1 0 91104 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_210
timestamp 1679581782
transform 1 0 91776 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_217
timestamp 1679581782
transform 1 0 92448 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_224
timestamp 1679581782
transform 1 0 93120 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_231
timestamp 1679581782
transform 1 0 93792 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_238
timestamp 1679581782
transform 1 0 94464 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_245
timestamp 1679581782
transform 1 0 95136 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_252
timestamp 1679581782
transform 1 0 95808 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_259
timestamp 1679581782
transform 1 0 96480 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_266
timestamp 1679581782
transform 1 0 97152 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_273
timestamp 1679581782
transform 1 0 97824 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_280
timestamp 1679581782
transform 1 0 98496 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_287
timestamp 1679581782
transform 1 0 99168 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_294
timestamp 1679581782
transform 1 0 99840 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_301
timestamp 1679581782
transform 1 0 100512 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_308
timestamp 1679581782
transform 1 0 101184 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_315
timestamp 1679581782
transform 1 0 101856 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_322
timestamp 1679581782
transform 1 0 102528 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_329
timestamp 1679581782
transform 1 0 103200 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_336
timestamp 1679581782
transform 1 0 103872 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_343
timestamp 1679581782
transform 1 0 104544 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_350
timestamp 1679581782
transform 1 0 105216 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_357
timestamp 1679581782
transform 1 0 105888 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_364
timestamp 1679581782
transform 1 0 106560 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_371
timestamp 1679581782
transform 1 0 107232 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_378
timestamp 1679581782
transform 1 0 107904 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_385
timestamp 1679581782
transform 1 0 108576 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_392
timestamp 1679581782
transform 1 0 109248 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_399
timestamp 1679581782
transform 1 0 109920 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_406
timestamp 1679581782
transform 1 0 110592 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_413
timestamp 1679581782
transform 1 0 111264 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_420
timestamp 1679581782
transform 1 0 111936 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_427
timestamp 1679581782
transform 1 0 112608 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_434
timestamp 1679581782
transform 1 0 113280 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_441
timestamp 1679581782
transform 1 0 113952 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_448
timestamp 1679581782
transform 1 0 114624 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_455
timestamp 1679581782
transform 1 0 115296 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_462
timestamp 1679581782
transform 1 0 115968 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_469
timestamp 1679581782
transform 1 0 116640 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_476
timestamp 1679581782
transform 1 0 117312 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_483
timestamp 1679581782
transform 1 0 117984 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_490
timestamp 1679581782
transform 1 0 118656 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_497
timestamp 1679581782
transform 1 0 119328 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_504
timestamp 1679581782
transform 1 0 120000 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_511
timestamp 1679581782
transform 1 0 120672 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_518
timestamp 1679581782
transform 1 0 121344 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_525
timestamp 1679581782
transform 1 0 122016 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_532
timestamp 1679581782
transform 1 0 122688 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_539
timestamp 1679581782
transform 1 0 123360 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_546
timestamp 1679581782
transform 1 0 124032 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_553
timestamp 1679581782
transform 1 0 124704 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_560
timestamp 1679581782
transform 1 0 125376 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_567
timestamp 1679581782
transform 1 0 126048 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_574
timestamp 1679581782
transform 1 0 126720 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_581
timestamp 1679581782
transform 1 0 127392 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_588
timestamp 1679581782
transform 1 0 128064 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_595
timestamp 1679581782
transform 1 0 128736 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_602
timestamp 1679581782
transform 1 0 129408 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_609
timestamp 1679581782
transform 1 0 130080 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_616
timestamp 1679581782
transform 1 0 130752 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_623
timestamp 1679581782
transform 1 0 131424 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_630
timestamp 1679581782
transform 1 0 132096 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_637
timestamp 1679581782
transform 1 0 132768 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_644
timestamp 1679581782
transform 1 0 133440 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_651
timestamp 1679581782
transform 1 0 134112 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_658
timestamp 1679581782
transform 1 0 134784 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_665
timestamp 1679581782
transform 1 0 135456 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_672
timestamp 1679581782
transform 1 0 136128 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_679
timestamp 1679581782
transform 1 0 136800 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_686
timestamp 1679581782
transform 1 0 137472 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_693
timestamp 1679581782
transform 1 0 138144 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_700
timestamp 1679581782
transform 1 0 138816 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_707
timestamp 1679581782
transform 1 0 139488 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_714
timestamp 1679581782
transform 1 0 140160 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_721
timestamp 1679581782
transform 1 0 140832 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_728
timestamp 1679581782
transform 1 0 141504 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_735
timestamp 1679581782
transform 1 0 142176 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_742
timestamp 1679581782
transform 1 0 142848 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_749
timestamp 1679581782
transform 1 0 143520 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_756
timestamp 1679581782
transform 1 0 144192 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_763
timestamp 1679581782
transform 1 0 144864 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_770
timestamp 1679581782
transform 1 0 145536 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_777
timestamp 1679581782
transform 1 0 146208 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_784
timestamp 1679581782
transform 1 0 146880 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_791
timestamp 1679581782
transform 1 0 147552 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_798
timestamp 1679581782
transform 1 0 148224 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_805
timestamp 1679581782
transform 1 0 148896 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_812
timestamp 1679581782
transform 1 0 149568 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_819
timestamp 1679581782
transform 1 0 150240 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_826
timestamp 1679581782
transform 1 0 150912 0 -1 151956
box -48 -56 720 834
use sg13g2_decap_8  FILLER_105_833
timestamp 1679581782
transform 1 0 151584 0 -1 151956
box -48 -56 720 834
use sg13g2_fill_1  FILLER_105_840
timestamp 1677579658
transform 1 0 152256 0 -1 151956
box -48 -56 144 834
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[0\].ui
timestamp 1544787571
transform 0 1 14000 1 0 65000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[1\].ui
timestamp 1544787571
transform 0 1 14000 1 0 81000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[2\].ui
timestamp 1544787571
transform 0 1 14000 1 0 97000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[3\].ui
timestamp 1544787571
transform 0 1 14000 1 0 113000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[4\].ui
timestamp 1544787571
transform 0 1 14000 1 0 129000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[5\].ui
timestamp 1544787571
transform 0 1 14000 1 0 145000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[6\].ui
timestamp 1544787571
transform 1 0 65000 0 1 14000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[7\].ui
timestamp 1544787571
transform 1 0 81000 0 1 14000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[8\].ui
timestamp 1544787571
transform 1 0 97000 0 1 14000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIn_ui\[9\].ui
timestamp 1544787571
transform 1 0 113000 0 1 14000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIOVdd_north
timestamp 1544787571
transform 1 0 65000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadIOVss_north
timestamp 1544787571
transform 1 0 81000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[0\].uo
timestamp 1544787571
transform 0 -1 210000 1 0 65000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[1\].uo
timestamp 1544787571
transform 0 -1 210000 1 0 81000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[2\].uo
timestamp 1544787571
transform 0 -1 210000 1 0 97000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[3\].uo
timestamp 1544787571
transform 0 -1 210000 1 0 113000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[4\].uo
timestamp 1544787571
transform 0 -1 210000 1 0 129000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[5\].uo
timestamp 1544787571
transform 0 -1 210000 1 0 145000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[6\].uo
timestamp 1544787571
transform 1 0 97000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[7\].uo
timestamp 1544787571
transform 1 0 113000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[8\].uo
timestamp 1544787571
transform 1 0 129000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadOut30mA_uo\[9\].uo
timestamp 1544787571
transform 1 0 145000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadVdd_south
timestamp 1544787571
transform 1 0 129000 0 1 14000
box 0 0 14000 14000
use bondpad_70x70  IO_BOND_sg13g2_IOPadVss_south
timestamp 1544787571
transform 1 0 145000 0 1 14000
box 0 0 14000 14000
use sg13g2_Corner  IO_CORNER_NORTH_EAST_INST
timestamp 1716375578
transform -1 0 196000 0 -1 196000
box 1076 1076 36124 36124
use sg13g2_Corner  IO_CORNER_NORTH_WEST_INST
timestamp 1716375578
transform 1 0 28000 0 -1 196000
box 1076 1076 36124 36124
use sg13g2_Corner  IO_CORNER_SOUTH_EAST_INST
timestamp 1716375578
transform -1 0 196000 0 1 28000
box 1076 1076 36124 36124
use sg13g2_Corner  IO_CORNER_SOUTH_WEST_INST
timestamp 1716375578
transform 1 0 28000 0 1 28000
box 1076 1076 36124 36124
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[0\].ui
timestamp 1716375577
transform 0 1 28000 1 0 64000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[1\].ui
timestamp 1716375577
transform 0 1 28000 1 0 80000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[2\].ui
timestamp 1716375577
transform 0 1 28000 1 0 96000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[3\].ui
timestamp 1716375577
transform 0 1 28000 1 0 112000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[4\].ui
timestamp 1716375577
transform 0 1 28000 1 0 128000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[5\].ui
timestamp 1716375577
transform 0 1 28000 1 0 144000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[6\].ui
timestamp 1716375577
transform 1 0 64000 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[7\].ui
timestamp 1716375577
transform 1 0 80000 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[8\].ui
timestamp 1716375577
transform 1 0 96000 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  sg13g2_IOPadIn_ui\[9\].ui
timestamp 1716375577
transform 1 0 112000 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIOVdd  sg13g2_IOPadIOVdd_north
timestamp 1716375578
transform 1 0 64000 0 -1 196000
box -124 0 16124 35600
use sg13g2_IOPadIOVss  sg13g2_IOPadIOVss_north
timestamp 1716375577
transform 1 0 80000 0 -1 196000
box -124 0 16124 35600
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[0\].uo
timestamp 1716375577
transform 0 -1 196000 1 0 64000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[1\].uo
timestamp 1716375577
transform 0 -1 196000 1 0 80000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[2\].uo
timestamp 1716375577
transform 0 -1 196000 1 0 96000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[3\].uo
timestamp 1716375577
transform 0 -1 196000 1 0 112000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[4\].uo
timestamp 1716375577
transform 0 -1 196000 1 0 128000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[5\].uo
timestamp 1716375577
transform 0 -1 196000 1 0 144000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[6\].uo
timestamp 1716375577
transform 1 0 96000 0 -1 196000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[7\].uo
timestamp 1716375577
transform 1 0 112000 0 -1 196000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[8\].uo
timestamp 1716375577
transform 1 0 128000 0 -1 196000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  sg13g2_IOPadOut30mA_uo\[9\].uo
timestamp 1716375577
transform 1 0 144000 0 -1 196000
box -124 0 16124 36000
use sg13g2_IOPadVdd  sg13g2_IOPadVdd_south
timestamp 1716375577
transform 1 0 128000 0 1 28000
box -124 0 16124 35600
use sg13g2_IOPadVss  sg13g2_IOPadVss_south
timestamp 1716375577
transform 1 0 144000 0 1 28000
box -124 0 16124 35600
<< labels >>
flabel metal7 s 65000 196000 79000 210000 0 FreeSans 102400 0 0 0 IO_CORNER_NORTH_WEST_INST.iovdd_RING
port 0 nsew power input
flabel metal7 s 81000 196000 95000 210000 0 FreeSans 102400 0 0 0 IO_CORNER_NORTH_WEST_INST.iovss_RING
port 1 nsew ground input
flabel metal7 s 129000 14000 143000 28000 0 FreeSans 102400 0 0 0 IO_CORNER_NORTH_WEST_INST.vdd_RING
port 2 nsew power input
flabel metal7 s 145000 14000 159000 28000 0 FreeSans 102400 0 0 0 IO_CORNER_NORTH_WEST_INST.vss_RING
port 3 nsew ground input
flabel metal6 s 69716 69920 70716 153856 0 FreeSans 5248 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 69716 69920 154252 70920 0 FreeSans 6400 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 69716 152856 154252 153856 0 FreeSans 6400 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal6 s 153252 69920 154252 153856 0 FreeSans 5248 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 146666 56000 149332 68120 0 FreeSans 12800 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 146666 155656 149332 168000 0 FreeSans 12800 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 130666 155656 133332 168000 0 FreeSans 12800 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 114666 155656 117332 168000 0 FreeSans 12800 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 98666 155656 101332 168000 0 FreeSans 12800 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 153252 146666 168000 149332 0 FreeSans 12800 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 153252 130666 168000 133332 0 FreeSans 12800 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 153252 114666 168000 117332 0 FreeSans 12800 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 153252 98666 168000 101332 0 FreeSans 12800 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 153252 82666 168000 85332 0 FreeSans 12800 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 114666 56000 117332 68120 0 FreeSans 12800 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 98666 56000 101332 68120 0 FreeSans 12800 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 82666 56000 85332 68120 0 FreeSans 12800 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 56000 146666 70716 149332 0 FreeSans 12800 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 56000 130666 70716 133332 0 FreeSans 12800 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 56000 114666 70716 117332 0 FreeSans 12800 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 56000 98666 70716 101332 0 FreeSans 12800 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 56000 82666 70716 85332 0 FreeSans 12800 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 82666 155656 85332 168000 0 FreeSans 12800 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal6 s 74116 68520 74556 155256 0 FreeSans 2624 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal6 s 89236 68520 89676 155256 0 FreeSans 2624 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal6 s 104356 68520 104796 155256 0 FreeSans 2624 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal6 s 119476 68520 119916 155256 0 FreeSans 2624 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal6 s 134596 68520 135036 155256 0 FreeSans 2624 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal6 s 149716 68520 150156 155256 0 FreeSans 2624 90 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 69716 74320 154252 74760 0 FreeSans 3200 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 69716 89440 154252 89880 0 FreeSans 3200 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 69716 104560 154252 105000 0 FreeSans 3200 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 69716 119680 154252 120120 0 FreeSans 3200 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 69716 134800 154252 135240 0 FreeSans 3200 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal7 s 71116 149920 152852 150360 0 FreeSans 3200 0 0 0 VDD
port 4 nsew power bidirectional
flabel metal6 s 68316 68520 69316 155256 0 FreeSans 5248 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 68316 68520 155652 69520 0 FreeSans 6400 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 68316 154256 155652 155256 0 FreeSans 6400 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal6 s 154652 68520 155652 155256 0 FreeSans 5248 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 151998 60000 154664 68120 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 132000 60000 136000 68120 0 FreeSans 25600 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 151998 155656 154664 164000 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 135998 155656 138664 164000 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 119998 155656 122664 164000 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 103998 155656 106664 164000 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 156052 151998 164000 154664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 154652 135998 164000 138664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 154652 119998 164000 122664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 154652 103998 164000 106664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 154652 87998 164000 90664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 154652 71998 164000 74664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 119998 60000 122664 68120 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 103998 60000 106664 68120 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 87998 60000 90664 68120 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 71998 60000 74664 68120 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 60000 151998 67916 154664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 60000 135998 69316 138664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 60000 119998 69316 122664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 60000 103998 69316 106664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 60000 87998 69316 90664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 60000 71998 69316 74664 0 FreeSans 12800 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 87998 155656 90664 164000 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 71998 155656 74664 164000 0 FreeSans 12800 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal6 s 75356 68520 75796 155256 0 FreeSans 2624 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal6 s 90476 68520 90916 155256 0 FreeSans 2624 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal6 s 105596 68520 106036 155256 0 FreeSans 2624 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal6 s 120716 68520 121156 155256 0 FreeSans 2624 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal6 s 135836 68520 136276 155256 0 FreeSans 2624 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal6 s 150956 68520 151396 155256 0 FreeSans 2624 90 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 68316 75560 155652 76000 0 FreeSans 3200 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 68316 151160 155652 151600 0 FreeSans 3200 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 69716 90680 154252 91120 0 FreeSans 3200 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 69716 105800 154252 106240 0 FreeSans 3200 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 69716 120920 154252 121360 0 FreeSans 3200 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 69716 136040 154252 136480 0 FreeSans 3200 0 0 0 VSS
port 5 nsew ground bidirectional
flabel metal7 s 14000 65000 28000 79000 0 FreeSans 102400 0 0 0 ui_PAD[0]
port 6 nsew signal bidirectional
flabel metal7 s 14000 81000 28000 95000 0 FreeSans 102400 0 0 0 ui_PAD[1]
port 7 nsew signal bidirectional
flabel metal7 s 14000 97000 28000 111000 0 FreeSans 102400 0 0 0 ui_PAD[2]
port 8 nsew signal bidirectional
flabel metal7 s 14000 113000 28000 127000 0 FreeSans 102400 0 0 0 ui_PAD[3]
port 9 nsew signal bidirectional
flabel metal7 s 14000 129000 28000 143000 0 FreeSans 102400 0 0 0 ui_PAD[4]
port 10 nsew signal bidirectional
flabel metal7 s 14000 145000 28000 159000 0 FreeSans 102400 0 0 0 ui_PAD[5]
port 11 nsew signal bidirectional
flabel metal7 s 65000 14000 79000 28000 0 FreeSans 102400 0 0 0 ui_PAD[6]
port 12 nsew signal bidirectional
flabel metal7 s 81000 14000 95000 28000 0 FreeSans 102400 0 0 0 ui_PAD[7]
port 13 nsew signal bidirectional
flabel metal7 s 97000 14000 111000 28000 0 FreeSans 102400 0 0 0 ui_PAD[8]
port 14 nsew signal bidirectional
flabel metal7 s 113000 14000 127000 28000 0 FreeSans 102400 0 0 0 ui_PAD[9]
port 15 nsew signal bidirectional
flabel metal7 s 196000 65000 210000 79000 0 FreeSans 102400 0 0 0 uo_PAD[0]
port 16 nsew signal bidirectional
flabel metal7 s 196000 81000 210000 95000 0 FreeSans 102400 0 0 0 uo_PAD[1]
port 17 nsew signal bidirectional
flabel metal7 s 196000 97000 210000 111000 0 FreeSans 102400 0 0 0 uo_PAD[2]
port 18 nsew signal bidirectional
flabel metal7 s 196000 113000 210000 127000 0 FreeSans 102400 0 0 0 uo_PAD[3]
port 19 nsew signal bidirectional
flabel metal7 s 196000 129000 210000 143000 0 FreeSans 102400 0 0 0 uo_PAD[4]
port 20 nsew signal bidirectional
flabel metal7 s 196000 145000 210000 159000 0 FreeSans 102400 0 0 0 uo_PAD[5]
port 21 nsew signal bidirectional
flabel metal7 s 97000 196000 111000 210000 0 FreeSans 102400 0 0 0 uo_PAD[6]
port 22 nsew signal bidirectional
flabel metal7 s 113000 196000 127000 210000 0 FreeSans 102400 0 0 0 uo_PAD[7]
port 23 nsew signal bidirectional
flabel metal7 s 129000 196000 143000 210000 0 FreeSans 102400 0 0 0 uo_PAD[8]
port 24 nsew signal bidirectional
flabel metal7 s 145000 196000 159000 210000 0 FreeSans 102400 0 0 0 uo_PAD[9]
port 25 nsew signal bidirectional
rlabel metal7 111984 150140 111984 150140 0 VDD
rlabel metal7 111984 136260 111984 136260 0 VSS
rlabel metal2 64066 71988 64066 71988 0 ui_PAD2CORE\[0\]
rlabel metal2 64128 88011 64128 88011 0 ui_PAD2CORE\[1\]
rlabel metal2 64066 103992 64066 103992 0 ui_PAD2CORE\[2\]
rlabel metal2 64128 120015 64128 120015 0 ui_PAD2CORE\[3\]
rlabel metal2 64066 135996 64066 135996 0 ui_PAD2CORE\[4\]
rlabel metal2 64128 152019 64128 152019 0 ui_PAD2CORE\[5\]
rlabel metal2 71997 64344 71997 64344 0 ui_PAD2CORE\[6\]
rlabel metal2 119712 159674 119712 159674 0 ui_PAD2CORE\[7\]
rlabel metal2 135744 159716 135744 159716 0 ui_PAD2CORE\[8\]
rlabel metal2 151632 158760 151632 158760 0 ui_PAD2CORE\[9\]
<< properties >>
string FIXED_BBOX 0 0 224000 224000
<< end >>
