magic
tech ihp-sg13g2
magscale 1 2
timestamp 1771591880
<< metal1 >>
rect 75648 148196 148320 148220
rect 75648 148156 79424 148196
rect 79464 148156 79506 148196
rect 79546 148156 79588 148196
rect 79628 148156 79670 148196
rect 79710 148156 79752 148196
rect 79792 148156 94544 148196
rect 94584 148156 94626 148196
rect 94666 148156 94708 148196
rect 94748 148156 94790 148196
rect 94830 148156 94872 148196
rect 94912 148156 109664 148196
rect 109704 148156 109746 148196
rect 109786 148156 109828 148196
rect 109868 148156 109910 148196
rect 109950 148156 109992 148196
rect 110032 148156 124784 148196
rect 124824 148156 124866 148196
rect 124906 148156 124948 148196
rect 124988 148156 125030 148196
rect 125070 148156 125112 148196
rect 125152 148156 139904 148196
rect 139944 148156 139986 148196
rect 140026 148156 140068 148196
rect 140108 148156 140150 148196
rect 140190 148156 140232 148196
rect 140272 148156 148320 148196
rect 75648 148132 148320 148156
rect 75648 147440 148320 147464
rect 75648 147400 78184 147440
rect 78224 147400 78266 147440
rect 78306 147400 78348 147440
rect 78388 147400 78430 147440
rect 78470 147400 78512 147440
rect 78552 147400 93304 147440
rect 93344 147400 93386 147440
rect 93426 147400 93468 147440
rect 93508 147400 93550 147440
rect 93590 147400 93632 147440
rect 93672 147400 108424 147440
rect 108464 147400 108506 147440
rect 108546 147400 108588 147440
rect 108628 147400 108670 147440
rect 108710 147400 108752 147440
rect 108792 147400 123544 147440
rect 123584 147400 123626 147440
rect 123666 147400 123708 147440
rect 123748 147400 123790 147440
rect 123830 147400 123872 147440
rect 123912 147400 138664 147440
rect 138704 147400 138746 147440
rect 138786 147400 138828 147440
rect 138868 147400 138910 147440
rect 138950 147400 138992 147440
rect 139032 147400 148320 147440
rect 75648 147376 148320 147400
rect 75648 146684 148320 146708
rect 75648 146644 79424 146684
rect 79464 146644 79506 146684
rect 79546 146644 79588 146684
rect 79628 146644 79670 146684
rect 79710 146644 79752 146684
rect 79792 146644 94544 146684
rect 94584 146644 94626 146684
rect 94666 146644 94708 146684
rect 94748 146644 94790 146684
rect 94830 146644 94872 146684
rect 94912 146644 109664 146684
rect 109704 146644 109746 146684
rect 109786 146644 109828 146684
rect 109868 146644 109910 146684
rect 109950 146644 109992 146684
rect 110032 146644 124784 146684
rect 124824 146644 124866 146684
rect 124906 146644 124948 146684
rect 124988 146644 125030 146684
rect 125070 146644 125112 146684
rect 125152 146644 139904 146684
rect 139944 146644 139986 146684
rect 140026 146644 140068 146684
rect 140108 146644 140150 146684
rect 140190 146644 140232 146684
rect 140272 146644 148320 146684
rect 75648 146620 148320 146644
rect 75648 145928 148320 145952
rect 75648 145888 78184 145928
rect 78224 145888 78266 145928
rect 78306 145888 78348 145928
rect 78388 145888 78430 145928
rect 78470 145888 78512 145928
rect 78552 145888 93304 145928
rect 93344 145888 93386 145928
rect 93426 145888 93468 145928
rect 93508 145888 93550 145928
rect 93590 145888 93632 145928
rect 93672 145888 108424 145928
rect 108464 145888 108506 145928
rect 108546 145888 108588 145928
rect 108628 145888 108670 145928
rect 108710 145888 108752 145928
rect 108792 145888 123544 145928
rect 123584 145888 123626 145928
rect 123666 145888 123708 145928
rect 123748 145888 123790 145928
rect 123830 145888 123872 145928
rect 123912 145888 138664 145928
rect 138704 145888 138746 145928
rect 138786 145888 138828 145928
rect 138868 145888 138910 145928
rect 138950 145888 138992 145928
rect 139032 145888 148320 145928
rect 75648 145864 148320 145888
rect 75648 145172 148320 145196
rect 75648 145132 79424 145172
rect 79464 145132 79506 145172
rect 79546 145132 79588 145172
rect 79628 145132 79670 145172
rect 79710 145132 79752 145172
rect 79792 145132 94544 145172
rect 94584 145132 94626 145172
rect 94666 145132 94708 145172
rect 94748 145132 94790 145172
rect 94830 145132 94872 145172
rect 94912 145132 109664 145172
rect 109704 145132 109746 145172
rect 109786 145132 109828 145172
rect 109868 145132 109910 145172
rect 109950 145132 109992 145172
rect 110032 145132 124784 145172
rect 124824 145132 124866 145172
rect 124906 145132 124948 145172
rect 124988 145132 125030 145172
rect 125070 145132 125112 145172
rect 125152 145132 139904 145172
rect 139944 145132 139986 145172
rect 140026 145132 140068 145172
rect 140108 145132 140150 145172
rect 140190 145132 140232 145172
rect 140272 145132 148320 145172
rect 75648 145108 148320 145132
rect 75648 144416 148320 144440
rect 75648 144376 78184 144416
rect 78224 144376 78266 144416
rect 78306 144376 78348 144416
rect 78388 144376 78430 144416
rect 78470 144376 78512 144416
rect 78552 144376 93304 144416
rect 93344 144376 93386 144416
rect 93426 144376 93468 144416
rect 93508 144376 93550 144416
rect 93590 144376 93632 144416
rect 93672 144376 108424 144416
rect 108464 144376 108506 144416
rect 108546 144376 108588 144416
rect 108628 144376 108670 144416
rect 108710 144376 108752 144416
rect 108792 144376 123544 144416
rect 123584 144376 123626 144416
rect 123666 144376 123708 144416
rect 123748 144376 123790 144416
rect 123830 144376 123872 144416
rect 123912 144376 138664 144416
rect 138704 144376 138746 144416
rect 138786 144376 138828 144416
rect 138868 144376 138910 144416
rect 138950 144376 138992 144416
rect 139032 144376 148320 144416
rect 75648 144352 148320 144376
rect 75648 143660 148320 143684
rect 75648 143620 79424 143660
rect 79464 143620 79506 143660
rect 79546 143620 79588 143660
rect 79628 143620 79670 143660
rect 79710 143620 79752 143660
rect 79792 143620 94544 143660
rect 94584 143620 94626 143660
rect 94666 143620 94708 143660
rect 94748 143620 94790 143660
rect 94830 143620 94872 143660
rect 94912 143620 109664 143660
rect 109704 143620 109746 143660
rect 109786 143620 109828 143660
rect 109868 143620 109910 143660
rect 109950 143620 109992 143660
rect 110032 143620 124784 143660
rect 124824 143620 124866 143660
rect 124906 143620 124948 143660
rect 124988 143620 125030 143660
rect 125070 143620 125112 143660
rect 125152 143620 139904 143660
rect 139944 143620 139986 143660
rect 140026 143620 140068 143660
rect 140108 143620 140150 143660
rect 140190 143620 140232 143660
rect 140272 143620 148320 143660
rect 75648 143596 148320 143620
rect 75648 142904 148320 142928
rect 75648 142864 78184 142904
rect 78224 142864 78266 142904
rect 78306 142864 78348 142904
rect 78388 142864 78430 142904
rect 78470 142864 78512 142904
rect 78552 142864 93304 142904
rect 93344 142864 93386 142904
rect 93426 142864 93468 142904
rect 93508 142864 93550 142904
rect 93590 142864 93632 142904
rect 93672 142864 108424 142904
rect 108464 142864 108506 142904
rect 108546 142864 108588 142904
rect 108628 142864 108670 142904
rect 108710 142864 108752 142904
rect 108792 142864 123544 142904
rect 123584 142864 123626 142904
rect 123666 142864 123708 142904
rect 123748 142864 123790 142904
rect 123830 142864 123872 142904
rect 123912 142864 138664 142904
rect 138704 142864 138746 142904
rect 138786 142864 138828 142904
rect 138868 142864 138910 142904
rect 138950 142864 138992 142904
rect 139032 142864 148320 142904
rect 75648 142840 148320 142864
rect 75648 142148 148320 142172
rect 75648 142108 79424 142148
rect 79464 142108 79506 142148
rect 79546 142108 79588 142148
rect 79628 142108 79670 142148
rect 79710 142108 79752 142148
rect 79792 142108 94544 142148
rect 94584 142108 94626 142148
rect 94666 142108 94708 142148
rect 94748 142108 94790 142148
rect 94830 142108 94872 142148
rect 94912 142108 109664 142148
rect 109704 142108 109746 142148
rect 109786 142108 109828 142148
rect 109868 142108 109910 142148
rect 109950 142108 109992 142148
rect 110032 142108 124784 142148
rect 124824 142108 124866 142148
rect 124906 142108 124948 142148
rect 124988 142108 125030 142148
rect 125070 142108 125112 142148
rect 125152 142108 139904 142148
rect 139944 142108 139986 142148
rect 140026 142108 140068 142148
rect 140108 142108 140150 142148
rect 140190 142108 140232 142148
rect 140272 142108 148320 142148
rect 75648 142084 148320 142108
rect 75648 141392 148320 141416
rect 75648 141352 78184 141392
rect 78224 141352 78266 141392
rect 78306 141352 78348 141392
rect 78388 141352 78430 141392
rect 78470 141352 78512 141392
rect 78552 141352 93304 141392
rect 93344 141352 93386 141392
rect 93426 141352 93468 141392
rect 93508 141352 93550 141392
rect 93590 141352 93632 141392
rect 93672 141352 108424 141392
rect 108464 141352 108506 141392
rect 108546 141352 108588 141392
rect 108628 141352 108670 141392
rect 108710 141352 108752 141392
rect 108792 141352 123544 141392
rect 123584 141352 123626 141392
rect 123666 141352 123708 141392
rect 123748 141352 123790 141392
rect 123830 141352 123872 141392
rect 123912 141352 138664 141392
rect 138704 141352 138746 141392
rect 138786 141352 138828 141392
rect 138868 141352 138910 141392
rect 138950 141352 138992 141392
rect 139032 141352 148320 141392
rect 75648 141328 148320 141352
rect 75648 140636 148320 140660
rect 75648 140596 79424 140636
rect 79464 140596 79506 140636
rect 79546 140596 79588 140636
rect 79628 140596 79670 140636
rect 79710 140596 79752 140636
rect 79792 140596 94544 140636
rect 94584 140596 94626 140636
rect 94666 140596 94708 140636
rect 94748 140596 94790 140636
rect 94830 140596 94872 140636
rect 94912 140596 109664 140636
rect 109704 140596 109746 140636
rect 109786 140596 109828 140636
rect 109868 140596 109910 140636
rect 109950 140596 109992 140636
rect 110032 140596 124784 140636
rect 124824 140596 124866 140636
rect 124906 140596 124948 140636
rect 124988 140596 125030 140636
rect 125070 140596 125112 140636
rect 125152 140596 139904 140636
rect 139944 140596 139986 140636
rect 140026 140596 140068 140636
rect 140108 140596 140150 140636
rect 140190 140596 140232 140636
rect 140272 140596 148320 140636
rect 75648 140572 148320 140596
rect 75648 139880 148320 139904
rect 75648 139840 78184 139880
rect 78224 139840 78266 139880
rect 78306 139840 78348 139880
rect 78388 139840 78430 139880
rect 78470 139840 78512 139880
rect 78552 139840 93304 139880
rect 93344 139840 93386 139880
rect 93426 139840 93468 139880
rect 93508 139840 93550 139880
rect 93590 139840 93632 139880
rect 93672 139840 108424 139880
rect 108464 139840 108506 139880
rect 108546 139840 108588 139880
rect 108628 139840 108670 139880
rect 108710 139840 108752 139880
rect 108792 139840 123544 139880
rect 123584 139840 123626 139880
rect 123666 139840 123708 139880
rect 123748 139840 123790 139880
rect 123830 139840 123872 139880
rect 123912 139840 138664 139880
rect 138704 139840 138746 139880
rect 138786 139840 138828 139880
rect 138868 139840 138910 139880
rect 138950 139840 138992 139880
rect 139032 139840 148320 139880
rect 75648 139816 148320 139840
rect 75648 139124 148320 139148
rect 75648 139084 79424 139124
rect 79464 139084 79506 139124
rect 79546 139084 79588 139124
rect 79628 139084 79670 139124
rect 79710 139084 79752 139124
rect 79792 139084 94544 139124
rect 94584 139084 94626 139124
rect 94666 139084 94708 139124
rect 94748 139084 94790 139124
rect 94830 139084 94872 139124
rect 94912 139084 109664 139124
rect 109704 139084 109746 139124
rect 109786 139084 109828 139124
rect 109868 139084 109910 139124
rect 109950 139084 109992 139124
rect 110032 139084 124784 139124
rect 124824 139084 124866 139124
rect 124906 139084 124948 139124
rect 124988 139084 125030 139124
rect 125070 139084 125112 139124
rect 125152 139084 139904 139124
rect 139944 139084 139986 139124
rect 140026 139084 140068 139124
rect 140108 139084 140150 139124
rect 140190 139084 140232 139124
rect 140272 139084 148320 139124
rect 75648 139060 148320 139084
rect 75648 138368 148320 138392
rect 75648 138328 78184 138368
rect 78224 138328 78266 138368
rect 78306 138328 78348 138368
rect 78388 138328 78430 138368
rect 78470 138328 78512 138368
rect 78552 138328 93304 138368
rect 93344 138328 93386 138368
rect 93426 138328 93468 138368
rect 93508 138328 93550 138368
rect 93590 138328 93632 138368
rect 93672 138328 108424 138368
rect 108464 138328 108506 138368
rect 108546 138328 108588 138368
rect 108628 138328 108670 138368
rect 108710 138328 108752 138368
rect 108792 138328 123544 138368
rect 123584 138328 123626 138368
rect 123666 138328 123708 138368
rect 123748 138328 123790 138368
rect 123830 138328 123872 138368
rect 123912 138328 138664 138368
rect 138704 138328 138746 138368
rect 138786 138328 138828 138368
rect 138868 138328 138910 138368
rect 138950 138328 138992 138368
rect 139032 138328 148320 138368
rect 75648 138304 148320 138328
rect 75648 137612 148320 137636
rect 75648 137572 79424 137612
rect 79464 137572 79506 137612
rect 79546 137572 79588 137612
rect 79628 137572 79670 137612
rect 79710 137572 79752 137612
rect 79792 137572 94544 137612
rect 94584 137572 94626 137612
rect 94666 137572 94708 137612
rect 94748 137572 94790 137612
rect 94830 137572 94872 137612
rect 94912 137572 109664 137612
rect 109704 137572 109746 137612
rect 109786 137572 109828 137612
rect 109868 137572 109910 137612
rect 109950 137572 109992 137612
rect 110032 137572 124784 137612
rect 124824 137572 124866 137612
rect 124906 137572 124948 137612
rect 124988 137572 125030 137612
rect 125070 137572 125112 137612
rect 125152 137572 139904 137612
rect 139944 137572 139986 137612
rect 140026 137572 140068 137612
rect 140108 137572 140150 137612
rect 140190 137572 140232 137612
rect 140272 137572 148320 137612
rect 75648 137548 148320 137572
rect 75648 136856 148320 136880
rect 75648 136816 78184 136856
rect 78224 136816 78266 136856
rect 78306 136816 78348 136856
rect 78388 136816 78430 136856
rect 78470 136816 78512 136856
rect 78552 136816 93304 136856
rect 93344 136816 93386 136856
rect 93426 136816 93468 136856
rect 93508 136816 93550 136856
rect 93590 136816 93632 136856
rect 93672 136816 108424 136856
rect 108464 136816 108506 136856
rect 108546 136816 108588 136856
rect 108628 136816 108670 136856
rect 108710 136816 108752 136856
rect 108792 136816 123544 136856
rect 123584 136816 123626 136856
rect 123666 136816 123708 136856
rect 123748 136816 123790 136856
rect 123830 136816 123872 136856
rect 123912 136816 138664 136856
rect 138704 136816 138746 136856
rect 138786 136816 138828 136856
rect 138868 136816 138910 136856
rect 138950 136816 138992 136856
rect 139032 136816 148320 136856
rect 75648 136792 148320 136816
rect 75648 136100 148320 136124
rect 75648 136060 79424 136100
rect 79464 136060 79506 136100
rect 79546 136060 79588 136100
rect 79628 136060 79670 136100
rect 79710 136060 79752 136100
rect 79792 136060 94544 136100
rect 94584 136060 94626 136100
rect 94666 136060 94708 136100
rect 94748 136060 94790 136100
rect 94830 136060 94872 136100
rect 94912 136060 109664 136100
rect 109704 136060 109746 136100
rect 109786 136060 109828 136100
rect 109868 136060 109910 136100
rect 109950 136060 109992 136100
rect 110032 136060 124784 136100
rect 124824 136060 124866 136100
rect 124906 136060 124948 136100
rect 124988 136060 125030 136100
rect 125070 136060 125112 136100
rect 125152 136060 139904 136100
rect 139944 136060 139986 136100
rect 140026 136060 140068 136100
rect 140108 136060 140150 136100
rect 140190 136060 140232 136100
rect 140272 136060 148320 136100
rect 75648 136036 148320 136060
rect 75648 135344 148320 135368
rect 75648 135304 78184 135344
rect 78224 135304 78266 135344
rect 78306 135304 78348 135344
rect 78388 135304 78430 135344
rect 78470 135304 78512 135344
rect 78552 135304 93304 135344
rect 93344 135304 93386 135344
rect 93426 135304 93468 135344
rect 93508 135304 93550 135344
rect 93590 135304 93632 135344
rect 93672 135304 108424 135344
rect 108464 135304 108506 135344
rect 108546 135304 108588 135344
rect 108628 135304 108670 135344
rect 108710 135304 108752 135344
rect 108792 135304 123544 135344
rect 123584 135304 123626 135344
rect 123666 135304 123708 135344
rect 123748 135304 123790 135344
rect 123830 135304 123872 135344
rect 123912 135304 138664 135344
rect 138704 135304 138746 135344
rect 138786 135304 138828 135344
rect 138868 135304 138910 135344
rect 138950 135304 138992 135344
rect 139032 135304 148320 135344
rect 75648 135280 148320 135304
rect 75648 134588 148320 134612
rect 75648 134548 79424 134588
rect 79464 134548 79506 134588
rect 79546 134548 79588 134588
rect 79628 134548 79670 134588
rect 79710 134548 79752 134588
rect 79792 134548 94544 134588
rect 94584 134548 94626 134588
rect 94666 134548 94708 134588
rect 94748 134548 94790 134588
rect 94830 134548 94872 134588
rect 94912 134548 109664 134588
rect 109704 134548 109746 134588
rect 109786 134548 109828 134588
rect 109868 134548 109910 134588
rect 109950 134548 109992 134588
rect 110032 134548 124784 134588
rect 124824 134548 124866 134588
rect 124906 134548 124948 134588
rect 124988 134548 125030 134588
rect 125070 134548 125112 134588
rect 125152 134548 139904 134588
rect 139944 134548 139986 134588
rect 140026 134548 140068 134588
rect 140108 134548 140150 134588
rect 140190 134548 140232 134588
rect 140272 134548 148320 134588
rect 75648 134524 148320 134548
rect 115939 134420 115997 134421
rect 115939 134380 115948 134420
rect 115988 134380 115997 134420
rect 115939 134379 115997 134380
rect 97419 134252 97461 134261
rect 97419 134212 97420 134252
rect 97460 134212 97461 134252
rect 97419 134203 97461 134212
rect 97795 134252 97853 134253
rect 97795 134212 97804 134252
rect 97844 134212 97853 134252
rect 97795 134211 97853 134212
rect 98659 134252 98717 134253
rect 98659 134212 98668 134252
rect 98708 134212 98717 134252
rect 98659 134211 98717 134212
rect 113547 134252 113589 134261
rect 113547 134212 113548 134252
rect 113588 134212 113589 134252
rect 113547 134203 113589 134212
rect 113923 134252 113981 134253
rect 113923 134212 113932 134252
rect 113972 134212 113981 134252
rect 113923 134211 113981 134212
rect 114787 134252 114845 134253
rect 114787 134212 114796 134252
rect 114836 134212 114845 134252
rect 114787 134211 114845 134212
rect 99811 134084 99869 134085
rect 99811 134044 99820 134084
rect 99860 134044 99869 134084
rect 99811 134043 99869 134044
rect 119883 134084 119925 134093
rect 119883 134044 119884 134084
rect 119924 134044 119925 134084
rect 119883 134035 119925 134044
rect 115939 134000 115997 134001
rect 115939 133960 115948 134000
rect 115988 133960 115997 134000
rect 115939 133959 115997 133960
rect 75648 133832 148320 133856
rect 75648 133792 78184 133832
rect 78224 133792 78266 133832
rect 78306 133792 78348 133832
rect 78388 133792 78430 133832
rect 78470 133792 78512 133832
rect 78552 133792 93304 133832
rect 93344 133792 93386 133832
rect 93426 133792 93468 133832
rect 93508 133792 93550 133832
rect 93590 133792 93632 133832
rect 93672 133792 108424 133832
rect 108464 133792 108506 133832
rect 108546 133792 108588 133832
rect 108628 133792 108670 133832
rect 108710 133792 108752 133832
rect 108792 133792 123544 133832
rect 123584 133792 123626 133832
rect 123666 133792 123708 133832
rect 123748 133792 123790 133832
rect 123830 133792 123872 133832
rect 123912 133792 138664 133832
rect 138704 133792 138746 133832
rect 138786 133792 138828 133832
rect 138868 133792 138910 133832
rect 138950 133792 138992 133832
rect 139032 133792 148320 133832
rect 75648 133768 148320 133792
rect 98179 133664 98237 133665
rect 98179 133624 98188 133664
rect 98228 133624 98237 133664
rect 98179 133623 98237 133624
rect 121795 133664 121853 133665
rect 121795 133624 121804 133664
rect 121844 133624 121853 133664
rect 121795 133623 121853 133624
rect 97803 133580 97845 133589
rect 97803 133540 97804 133580
rect 97844 133540 97845 133580
rect 97803 133531 97845 133540
rect 114027 133580 114069 133589
rect 114027 133540 114028 133580
rect 114068 133540 114069 133580
rect 114027 133531 114069 133540
rect 98851 133412 98909 133413
rect 98851 133372 98860 133412
rect 98900 133372 98909 133412
rect 98851 133371 98909 133372
rect 115075 133412 115133 133413
rect 115075 133372 115084 133412
rect 115124 133372 115133 133412
rect 115075 133371 115133 133372
rect 119779 133412 119837 133413
rect 119779 133372 119788 133412
rect 119828 133372 119837 133412
rect 119779 133371 119837 133372
rect 120643 133412 120701 133413
rect 120643 133372 120652 133412
rect 120692 133372 120701 133412
rect 120643 133371 120701 133372
rect 119403 133328 119445 133337
rect 119403 133288 119404 133328
rect 119444 133288 119445 133328
rect 119403 133279 119445 133288
rect 114403 133244 114461 133245
rect 114403 133204 114412 133244
rect 114452 133204 114461 133244
rect 114403 133203 114461 133204
rect 121795 133244 121853 133245
rect 121795 133204 121804 133244
rect 121844 133204 121853 133244
rect 121795 133203 121853 133204
rect 75648 133076 148320 133100
rect 75648 133036 79424 133076
rect 79464 133036 79506 133076
rect 79546 133036 79588 133076
rect 79628 133036 79670 133076
rect 79710 133036 79752 133076
rect 79792 133036 94544 133076
rect 94584 133036 94626 133076
rect 94666 133036 94708 133076
rect 94748 133036 94790 133076
rect 94830 133036 94872 133076
rect 94912 133036 109664 133076
rect 109704 133036 109746 133076
rect 109786 133036 109828 133076
rect 109868 133036 109910 133076
rect 109950 133036 109992 133076
rect 110032 133036 124784 133076
rect 124824 133036 124866 133076
rect 124906 133036 124948 133076
rect 124988 133036 125030 133076
rect 125070 133036 125112 133076
rect 125152 133036 139904 133076
rect 139944 133036 139986 133076
rect 140026 133036 140068 133076
rect 140108 133036 140150 133076
rect 140190 133036 140232 133076
rect 140272 133036 148320 133076
rect 75648 133012 148320 133036
rect 98659 132908 98717 132909
rect 98659 132868 98668 132908
rect 98708 132868 98717 132908
rect 98659 132867 98717 132868
rect 119395 132908 119453 132909
rect 119395 132868 119404 132908
rect 119444 132868 119453 132908
rect 119395 132867 119453 132868
rect 78595 132740 78653 132741
rect 78595 132700 78604 132740
rect 78644 132700 78653 132740
rect 78595 132699 78653 132700
rect 98571 132740 98613 132749
rect 98571 132700 98572 132740
rect 98612 132700 98613 132740
rect 98571 132691 98613 132700
rect 98763 132740 98805 132749
rect 98763 132700 98764 132740
rect 98804 132700 98805 132740
rect 98763 132691 98805 132700
rect 98851 132740 98909 132741
rect 98851 132700 98860 132740
rect 98900 132700 98909 132740
rect 98851 132699 98909 132700
rect 102979 132740 103037 132741
rect 102979 132700 102988 132740
rect 103028 132700 103037 132740
rect 102979 132699 103037 132700
rect 103659 132740 103701 132749
rect 103659 132700 103660 132740
rect 103700 132700 103701 132740
rect 103659 132691 103701 132700
rect 103851 132740 103893 132749
rect 103851 132700 103852 132740
rect 103892 132700 103893 132740
rect 103851 132691 103893 132700
rect 104227 132740 104285 132741
rect 104227 132700 104236 132740
rect 104276 132700 104285 132740
rect 104227 132699 104285 132700
rect 105091 132740 105149 132741
rect 105091 132700 105100 132740
rect 105140 132700 105149 132740
rect 105091 132699 105149 132700
rect 120067 132740 120125 132741
rect 120067 132700 120076 132740
rect 120116 132700 120125 132740
rect 120067 132699 120125 132700
rect 120931 132740 120989 132741
rect 120931 132700 120940 132740
rect 120980 132700 120989 132740
rect 120931 132699 120989 132700
rect 106251 132656 106293 132665
rect 106251 132616 106252 132656
rect 106292 132616 106293 132656
rect 106251 132607 106293 132616
rect 79267 132572 79325 132573
rect 79267 132532 79276 132572
rect 79316 132532 79325 132572
rect 79267 132531 79325 132532
rect 109899 132572 109941 132581
rect 109899 132532 109900 132572
rect 109940 132532 109941 132572
rect 109899 132523 109941 132532
rect 120259 132572 120317 132573
rect 120259 132532 120268 132572
rect 120308 132532 120317 132572
rect 120259 132531 120317 132532
rect 75648 132320 148320 132344
rect 75648 132280 78184 132320
rect 78224 132280 78266 132320
rect 78306 132280 78348 132320
rect 78388 132280 78430 132320
rect 78470 132280 78512 132320
rect 78552 132280 93304 132320
rect 93344 132280 93386 132320
rect 93426 132280 93468 132320
rect 93508 132280 93550 132320
rect 93590 132280 93632 132320
rect 93672 132280 108424 132320
rect 108464 132280 108506 132320
rect 108546 132280 108588 132320
rect 108628 132280 108670 132320
rect 108710 132280 108752 132320
rect 108792 132280 123544 132320
rect 123584 132280 123626 132320
rect 123666 132280 123708 132320
rect 123748 132280 123790 132320
rect 123830 132280 123872 132320
rect 123912 132280 138664 132320
rect 138704 132280 138746 132320
rect 138786 132280 138828 132320
rect 138868 132280 138910 132320
rect 138950 132280 138992 132320
rect 139032 132280 148320 132320
rect 75648 132256 148320 132280
rect 99043 132068 99101 132069
rect 99043 132028 99052 132068
rect 99092 132028 99101 132068
rect 99043 132027 99101 132028
rect 104331 132068 104373 132077
rect 104331 132028 104332 132068
rect 104372 132028 104373 132068
rect 104331 132019 104373 132028
rect 98371 131900 98429 131901
rect 98371 131860 98380 131900
rect 98420 131860 98429 131900
rect 98371 131859 98429 131860
rect 99243 131900 99285 131909
rect 99243 131860 99244 131900
rect 99284 131860 99285 131900
rect 99243 131851 99285 131860
rect 99339 131900 99381 131909
rect 99339 131860 99340 131900
rect 99380 131860 99381 131900
rect 99339 131851 99381 131860
rect 99435 131900 99477 131909
rect 99435 131860 99436 131900
rect 99476 131860 99477 131900
rect 99435 131851 99477 131860
rect 99531 131900 99573 131909
rect 99531 131860 99532 131900
rect 99572 131860 99573 131900
rect 99531 131851 99573 131860
rect 100011 131900 100053 131909
rect 100011 131860 100012 131900
rect 100052 131860 100053 131900
rect 100011 131851 100053 131860
rect 100195 131900 100253 131901
rect 100195 131860 100204 131900
rect 100244 131860 100253 131900
rect 100195 131859 100253 131860
rect 101059 131900 101117 131901
rect 101059 131860 101068 131900
rect 101108 131860 101117 131900
rect 101059 131859 101117 131860
rect 101163 131900 101205 131909
rect 101163 131860 101164 131900
rect 101204 131860 101205 131900
rect 101163 131851 101205 131860
rect 101355 131900 101397 131909
rect 101355 131860 101356 131900
rect 101396 131860 101397 131900
rect 101355 131851 101397 131860
rect 101635 131900 101693 131901
rect 101635 131860 101644 131900
rect 101684 131860 101693 131900
rect 101635 131859 101693 131860
rect 109795 131900 109853 131901
rect 109795 131860 109804 131900
rect 109844 131860 109853 131900
rect 109795 131859 109853 131860
rect 110659 131900 110717 131901
rect 110659 131860 110668 131900
rect 110708 131860 110717 131900
rect 110659 131859 110717 131860
rect 112203 131900 112245 131909
rect 112203 131860 112204 131900
rect 112244 131860 112245 131900
rect 112203 131851 112245 131860
rect 112299 131900 112341 131909
rect 112299 131860 112300 131900
rect 112340 131860 112341 131900
rect 112299 131851 112341 131860
rect 112771 131900 112829 131901
rect 112771 131860 112780 131900
rect 112820 131860 112829 131900
rect 112771 131859 112829 131860
rect 118531 131900 118589 131901
rect 118531 131860 118540 131900
rect 118580 131860 118589 131900
rect 118531 131859 118589 131860
rect 100107 131816 100149 131825
rect 100107 131776 100108 131816
rect 100148 131776 100149 131816
rect 100107 131767 100149 131776
rect 109419 131816 109461 131825
rect 109419 131776 109420 131816
rect 109460 131776 109461 131816
rect 109419 131767 109461 131776
rect 112395 131816 112453 131817
rect 112395 131776 112404 131816
rect 112444 131776 112453 131816
rect 112395 131775 112453 131776
rect 101251 131732 101309 131733
rect 101251 131692 101260 131732
rect 101300 131692 101309 131732
rect 101251 131691 101309 131692
rect 101547 131732 101589 131741
rect 101547 131692 101548 131732
rect 101588 131692 101589 131732
rect 101547 131683 101589 131692
rect 111811 131732 111869 131733
rect 111811 131692 111820 131732
rect 111860 131692 111869 131732
rect 111811 131691 111869 131692
rect 112483 131732 112541 131733
rect 112483 131692 112492 131732
rect 112532 131692 112541 131732
rect 112483 131691 112541 131692
rect 112587 131732 112629 131741
rect 112587 131692 112588 131732
rect 112628 131692 112629 131732
rect 112587 131683 112629 131692
rect 113443 131732 113501 131733
rect 113443 131692 113452 131732
rect 113492 131692 113501 131732
rect 113443 131691 113501 131692
rect 118443 131732 118485 131741
rect 118443 131692 118444 131732
rect 118484 131692 118485 131732
rect 118443 131683 118485 131692
rect 75648 131564 148320 131588
rect 75648 131524 79424 131564
rect 79464 131524 79506 131564
rect 79546 131524 79588 131564
rect 79628 131524 79670 131564
rect 79710 131524 79752 131564
rect 79792 131524 94544 131564
rect 94584 131524 94626 131564
rect 94666 131524 94708 131564
rect 94748 131524 94790 131564
rect 94830 131524 94872 131564
rect 94912 131524 109664 131564
rect 109704 131524 109746 131564
rect 109786 131524 109828 131564
rect 109868 131524 109910 131564
rect 109950 131524 109992 131564
rect 110032 131524 124784 131564
rect 124824 131524 124866 131564
rect 124906 131524 124948 131564
rect 124988 131524 125030 131564
rect 125070 131524 125112 131564
rect 125152 131524 139904 131564
rect 139944 131524 139986 131564
rect 140026 131524 140068 131564
rect 140108 131524 140150 131564
rect 140190 131524 140232 131564
rect 140272 131524 148320 131564
rect 75648 131500 148320 131524
rect 102219 131396 102261 131405
rect 102219 131356 102220 131396
rect 102260 131356 102261 131396
rect 102219 131347 102261 131356
rect 108835 131396 108893 131397
rect 108835 131356 108844 131396
rect 108884 131356 108893 131396
rect 108835 131355 108893 131356
rect 109795 131396 109853 131397
rect 109795 131356 109804 131396
rect 109844 131356 109853 131396
rect 109795 131355 109853 131356
rect 110755 131396 110813 131397
rect 110755 131356 110764 131396
rect 110804 131356 110813 131396
rect 110755 131355 110813 131356
rect 112291 131396 112349 131397
rect 112291 131356 112300 131396
rect 112340 131356 112349 131396
rect 112291 131355 112349 131356
rect 113059 131396 113117 131397
rect 113059 131356 113068 131396
rect 113108 131356 113117 131396
rect 113059 131355 113117 131356
rect 115171 131396 115229 131397
rect 115171 131356 115180 131396
rect 115220 131356 115229 131396
rect 115171 131355 115229 131356
rect 119299 131396 119357 131397
rect 119299 131356 119308 131396
rect 119348 131356 119357 131396
rect 119299 131355 119357 131356
rect 113347 131312 113405 131313
rect 113347 131272 113356 131312
rect 113396 131272 113405 131312
rect 113347 131271 113405 131272
rect 115075 131312 115133 131313
rect 115075 131272 115084 131312
rect 115124 131272 115133 131312
rect 115075 131271 115133 131272
rect 99907 131228 99965 131229
rect 99907 131188 99916 131228
rect 99956 131188 99965 131228
rect 99907 131187 99965 131188
rect 100587 131228 100629 131237
rect 100587 131188 100588 131228
rect 100628 131188 100629 131228
rect 100587 131179 100629 131188
rect 102027 131228 102069 131237
rect 102027 131188 102028 131228
rect 102068 131188 102069 131228
rect 102027 131179 102069 131188
rect 102123 131228 102165 131237
rect 102123 131188 102124 131228
rect 102164 131188 102165 131228
rect 102123 131179 102165 131188
rect 102315 131228 102357 131237
rect 102315 131188 102316 131228
rect 102356 131188 102357 131228
rect 102315 131179 102357 131188
rect 103171 131228 103229 131229
rect 103171 131188 103180 131228
rect 103220 131188 103229 131228
rect 103171 131187 103229 131188
rect 103363 131228 103421 131229
rect 103363 131188 103372 131228
rect 103412 131188 103421 131228
rect 103363 131187 103421 131188
rect 108939 131228 108981 131237
rect 108939 131188 108940 131228
rect 108980 131188 108981 131228
rect 108939 131179 108981 131188
rect 109035 131228 109077 131237
rect 109035 131188 109036 131228
rect 109076 131188 109077 131228
rect 109035 131179 109077 131188
rect 109131 131228 109173 131237
rect 109131 131188 109132 131228
rect 109172 131188 109173 131228
rect 109131 131179 109173 131188
rect 109323 131228 109365 131237
rect 109323 131188 109324 131228
rect 109364 131188 109365 131228
rect 109323 131179 109365 131188
rect 109419 131228 109461 131237
rect 109419 131188 109420 131228
rect 109460 131188 109461 131228
rect 109419 131179 109461 131188
rect 109611 131228 109653 131237
rect 109611 131188 109612 131228
rect 109652 131188 109653 131228
rect 109611 131179 109653 131188
rect 110467 131228 110525 131229
rect 110467 131188 110476 131228
rect 110516 131188 110525 131228
rect 110467 131187 110525 131188
rect 111427 131228 111485 131229
rect 111427 131188 111436 131228
rect 111476 131188 111485 131228
rect 111427 131187 111485 131188
rect 112491 131228 112533 131237
rect 112491 131188 112492 131228
rect 112532 131188 112533 131228
rect 112491 131179 112533 131188
rect 112587 131228 112629 131237
rect 112587 131188 112588 131228
rect 112628 131188 112629 131228
rect 112587 131179 112629 131188
rect 113067 131228 113109 131237
rect 113067 131188 113068 131228
rect 113108 131188 113109 131228
rect 113067 131179 113109 131188
rect 113163 131228 113205 131237
rect 113163 131188 113164 131228
rect 113204 131188 113205 131228
rect 113163 131179 113205 131188
rect 114891 131228 114933 131237
rect 114891 131188 114892 131228
rect 114932 131188 114933 131228
rect 114891 131179 114933 131188
rect 114987 131228 115029 131237
rect 114987 131188 114988 131228
rect 115028 131188 115029 131228
rect 114987 131179 115029 131188
rect 119107 131228 119165 131229
rect 119107 131188 119116 131228
rect 119156 131188 119165 131228
rect 119107 131187 119165 131188
rect 119211 131228 119253 131237
rect 119211 131188 119212 131228
rect 119252 131188 119253 131228
rect 119211 131179 119253 131188
rect 119403 131228 119445 131237
rect 119403 131188 119404 131228
rect 119444 131188 119445 131228
rect 119403 131179 119445 131188
rect 104035 131060 104093 131061
rect 104035 131020 104044 131060
rect 104084 131020 104093 131060
rect 104035 131019 104093 131020
rect 102499 130976 102557 130977
rect 102499 130936 102508 130976
rect 102548 130936 102557 130976
rect 102499 130935 102557 130936
rect 115179 130976 115221 130985
rect 115179 130936 115180 130976
rect 115220 130936 115221 130976
rect 115179 130927 115221 130936
rect 75648 130808 148320 130832
rect 75648 130768 78184 130808
rect 78224 130768 78266 130808
rect 78306 130768 78348 130808
rect 78388 130768 78430 130808
rect 78470 130768 78512 130808
rect 78552 130768 93304 130808
rect 93344 130768 93386 130808
rect 93426 130768 93468 130808
rect 93508 130768 93550 130808
rect 93590 130768 93632 130808
rect 93672 130768 108424 130808
rect 108464 130768 108506 130808
rect 108546 130768 108588 130808
rect 108628 130768 108670 130808
rect 108710 130768 108752 130808
rect 108792 130768 123544 130808
rect 123584 130768 123626 130808
rect 123666 130768 123708 130808
rect 123748 130768 123790 130808
rect 123830 130768 123872 130808
rect 123912 130768 138664 130808
rect 138704 130768 138746 130808
rect 138786 130768 138828 130808
rect 138868 130768 138910 130808
rect 138950 130768 138992 130808
rect 139032 130768 148320 130808
rect 75648 130744 148320 130768
rect 98091 130640 98133 130649
rect 98091 130600 98092 130640
rect 98132 130600 98133 130640
rect 98091 130591 98133 130600
rect 102603 130640 102645 130649
rect 102603 130600 102604 130640
rect 102644 130600 102645 130640
rect 102603 130591 102645 130600
rect 110475 130640 110517 130649
rect 110475 130600 110476 130640
rect 110516 130600 110517 130640
rect 110475 130591 110517 130600
rect 117579 130640 117621 130649
rect 117579 130600 117580 130640
rect 117620 130600 117621 130640
rect 117579 130591 117621 130600
rect 103075 130556 103133 130557
rect 103075 130516 103084 130556
rect 103124 130516 103133 130556
rect 103075 130515 103133 130516
rect 108739 130472 108797 130473
rect 108739 130432 108748 130472
rect 108788 130432 108797 130472
rect 108739 130431 108797 130432
rect 98091 130388 98133 130397
rect 97902 130377 97960 130378
rect 97902 130337 97911 130377
rect 97951 130337 97960 130377
rect 98091 130348 98092 130388
rect 98132 130348 98133 130388
rect 98091 130339 98133 130348
rect 102499 130388 102557 130389
rect 102499 130348 102508 130388
rect 102548 130348 102557 130388
rect 102499 130347 102557 130348
rect 102795 130388 102837 130397
rect 102795 130348 102796 130388
rect 102836 130348 102837 130388
rect 102795 130339 102837 130348
rect 102987 130388 103029 130397
rect 102987 130348 102988 130388
rect 103028 130348 103029 130388
rect 102987 130339 103029 130348
rect 103083 130388 103125 130397
rect 103083 130348 103084 130388
rect 103124 130348 103125 130388
rect 103083 130339 103125 130348
rect 105379 130388 105437 130389
rect 105379 130348 105388 130388
rect 105428 130348 105437 130388
rect 105379 130347 105437 130348
rect 110179 130388 110237 130389
rect 110179 130348 110188 130388
rect 110228 130348 110237 130388
rect 110179 130347 110237 130348
rect 110467 130388 110525 130389
rect 110467 130348 110476 130388
rect 110516 130348 110525 130388
rect 110467 130347 110525 130348
rect 110667 130388 110709 130397
rect 110667 130348 110668 130388
rect 110708 130348 110709 130388
rect 110667 130339 110709 130348
rect 110755 130388 110813 130389
rect 110755 130348 110764 130388
rect 110804 130348 110813 130388
rect 110755 130347 110813 130348
rect 117483 130388 117525 130397
rect 117483 130348 117484 130388
rect 117524 130348 117525 130388
rect 117483 130339 117525 130348
rect 117667 130388 117725 130389
rect 117667 130348 117676 130388
rect 117716 130348 117725 130388
rect 117667 130347 117725 130348
rect 97902 130336 97960 130337
rect 104707 130220 104765 130221
rect 104707 130180 104716 130220
rect 104756 130180 104765 130220
rect 104707 130179 104765 130180
rect 75648 130052 148320 130076
rect 75648 130012 79424 130052
rect 79464 130012 79506 130052
rect 79546 130012 79588 130052
rect 79628 130012 79670 130052
rect 79710 130012 79752 130052
rect 79792 130012 94544 130052
rect 94584 130012 94626 130052
rect 94666 130012 94708 130052
rect 94748 130012 94790 130052
rect 94830 130012 94872 130052
rect 94912 130012 109664 130052
rect 109704 130012 109746 130052
rect 109786 130012 109828 130052
rect 109868 130012 109910 130052
rect 109950 130012 109992 130052
rect 110032 130012 124784 130052
rect 124824 130012 124866 130052
rect 124906 130012 124948 130052
rect 124988 130012 125030 130052
rect 125070 130012 125112 130052
rect 125152 130012 139904 130052
rect 139944 130012 139986 130052
rect 140026 130012 140068 130052
rect 140108 130012 140150 130052
rect 140190 130012 140232 130052
rect 140272 130012 148320 130052
rect 75648 129988 148320 130012
rect 96835 129884 96893 129885
rect 96835 129844 96844 129884
rect 96884 129844 96893 129884
rect 96835 129843 96893 129844
rect 97227 129884 97269 129893
rect 97227 129844 97228 129884
rect 97268 129844 97269 129884
rect 97227 129835 97269 129844
rect 103179 129884 103221 129893
rect 103179 129844 103180 129884
rect 103220 129844 103221 129884
rect 103179 129835 103221 129844
rect 105955 129884 106013 129885
rect 105955 129844 105964 129884
rect 106004 129844 106013 129884
rect 105955 129843 106013 129844
rect 103563 129800 103605 129809
rect 103563 129760 103564 129800
rect 103604 129760 103605 129800
rect 103563 129751 103605 129760
rect 96163 129716 96221 129717
rect 96163 129676 96172 129716
rect 96212 129676 96221 129716
rect 96163 129675 96221 129676
rect 97131 129716 97173 129725
rect 97131 129676 97132 129716
rect 97172 129676 97173 129716
rect 97131 129667 97173 129676
rect 97323 129716 97365 129725
rect 97323 129676 97324 129716
rect 97364 129676 97365 129716
rect 97323 129667 97365 129676
rect 97419 129716 97461 129725
rect 97419 129676 97420 129716
rect 97460 129676 97461 129716
rect 97419 129667 97461 129676
rect 103083 129716 103125 129725
rect 103083 129676 103084 129716
rect 103124 129676 103125 129716
rect 103083 129667 103125 129676
rect 103275 129716 103317 129725
rect 103275 129676 103276 129716
rect 103316 129676 103317 129716
rect 103275 129667 103317 129676
rect 103939 129716 103997 129717
rect 103939 129676 103948 129716
rect 103988 129676 103997 129716
rect 103939 129675 103997 129676
rect 104803 129716 104861 129717
rect 104803 129676 104812 129716
rect 104852 129676 104861 129716
rect 104803 129675 104861 129676
rect 110563 129716 110621 129717
rect 110563 129676 110572 129716
rect 110612 129676 110621 129716
rect 110563 129675 110621 129676
rect 112011 129716 112053 129725
rect 112011 129676 112012 129716
rect 112052 129676 112053 129716
rect 112011 129667 112053 129676
rect 113923 129716 113981 129717
rect 113923 129676 113932 129716
rect 113972 129676 113981 129716
rect 113923 129675 113981 129676
rect 115371 129716 115413 129725
rect 115371 129676 115372 129716
rect 115412 129676 115413 129716
rect 115371 129667 115413 129676
rect 75648 129296 148320 129320
rect 75648 129256 78184 129296
rect 78224 129256 78266 129296
rect 78306 129256 78348 129296
rect 78388 129256 78430 129296
rect 78470 129256 78512 129296
rect 78552 129256 93304 129296
rect 93344 129256 93386 129296
rect 93426 129256 93468 129296
rect 93508 129256 93550 129296
rect 93590 129256 93632 129296
rect 93672 129256 108424 129296
rect 108464 129256 108506 129296
rect 108546 129256 108588 129296
rect 108628 129256 108670 129296
rect 108710 129256 108752 129296
rect 108792 129256 123544 129296
rect 123584 129256 123626 129296
rect 123666 129256 123708 129296
rect 123748 129256 123790 129296
rect 123830 129256 123872 129296
rect 123912 129256 138664 129296
rect 138704 129256 138746 129296
rect 138786 129256 138828 129296
rect 138868 129256 138910 129296
rect 138950 129256 138992 129296
rect 139032 129256 148320 129296
rect 75648 129232 148320 129256
rect 94155 129128 94197 129137
rect 94155 129088 94156 129128
rect 94196 129088 94197 129128
rect 94155 129079 94197 129088
rect 96739 129128 96797 129129
rect 96739 129088 96748 129128
rect 96788 129088 96797 129128
rect 96739 129087 96797 129088
rect 104043 129044 104085 129053
rect 104043 129004 104044 129044
rect 104084 129004 104085 129044
rect 104043 128995 104085 129004
rect 121227 129044 121269 129053
rect 121227 129004 121228 129044
rect 121268 129004 121269 129044
rect 121227 128995 121269 129004
rect 93867 128876 93909 128885
rect 93867 128836 93868 128876
rect 93908 128836 93909 128876
rect 93867 128827 93909 128836
rect 93963 128876 94005 128885
rect 93963 128836 93964 128876
rect 94004 128836 94005 128876
rect 93963 128827 94005 128836
rect 96067 128876 96125 128877
rect 96067 128836 96076 128876
rect 96116 128836 96125 128876
rect 96067 128835 96125 128836
rect 119491 128876 119549 128877
rect 119491 128836 119500 128876
rect 119540 128836 119549 128876
rect 119491 128835 119549 128836
rect 120355 128876 120413 128877
rect 120355 128836 120364 128876
rect 120404 128836 120413 128876
rect 120355 128835 120413 128836
rect 121987 128876 122045 128877
rect 121987 128836 121996 128876
rect 122036 128836 122045 128876
rect 121987 128835 122045 128836
rect 94051 128792 94109 128793
rect 94051 128752 94060 128792
rect 94100 128752 94109 128792
rect 94051 128751 94109 128752
rect 94147 128708 94205 128709
rect 94147 128668 94156 128708
rect 94196 128668 94205 128708
rect 94147 128667 94205 128668
rect 120163 128708 120221 128709
rect 120163 128668 120172 128708
rect 120212 128668 120221 128708
rect 120163 128667 120221 128668
rect 121027 128708 121085 128709
rect 121027 128668 121036 128708
rect 121076 128668 121085 128708
rect 121027 128667 121085 128668
rect 121899 128708 121941 128717
rect 121899 128668 121900 128708
rect 121940 128668 121941 128708
rect 121899 128659 121941 128668
rect 75648 128540 148320 128564
rect 75648 128500 79424 128540
rect 79464 128500 79506 128540
rect 79546 128500 79588 128540
rect 79628 128500 79670 128540
rect 79710 128500 79752 128540
rect 79792 128500 94544 128540
rect 94584 128500 94626 128540
rect 94666 128500 94708 128540
rect 94748 128500 94790 128540
rect 94830 128500 94872 128540
rect 94912 128500 109664 128540
rect 109704 128500 109746 128540
rect 109786 128500 109828 128540
rect 109868 128500 109910 128540
rect 109950 128500 109992 128540
rect 110032 128500 124784 128540
rect 124824 128500 124866 128540
rect 124906 128500 124948 128540
rect 124988 128500 125030 128540
rect 125070 128500 125112 128540
rect 125152 128500 139904 128540
rect 139944 128500 139986 128540
rect 140026 128500 140068 128540
rect 140108 128500 140150 128540
rect 140190 128500 140232 128540
rect 140272 128500 148320 128540
rect 75648 128476 148320 128500
rect 99147 128372 99189 128381
rect 99147 128332 99148 128372
rect 99188 128332 99189 128372
rect 99147 128323 99189 128332
rect 119299 128372 119357 128373
rect 119299 128332 119308 128372
rect 119348 128332 119357 128372
rect 119299 128331 119357 128332
rect 119779 128372 119837 128373
rect 119779 128332 119788 128372
rect 119828 128332 119837 128372
rect 119779 128331 119837 128332
rect 123139 128372 123197 128373
rect 123139 128332 123148 128372
rect 123188 128332 123197 128372
rect 123139 128331 123197 128332
rect 120747 128288 120789 128297
rect 120747 128248 120748 128288
rect 120788 128248 120789 128288
rect 120747 128239 120789 128248
rect 99147 128204 99189 128213
rect 99147 128164 99148 128204
rect 99188 128164 99189 128204
rect 99147 128155 99189 128164
rect 99235 128204 99293 128205
rect 99235 128164 99244 128204
rect 99284 128164 99293 128204
rect 99235 128163 99293 128164
rect 118243 128204 118301 128205
rect 118243 128164 118252 128204
rect 118292 128164 118301 128204
rect 118243 128163 118301 128164
rect 118443 128202 118485 128211
rect 118443 128162 118444 128202
rect 118484 128162 118485 128202
rect 118531 128204 118589 128205
rect 118531 128164 118540 128204
rect 118580 128164 118589 128204
rect 118531 128163 118589 128164
rect 118627 128204 118685 128205
rect 118627 128164 118636 128204
rect 118676 128164 118685 128204
rect 118627 128163 118685 128164
rect 119019 128204 119061 128213
rect 119019 128164 119020 128204
rect 119060 128164 119061 128204
rect 118443 128153 118485 128162
rect 119019 128155 119061 128164
rect 119115 128204 119157 128213
rect 119115 128164 119116 128204
rect 119156 128164 119157 128204
rect 119115 128155 119157 128164
rect 119211 128204 119253 128213
rect 119211 128164 119212 128204
rect 119252 128164 119253 128204
rect 119211 128155 119253 128164
rect 119587 128204 119645 128205
rect 119587 128164 119596 128204
rect 119636 128164 119645 128204
rect 119587 128163 119645 128164
rect 119691 128204 119733 128213
rect 119691 128164 119692 128204
rect 119732 128164 119733 128204
rect 119691 128155 119733 128164
rect 119883 128204 119925 128213
rect 119883 128164 119884 128204
rect 119924 128164 119925 128204
rect 119883 128155 119925 128164
rect 121123 128204 121181 128205
rect 121123 128164 121132 128204
rect 121172 128164 121181 128204
rect 121123 128163 121181 128164
rect 121987 128204 122045 128205
rect 121987 128164 121996 128204
rect 122036 128164 122045 128204
rect 121987 128163 122045 128164
rect 99051 128120 99093 128129
rect 99051 128080 99052 128120
rect 99092 128080 99093 128120
rect 99051 128071 99093 128080
rect 98955 128036 98997 128045
rect 98955 127996 98956 128036
rect 98996 127996 98997 128036
rect 98955 127987 98997 127996
rect 118827 127952 118869 127961
rect 118827 127912 118828 127952
rect 118868 127912 118869 127952
rect 118827 127903 118869 127912
rect 123139 127952 123197 127953
rect 123139 127912 123148 127952
rect 123188 127912 123197 127952
rect 123139 127911 123197 127912
rect 75648 127784 148320 127808
rect 75648 127744 78184 127784
rect 78224 127744 78266 127784
rect 78306 127744 78348 127784
rect 78388 127744 78430 127784
rect 78470 127744 78512 127784
rect 78552 127744 93304 127784
rect 93344 127744 93386 127784
rect 93426 127744 93468 127784
rect 93508 127744 93550 127784
rect 93590 127744 93632 127784
rect 93672 127744 108424 127784
rect 108464 127744 108506 127784
rect 108546 127744 108588 127784
rect 108628 127744 108670 127784
rect 108710 127744 108752 127784
rect 108792 127744 123544 127784
rect 123584 127744 123626 127784
rect 123666 127744 123708 127784
rect 123748 127744 123790 127784
rect 123830 127744 123872 127784
rect 123912 127744 138664 127784
rect 138704 127744 138746 127784
rect 138786 127744 138828 127784
rect 138868 127744 138910 127784
rect 138950 127744 138992 127784
rect 139032 127744 148320 127784
rect 75648 127720 148320 127744
rect 94827 127616 94869 127625
rect 94827 127576 94828 127616
rect 94868 127576 94869 127616
rect 94827 127567 94869 127576
rect 94598 127364 94640 127373
rect 94598 127324 94599 127364
rect 94639 127324 94640 127364
rect 94598 127315 94640 127324
rect 94703 127364 94761 127365
rect 94703 127324 94712 127364
rect 94752 127324 94761 127364
rect 94703 127323 94761 127324
rect 94827 127364 94869 127373
rect 94827 127324 94828 127364
rect 94868 127324 94869 127364
rect 94827 127315 94869 127324
rect 94923 127364 94965 127373
rect 94923 127324 94924 127364
rect 94964 127324 94965 127364
rect 94923 127315 94965 127324
rect 118827 127364 118869 127373
rect 118827 127324 118828 127364
rect 118868 127324 118869 127364
rect 118827 127315 118869 127324
rect 118923 127364 118965 127373
rect 118923 127324 118924 127364
rect 118964 127324 118965 127364
rect 118923 127315 118965 127324
rect 119019 127364 119061 127373
rect 119019 127324 119020 127364
rect 119060 127324 119061 127364
rect 119019 127315 119061 127324
rect 119107 127196 119165 127197
rect 119107 127156 119116 127196
rect 119156 127156 119165 127196
rect 119107 127155 119165 127156
rect 75648 127028 148320 127052
rect 75648 126988 79424 127028
rect 79464 126988 79506 127028
rect 79546 126988 79588 127028
rect 79628 126988 79670 127028
rect 79710 126988 79752 127028
rect 79792 126988 94544 127028
rect 94584 126988 94626 127028
rect 94666 126988 94708 127028
rect 94748 126988 94790 127028
rect 94830 126988 94872 127028
rect 94912 126988 109664 127028
rect 109704 126988 109746 127028
rect 109786 126988 109828 127028
rect 109868 126988 109910 127028
rect 109950 126988 109992 127028
rect 110032 126988 124784 127028
rect 124824 126988 124866 127028
rect 124906 126988 124948 127028
rect 124988 126988 125030 127028
rect 125070 126988 125112 127028
rect 125152 126988 139904 127028
rect 139944 126988 139986 127028
rect 140026 126988 140068 127028
rect 140108 126988 140150 127028
rect 140190 126988 140232 127028
rect 140272 126988 148320 127028
rect 75648 126964 148320 126988
rect 94627 126860 94685 126861
rect 94627 126820 94636 126860
rect 94676 126820 94685 126860
rect 94627 126819 94685 126820
rect 95499 126860 95541 126869
rect 95499 126820 95500 126860
rect 95540 126820 95541 126860
rect 95499 126811 95541 126820
rect 94723 126776 94781 126777
rect 94723 126736 94732 126776
rect 94772 126736 94781 126776
rect 94723 126735 94781 126736
rect 94827 126692 94869 126701
rect 94827 126652 94828 126692
rect 94868 126652 94869 126692
rect 94827 126643 94869 126652
rect 94923 126692 94965 126701
rect 94923 126652 94924 126692
rect 94964 126652 94965 126692
rect 94923 126643 94965 126652
rect 95558 126692 95600 126701
rect 95558 126652 95559 126692
rect 95599 126652 95600 126692
rect 95558 126643 95600 126652
rect 95663 126692 95721 126693
rect 95663 126652 95672 126692
rect 95712 126652 95721 126692
rect 95663 126651 95721 126652
rect 95787 126692 95829 126701
rect 95787 126652 95788 126692
rect 95828 126652 95829 126692
rect 95787 126643 95829 126652
rect 95883 126692 95925 126701
rect 95883 126652 95884 126692
rect 95924 126652 95925 126692
rect 95883 126643 95925 126652
rect 94827 126440 94869 126449
rect 94827 126400 94828 126440
rect 94868 126400 94869 126440
rect 94827 126391 94869 126400
rect 75648 126272 148320 126296
rect 75648 126232 78184 126272
rect 78224 126232 78266 126272
rect 78306 126232 78348 126272
rect 78388 126232 78430 126272
rect 78470 126232 78512 126272
rect 78552 126232 93304 126272
rect 93344 126232 93386 126272
rect 93426 126232 93468 126272
rect 93508 126232 93550 126272
rect 93590 126232 93632 126272
rect 93672 126232 108424 126272
rect 108464 126232 108506 126272
rect 108546 126232 108588 126272
rect 108628 126232 108670 126272
rect 108710 126232 108752 126272
rect 108792 126232 123544 126272
rect 123584 126232 123626 126272
rect 123666 126232 123708 126272
rect 123748 126232 123790 126272
rect 123830 126232 123872 126272
rect 123912 126232 138664 126272
rect 138704 126232 138746 126272
rect 138786 126232 138828 126272
rect 138868 126232 138910 126272
rect 138950 126232 138992 126272
rect 139032 126232 148320 126272
rect 75648 126208 148320 126232
rect 119211 125877 119253 125886
rect 119115 125852 119157 125861
rect 119115 125812 119116 125852
rect 119156 125812 119157 125852
rect 119211 125837 119212 125877
rect 119252 125837 119253 125877
rect 119211 125828 119253 125837
rect 119115 125803 119157 125812
rect 119395 125768 119453 125769
rect 119395 125728 119404 125768
rect 119444 125728 119453 125768
rect 119395 125727 119453 125728
rect 119107 125684 119165 125685
rect 119107 125644 119116 125684
rect 119156 125644 119165 125684
rect 119107 125643 119165 125644
rect 75648 125516 148320 125540
rect 75648 125476 79424 125516
rect 79464 125476 79506 125516
rect 79546 125476 79588 125516
rect 79628 125476 79670 125516
rect 79710 125476 79752 125516
rect 79792 125476 94544 125516
rect 94584 125476 94626 125516
rect 94666 125476 94708 125516
rect 94748 125476 94790 125516
rect 94830 125476 94872 125516
rect 94912 125476 109664 125516
rect 109704 125476 109746 125516
rect 109786 125476 109828 125516
rect 109868 125476 109910 125516
rect 109950 125476 109992 125516
rect 110032 125476 124784 125516
rect 124824 125476 124866 125516
rect 124906 125476 124948 125516
rect 124988 125476 125030 125516
rect 125070 125476 125112 125516
rect 125152 125476 139904 125516
rect 139944 125476 139986 125516
rect 140026 125476 140068 125516
rect 140108 125476 140150 125516
rect 140190 125476 140232 125516
rect 140272 125476 148320 125516
rect 75648 125452 148320 125476
rect 121035 125348 121077 125357
rect 121035 125308 121036 125348
rect 121076 125308 121077 125348
rect 121035 125299 121077 125308
rect 121123 125180 121181 125181
rect 121123 125140 121132 125180
rect 121172 125140 121181 125180
rect 121123 125139 121181 125140
rect 121515 125180 121557 125189
rect 121515 125140 121516 125180
rect 121556 125140 121557 125180
rect 121515 125131 121557 125140
rect 122179 125180 122237 125181
rect 122179 125140 122188 125180
rect 122228 125140 122237 125180
rect 122179 125139 122237 125140
rect 75648 124760 148320 124784
rect 75648 124720 78184 124760
rect 78224 124720 78266 124760
rect 78306 124720 78348 124760
rect 78388 124720 78430 124760
rect 78470 124720 78512 124760
rect 78552 124720 93304 124760
rect 93344 124720 93386 124760
rect 93426 124720 93468 124760
rect 93508 124720 93550 124760
rect 93590 124720 93632 124760
rect 93672 124720 108424 124760
rect 108464 124720 108506 124760
rect 108546 124720 108588 124760
rect 108628 124720 108670 124760
rect 108710 124720 108752 124760
rect 108792 124720 123544 124760
rect 123584 124720 123626 124760
rect 123666 124720 123708 124760
rect 123748 124720 123790 124760
rect 123830 124720 123872 124760
rect 123912 124720 138664 124760
rect 138704 124720 138746 124760
rect 138786 124720 138828 124760
rect 138868 124720 138910 124760
rect 138950 124720 138992 124760
rect 139032 124720 148320 124760
rect 75648 124696 148320 124720
rect 79555 124592 79613 124593
rect 79555 124552 79564 124592
rect 79604 124552 79613 124592
rect 79555 124551 79613 124552
rect 78883 124340 78941 124341
rect 78883 124300 78892 124340
rect 78932 124300 78941 124340
rect 78883 124299 78941 124300
rect 75648 124004 148320 124028
rect 75648 123964 79424 124004
rect 79464 123964 79506 124004
rect 79546 123964 79588 124004
rect 79628 123964 79670 124004
rect 79710 123964 79752 124004
rect 79792 123964 94544 124004
rect 94584 123964 94626 124004
rect 94666 123964 94708 124004
rect 94748 123964 94790 124004
rect 94830 123964 94872 124004
rect 94912 123964 109664 124004
rect 109704 123964 109746 124004
rect 109786 123964 109828 124004
rect 109868 123964 109910 124004
rect 109950 123964 109992 124004
rect 110032 123964 124784 124004
rect 124824 123964 124866 124004
rect 124906 123964 124948 124004
rect 124988 123964 125030 124004
rect 125070 123964 125112 124004
rect 125152 123964 139904 124004
rect 139944 123964 139986 124004
rect 140026 123964 140068 124004
rect 140108 123964 140150 124004
rect 140190 123964 140232 124004
rect 140272 123964 148320 124004
rect 75648 123940 148320 123964
rect 121603 123836 121661 123837
rect 121603 123796 121612 123836
rect 121652 123796 121661 123836
rect 121603 123795 121661 123796
rect 119211 123752 119253 123761
rect 119211 123712 119212 123752
rect 119252 123712 119253 123752
rect 119211 123703 119253 123712
rect 119587 123668 119645 123669
rect 119587 123628 119596 123668
rect 119636 123628 119645 123668
rect 119587 123627 119645 123628
rect 120451 123668 120509 123669
rect 120451 123628 120460 123668
rect 120500 123628 120509 123668
rect 120451 123627 120509 123628
rect 121603 123416 121661 123417
rect 121603 123376 121612 123416
rect 121652 123376 121661 123416
rect 121603 123375 121661 123376
rect 75648 123248 148320 123272
rect 75648 123208 78184 123248
rect 78224 123208 78266 123248
rect 78306 123208 78348 123248
rect 78388 123208 78430 123248
rect 78470 123208 78512 123248
rect 78552 123208 93304 123248
rect 93344 123208 93386 123248
rect 93426 123208 93468 123248
rect 93508 123208 93550 123248
rect 93590 123208 93632 123248
rect 93672 123208 108424 123248
rect 108464 123208 108506 123248
rect 108546 123208 108588 123248
rect 108628 123208 108670 123248
rect 108710 123208 108752 123248
rect 108792 123208 123544 123248
rect 123584 123208 123626 123248
rect 123666 123208 123708 123248
rect 123748 123208 123790 123248
rect 123830 123208 123872 123248
rect 123912 123208 138664 123248
rect 138704 123208 138746 123248
rect 138786 123208 138828 123248
rect 138868 123208 138910 123248
rect 138950 123208 138992 123248
rect 139032 123208 148320 123248
rect 75648 123184 148320 123208
rect 119691 122996 119733 123005
rect 119691 122956 119692 122996
rect 119732 122956 119733 122996
rect 119691 122947 119733 122956
rect 75648 122492 148320 122516
rect 75648 122452 79424 122492
rect 79464 122452 79506 122492
rect 79546 122452 79588 122492
rect 79628 122452 79670 122492
rect 79710 122452 79752 122492
rect 79792 122452 94544 122492
rect 94584 122452 94626 122492
rect 94666 122452 94708 122492
rect 94748 122452 94790 122492
rect 94830 122452 94872 122492
rect 94912 122452 109664 122492
rect 109704 122452 109746 122492
rect 109786 122452 109828 122492
rect 109868 122452 109910 122492
rect 109950 122452 109992 122492
rect 110032 122452 124784 122492
rect 124824 122452 124866 122492
rect 124906 122452 124948 122492
rect 124988 122452 125030 122492
rect 125070 122452 125112 122492
rect 125152 122452 139904 122492
rect 139944 122452 139986 122492
rect 140026 122452 140068 122492
rect 140108 122452 140150 122492
rect 140190 122452 140232 122492
rect 140272 122452 148320 122492
rect 75648 122428 148320 122452
rect 75648 121736 148320 121760
rect 75648 121696 78184 121736
rect 78224 121696 78266 121736
rect 78306 121696 78348 121736
rect 78388 121696 78430 121736
rect 78470 121696 78512 121736
rect 78552 121696 93304 121736
rect 93344 121696 93386 121736
rect 93426 121696 93468 121736
rect 93508 121696 93550 121736
rect 93590 121696 93632 121736
rect 93672 121696 108424 121736
rect 108464 121696 108506 121736
rect 108546 121696 108588 121736
rect 108628 121696 108670 121736
rect 108710 121696 108752 121736
rect 108792 121696 123544 121736
rect 123584 121696 123626 121736
rect 123666 121696 123708 121736
rect 123748 121696 123790 121736
rect 123830 121696 123872 121736
rect 123912 121696 138664 121736
rect 138704 121696 138746 121736
rect 138786 121696 138828 121736
rect 138868 121696 138910 121736
rect 138950 121696 138992 121736
rect 139032 121696 148320 121736
rect 75648 121672 148320 121696
rect 75648 120980 148320 121004
rect 75648 120940 79424 120980
rect 79464 120940 79506 120980
rect 79546 120940 79588 120980
rect 79628 120940 79670 120980
rect 79710 120940 79752 120980
rect 79792 120940 94544 120980
rect 94584 120940 94626 120980
rect 94666 120940 94708 120980
rect 94748 120940 94790 120980
rect 94830 120940 94872 120980
rect 94912 120940 109664 120980
rect 109704 120940 109746 120980
rect 109786 120940 109828 120980
rect 109868 120940 109910 120980
rect 109950 120940 109992 120980
rect 110032 120940 124784 120980
rect 124824 120940 124866 120980
rect 124906 120940 124948 120980
rect 124988 120940 125030 120980
rect 125070 120940 125112 120980
rect 125152 120940 139904 120980
rect 139944 120940 139986 120980
rect 140026 120940 140068 120980
rect 140108 120940 140150 120980
rect 140190 120940 140232 120980
rect 140272 120940 148320 120980
rect 75648 120916 148320 120940
rect 75648 120224 148320 120248
rect 75648 120184 78184 120224
rect 78224 120184 78266 120224
rect 78306 120184 78348 120224
rect 78388 120184 78430 120224
rect 78470 120184 78512 120224
rect 78552 120184 93304 120224
rect 93344 120184 93386 120224
rect 93426 120184 93468 120224
rect 93508 120184 93550 120224
rect 93590 120184 93632 120224
rect 93672 120184 108424 120224
rect 108464 120184 108506 120224
rect 108546 120184 108588 120224
rect 108628 120184 108670 120224
rect 108710 120184 108752 120224
rect 108792 120184 123544 120224
rect 123584 120184 123626 120224
rect 123666 120184 123708 120224
rect 123748 120184 123790 120224
rect 123830 120184 123872 120224
rect 123912 120184 138664 120224
rect 138704 120184 138746 120224
rect 138786 120184 138828 120224
rect 138868 120184 138910 120224
rect 138950 120184 138992 120224
rect 139032 120184 148320 120224
rect 75648 120160 148320 120184
rect 75648 119468 148320 119492
rect 75648 119428 79424 119468
rect 79464 119428 79506 119468
rect 79546 119428 79588 119468
rect 79628 119428 79670 119468
rect 79710 119428 79752 119468
rect 79792 119428 94544 119468
rect 94584 119428 94626 119468
rect 94666 119428 94708 119468
rect 94748 119428 94790 119468
rect 94830 119428 94872 119468
rect 94912 119428 109664 119468
rect 109704 119428 109746 119468
rect 109786 119428 109828 119468
rect 109868 119428 109910 119468
rect 109950 119428 109992 119468
rect 110032 119428 124784 119468
rect 124824 119428 124866 119468
rect 124906 119428 124948 119468
rect 124988 119428 125030 119468
rect 125070 119428 125112 119468
rect 125152 119428 139904 119468
rect 139944 119428 139986 119468
rect 140026 119428 140068 119468
rect 140108 119428 140150 119468
rect 140190 119428 140232 119468
rect 140272 119428 148320 119468
rect 75648 119404 148320 119428
rect 75648 118712 148320 118736
rect 75648 118672 78184 118712
rect 78224 118672 78266 118712
rect 78306 118672 78348 118712
rect 78388 118672 78430 118712
rect 78470 118672 78512 118712
rect 78552 118672 93304 118712
rect 93344 118672 93386 118712
rect 93426 118672 93468 118712
rect 93508 118672 93550 118712
rect 93590 118672 93632 118712
rect 93672 118672 108424 118712
rect 108464 118672 108506 118712
rect 108546 118672 108588 118712
rect 108628 118672 108670 118712
rect 108710 118672 108752 118712
rect 108792 118672 123544 118712
rect 123584 118672 123626 118712
rect 123666 118672 123708 118712
rect 123748 118672 123790 118712
rect 123830 118672 123872 118712
rect 123912 118672 138664 118712
rect 138704 118672 138746 118712
rect 138786 118672 138828 118712
rect 138868 118672 138910 118712
rect 138950 118672 138992 118712
rect 139032 118672 148320 118712
rect 75648 118648 148320 118672
rect 75648 117956 148320 117980
rect 75648 117916 79424 117956
rect 79464 117916 79506 117956
rect 79546 117916 79588 117956
rect 79628 117916 79670 117956
rect 79710 117916 79752 117956
rect 79792 117916 94544 117956
rect 94584 117916 94626 117956
rect 94666 117916 94708 117956
rect 94748 117916 94790 117956
rect 94830 117916 94872 117956
rect 94912 117916 109664 117956
rect 109704 117916 109746 117956
rect 109786 117916 109828 117956
rect 109868 117916 109910 117956
rect 109950 117916 109992 117956
rect 110032 117916 124784 117956
rect 124824 117916 124866 117956
rect 124906 117916 124948 117956
rect 124988 117916 125030 117956
rect 125070 117916 125112 117956
rect 125152 117916 139904 117956
rect 139944 117916 139986 117956
rect 140026 117916 140068 117956
rect 140108 117916 140150 117956
rect 140190 117916 140232 117956
rect 140272 117916 148320 117956
rect 75648 117892 148320 117916
rect 75648 117200 148320 117224
rect 75648 117160 78184 117200
rect 78224 117160 78266 117200
rect 78306 117160 78348 117200
rect 78388 117160 78430 117200
rect 78470 117160 78512 117200
rect 78552 117160 93304 117200
rect 93344 117160 93386 117200
rect 93426 117160 93468 117200
rect 93508 117160 93550 117200
rect 93590 117160 93632 117200
rect 93672 117160 108424 117200
rect 108464 117160 108506 117200
rect 108546 117160 108588 117200
rect 108628 117160 108670 117200
rect 108710 117160 108752 117200
rect 108792 117160 123544 117200
rect 123584 117160 123626 117200
rect 123666 117160 123708 117200
rect 123748 117160 123790 117200
rect 123830 117160 123872 117200
rect 123912 117160 138664 117200
rect 138704 117160 138746 117200
rect 138786 117160 138828 117200
rect 138868 117160 138910 117200
rect 138950 117160 138992 117200
rect 139032 117160 148320 117200
rect 75648 117136 148320 117160
rect 75648 116444 148320 116468
rect 75648 116404 79424 116444
rect 79464 116404 79506 116444
rect 79546 116404 79588 116444
rect 79628 116404 79670 116444
rect 79710 116404 79752 116444
rect 79792 116404 94544 116444
rect 94584 116404 94626 116444
rect 94666 116404 94708 116444
rect 94748 116404 94790 116444
rect 94830 116404 94872 116444
rect 94912 116404 109664 116444
rect 109704 116404 109746 116444
rect 109786 116404 109828 116444
rect 109868 116404 109910 116444
rect 109950 116404 109992 116444
rect 110032 116404 124784 116444
rect 124824 116404 124866 116444
rect 124906 116404 124948 116444
rect 124988 116404 125030 116444
rect 125070 116404 125112 116444
rect 125152 116404 139904 116444
rect 139944 116404 139986 116444
rect 140026 116404 140068 116444
rect 140108 116404 140150 116444
rect 140190 116404 140232 116444
rect 140272 116404 148320 116444
rect 75648 116380 148320 116404
rect 75648 115688 148320 115712
rect 75648 115648 78184 115688
rect 78224 115648 78266 115688
rect 78306 115648 78348 115688
rect 78388 115648 78430 115688
rect 78470 115648 78512 115688
rect 78552 115648 93304 115688
rect 93344 115648 93386 115688
rect 93426 115648 93468 115688
rect 93508 115648 93550 115688
rect 93590 115648 93632 115688
rect 93672 115648 108424 115688
rect 108464 115648 108506 115688
rect 108546 115648 108588 115688
rect 108628 115648 108670 115688
rect 108710 115648 108752 115688
rect 108792 115648 123544 115688
rect 123584 115648 123626 115688
rect 123666 115648 123708 115688
rect 123748 115648 123790 115688
rect 123830 115648 123872 115688
rect 123912 115648 138664 115688
rect 138704 115648 138746 115688
rect 138786 115648 138828 115688
rect 138868 115648 138910 115688
rect 138950 115648 138992 115688
rect 139032 115648 148320 115688
rect 75648 115624 148320 115648
rect 75648 114932 148320 114956
rect 75648 114892 79424 114932
rect 79464 114892 79506 114932
rect 79546 114892 79588 114932
rect 79628 114892 79670 114932
rect 79710 114892 79752 114932
rect 79792 114892 94544 114932
rect 94584 114892 94626 114932
rect 94666 114892 94708 114932
rect 94748 114892 94790 114932
rect 94830 114892 94872 114932
rect 94912 114892 109664 114932
rect 109704 114892 109746 114932
rect 109786 114892 109828 114932
rect 109868 114892 109910 114932
rect 109950 114892 109992 114932
rect 110032 114892 124784 114932
rect 124824 114892 124866 114932
rect 124906 114892 124948 114932
rect 124988 114892 125030 114932
rect 125070 114892 125112 114932
rect 125152 114892 139904 114932
rect 139944 114892 139986 114932
rect 140026 114892 140068 114932
rect 140108 114892 140150 114932
rect 140190 114892 140232 114932
rect 140272 114892 148320 114932
rect 75648 114868 148320 114892
rect 75648 114176 148320 114200
rect 75648 114136 78184 114176
rect 78224 114136 78266 114176
rect 78306 114136 78348 114176
rect 78388 114136 78430 114176
rect 78470 114136 78512 114176
rect 78552 114136 93304 114176
rect 93344 114136 93386 114176
rect 93426 114136 93468 114176
rect 93508 114136 93550 114176
rect 93590 114136 93632 114176
rect 93672 114136 108424 114176
rect 108464 114136 108506 114176
rect 108546 114136 108588 114176
rect 108628 114136 108670 114176
rect 108710 114136 108752 114176
rect 108792 114136 123544 114176
rect 123584 114136 123626 114176
rect 123666 114136 123708 114176
rect 123748 114136 123790 114176
rect 123830 114136 123872 114176
rect 123912 114136 138664 114176
rect 138704 114136 138746 114176
rect 138786 114136 138828 114176
rect 138868 114136 138910 114176
rect 138950 114136 138992 114176
rect 139032 114136 148320 114176
rect 75648 114112 148320 114136
rect 75648 113420 148320 113444
rect 75648 113380 79424 113420
rect 79464 113380 79506 113420
rect 79546 113380 79588 113420
rect 79628 113380 79670 113420
rect 79710 113380 79752 113420
rect 79792 113380 94544 113420
rect 94584 113380 94626 113420
rect 94666 113380 94708 113420
rect 94748 113380 94790 113420
rect 94830 113380 94872 113420
rect 94912 113380 109664 113420
rect 109704 113380 109746 113420
rect 109786 113380 109828 113420
rect 109868 113380 109910 113420
rect 109950 113380 109992 113420
rect 110032 113380 124784 113420
rect 124824 113380 124866 113420
rect 124906 113380 124948 113420
rect 124988 113380 125030 113420
rect 125070 113380 125112 113420
rect 125152 113380 139904 113420
rect 139944 113380 139986 113420
rect 140026 113380 140068 113420
rect 140108 113380 140150 113420
rect 140190 113380 140232 113420
rect 140272 113380 148320 113420
rect 75648 113356 148320 113380
rect 75648 112664 148320 112688
rect 75648 112624 78184 112664
rect 78224 112624 78266 112664
rect 78306 112624 78348 112664
rect 78388 112624 78430 112664
rect 78470 112624 78512 112664
rect 78552 112624 93304 112664
rect 93344 112624 93386 112664
rect 93426 112624 93468 112664
rect 93508 112624 93550 112664
rect 93590 112624 93632 112664
rect 93672 112624 108424 112664
rect 108464 112624 108506 112664
rect 108546 112624 108588 112664
rect 108628 112624 108670 112664
rect 108710 112624 108752 112664
rect 108792 112624 123544 112664
rect 123584 112624 123626 112664
rect 123666 112624 123708 112664
rect 123748 112624 123790 112664
rect 123830 112624 123872 112664
rect 123912 112624 138664 112664
rect 138704 112624 138746 112664
rect 138786 112624 138828 112664
rect 138868 112624 138910 112664
rect 138950 112624 138992 112664
rect 139032 112624 148320 112664
rect 75648 112600 148320 112624
rect 75648 111908 148320 111932
rect 75648 111868 79424 111908
rect 79464 111868 79506 111908
rect 79546 111868 79588 111908
rect 79628 111868 79670 111908
rect 79710 111868 79752 111908
rect 79792 111868 94544 111908
rect 94584 111868 94626 111908
rect 94666 111868 94708 111908
rect 94748 111868 94790 111908
rect 94830 111868 94872 111908
rect 94912 111868 109664 111908
rect 109704 111868 109746 111908
rect 109786 111868 109828 111908
rect 109868 111868 109910 111908
rect 109950 111868 109992 111908
rect 110032 111868 124784 111908
rect 124824 111868 124866 111908
rect 124906 111868 124948 111908
rect 124988 111868 125030 111908
rect 125070 111868 125112 111908
rect 125152 111868 139904 111908
rect 139944 111868 139986 111908
rect 140026 111868 140068 111908
rect 140108 111868 140150 111908
rect 140190 111868 140232 111908
rect 140272 111868 148320 111908
rect 75648 111844 148320 111868
rect 75648 111152 148320 111176
rect 75648 111112 78184 111152
rect 78224 111112 78266 111152
rect 78306 111112 78348 111152
rect 78388 111112 78430 111152
rect 78470 111112 78512 111152
rect 78552 111112 93304 111152
rect 93344 111112 93386 111152
rect 93426 111112 93468 111152
rect 93508 111112 93550 111152
rect 93590 111112 93632 111152
rect 93672 111112 108424 111152
rect 108464 111112 108506 111152
rect 108546 111112 108588 111152
rect 108628 111112 108670 111152
rect 108710 111112 108752 111152
rect 108792 111112 123544 111152
rect 123584 111112 123626 111152
rect 123666 111112 123708 111152
rect 123748 111112 123790 111152
rect 123830 111112 123872 111152
rect 123912 111112 138664 111152
rect 138704 111112 138746 111152
rect 138786 111112 138828 111152
rect 138868 111112 138910 111152
rect 138950 111112 138992 111152
rect 139032 111112 148320 111152
rect 75648 111088 148320 111112
rect 75648 110396 148320 110420
rect 75648 110356 79424 110396
rect 79464 110356 79506 110396
rect 79546 110356 79588 110396
rect 79628 110356 79670 110396
rect 79710 110356 79752 110396
rect 79792 110356 94544 110396
rect 94584 110356 94626 110396
rect 94666 110356 94708 110396
rect 94748 110356 94790 110396
rect 94830 110356 94872 110396
rect 94912 110356 109664 110396
rect 109704 110356 109746 110396
rect 109786 110356 109828 110396
rect 109868 110356 109910 110396
rect 109950 110356 109992 110396
rect 110032 110356 124784 110396
rect 124824 110356 124866 110396
rect 124906 110356 124948 110396
rect 124988 110356 125030 110396
rect 125070 110356 125112 110396
rect 125152 110356 139904 110396
rect 139944 110356 139986 110396
rect 140026 110356 140068 110396
rect 140108 110356 140150 110396
rect 140190 110356 140232 110396
rect 140272 110356 148320 110396
rect 75648 110332 148320 110356
rect 75648 109640 148320 109664
rect 75648 109600 78184 109640
rect 78224 109600 78266 109640
rect 78306 109600 78348 109640
rect 78388 109600 78430 109640
rect 78470 109600 78512 109640
rect 78552 109600 93304 109640
rect 93344 109600 93386 109640
rect 93426 109600 93468 109640
rect 93508 109600 93550 109640
rect 93590 109600 93632 109640
rect 93672 109600 108424 109640
rect 108464 109600 108506 109640
rect 108546 109600 108588 109640
rect 108628 109600 108670 109640
rect 108710 109600 108752 109640
rect 108792 109600 123544 109640
rect 123584 109600 123626 109640
rect 123666 109600 123708 109640
rect 123748 109600 123790 109640
rect 123830 109600 123872 109640
rect 123912 109600 138664 109640
rect 138704 109600 138746 109640
rect 138786 109600 138828 109640
rect 138868 109600 138910 109640
rect 138950 109600 138992 109640
rect 139032 109600 148320 109640
rect 75648 109576 148320 109600
rect 75648 108884 148320 108908
rect 75648 108844 79424 108884
rect 79464 108844 79506 108884
rect 79546 108844 79588 108884
rect 79628 108844 79670 108884
rect 79710 108844 79752 108884
rect 79792 108844 94544 108884
rect 94584 108844 94626 108884
rect 94666 108844 94708 108884
rect 94748 108844 94790 108884
rect 94830 108844 94872 108884
rect 94912 108844 109664 108884
rect 109704 108844 109746 108884
rect 109786 108844 109828 108884
rect 109868 108844 109910 108884
rect 109950 108844 109992 108884
rect 110032 108844 124784 108884
rect 124824 108844 124866 108884
rect 124906 108844 124948 108884
rect 124988 108844 125030 108884
rect 125070 108844 125112 108884
rect 125152 108844 139904 108884
rect 139944 108844 139986 108884
rect 140026 108844 140068 108884
rect 140108 108844 140150 108884
rect 140190 108844 140232 108884
rect 140272 108844 148320 108884
rect 75648 108820 148320 108844
rect 75648 108128 148320 108152
rect 75648 108088 78184 108128
rect 78224 108088 78266 108128
rect 78306 108088 78348 108128
rect 78388 108088 78430 108128
rect 78470 108088 78512 108128
rect 78552 108088 93304 108128
rect 93344 108088 93386 108128
rect 93426 108088 93468 108128
rect 93508 108088 93550 108128
rect 93590 108088 93632 108128
rect 93672 108088 108424 108128
rect 108464 108088 108506 108128
rect 108546 108088 108588 108128
rect 108628 108088 108670 108128
rect 108710 108088 108752 108128
rect 108792 108088 123544 108128
rect 123584 108088 123626 108128
rect 123666 108088 123708 108128
rect 123748 108088 123790 108128
rect 123830 108088 123872 108128
rect 123912 108088 138664 108128
rect 138704 108088 138746 108128
rect 138786 108088 138828 108128
rect 138868 108088 138910 108128
rect 138950 108088 138992 108128
rect 139032 108088 148320 108128
rect 75648 108064 148320 108088
rect 75648 107372 148320 107396
rect 75648 107332 79424 107372
rect 79464 107332 79506 107372
rect 79546 107332 79588 107372
rect 79628 107332 79670 107372
rect 79710 107332 79752 107372
rect 79792 107332 94544 107372
rect 94584 107332 94626 107372
rect 94666 107332 94708 107372
rect 94748 107332 94790 107372
rect 94830 107332 94872 107372
rect 94912 107332 109664 107372
rect 109704 107332 109746 107372
rect 109786 107332 109828 107372
rect 109868 107332 109910 107372
rect 109950 107332 109992 107372
rect 110032 107332 124784 107372
rect 124824 107332 124866 107372
rect 124906 107332 124948 107372
rect 124988 107332 125030 107372
rect 125070 107332 125112 107372
rect 125152 107332 139904 107372
rect 139944 107332 139986 107372
rect 140026 107332 140068 107372
rect 140108 107332 140150 107372
rect 140190 107332 140232 107372
rect 140272 107332 148320 107372
rect 75648 107308 148320 107332
rect 75648 106616 148320 106640
rect 75648 106576 78184 106616
rect 78224 106576 78266 106616
rect 78306 106576 78348 106616
rect 78388 106576 78430 106616
rect 78470 106576 78512 106616
rect 78552 106576 93304 106616
rect 93344 106576 93386 106616
rect 93426 106576 93468 106616
rect 93508 106576 93550 106616
rect 93590 106576 93632 106616
rect 93672 106576 108424 106616
rect 108464 106576 108506 106616
rect 108546 106576 108588 106616
rect 108628 106576 108670 106616
rect 108710 106576 108752 106616
rect 108792 106576 123544 106616
rect 123584 106576 123626 106616
rect 123666 106576 123708 106616
rect 123748 106576 123790 106616
rect 123830 106576 123872 106616
rect 123912 106576 138664 106616
rect 138704 106576 138746 106616
rect 138786 106576 138828 106616
rect 138868 106576 138910 106616
rect 138950 106576 138992 106616
rect 139032 106576 148320 106616
rect 75648 106552 148320 106576
rect 75648 105860 148320 105884
rect 75648 105820 79424 105860
rect 79464 105820 79506 105860
rect 79546 105820 79588 105860
rect 79628 105820 79670 105860
rect 79710 105820 79752 105860
rect 79792 105820 94544 105860
rect 94584 105820 94626 105860
rect 94666 105820 94708 105860
rect 94748 105820 94790 105860
rect 94830 105820 94872 105860
rect 94912 105820 109664 105860
rect 109704 105820 109746 105860
rect 109786 105820 109828 105860
rect 109868 105820 109910 105860
rect 109950 105820 109992 105860
rect 110032 105820 124784 105860
rect 124824 105820 124866 105860
rect 124906 105820 124948 105860
rect 124988 105820 125030 105860
rect 125070 105820 125112 105860
rect 125152 105820 139904 105860
rect 139944 105820 139986 105860
rect 140026 105820 140068 105860
rect 140108 105820 140150 105860
rect 140190 105820 140232 105860
rect 140272 105820 148320 105860
rect 75648 105796 148320 105820
rect 75648 105104 148320 105128
rect 75648 105064 78184 105104
rect 78224 105064 78266 105104
rect 78306 105064 78348 105104
rect 78388 105064 78430 105104
rect 78470 105064 78512 105104
rect 78552 105064 93304 105104
rect 93344 105064 93386 105104
rect 93426 105064 93468 105104
rect 93508 105064 93550 105104
rect 93590 105064 93632 105104
rect 93672 105064 108424 105104
rect 108464 105064 108506 105104
rect 108546 105064 108588 105104
rect 108628 105064 108670 105104
rect 108710 105064 108752 105104
rect 108792 105064 123544 105104
rect 123584 105064 123626 105104
rect 123666 105064 123708 105104
rect 123748 105064 123790 105104
rect 123830 105064 123872 105104
rect 123912 105064 138664 105104
rect 138704 105064 138746 105104
rect 138786 105064 138828 105104
rect 138868 105064 138910 105104
rect 138950 105064 138992 105104
rect 139032 105064 148320 105104
rect 75648 105040 148320 105064
rect 75648 104348 148320 104372
rect 75648 104308 79424 104348
rect 79464 104308 79506 104348
rect 79546 104308 79588 104348
rect 79628 104308 79670 104348
rect 79710 104308 79752 104348
rect 79792 104308 94544 104348
rect 94584 104308 94626 104348
rect 94666 104308 94708 104348
rect 94748 104308 94790 104348
rect 94830 104308 94872 104348
rect 94912 104308 109664 104348
rect 109704 104308 109746 104348
rect 109786 104308 109828 104348
rect 109868 104308 109910 104348
rect 109950 104308 109992 104348
rect 110032 104308 124784 104348
rect 124824 104308 124866 104348
rect 124906 104308 124948 104348
rect 124988 104308 125030 104348
rect 125070 104308 125112 104348
rect 125152 104308 139904 104348
rect 139944 104308 139986 104348
rect 140026 104308 140068 104348
rect 140108 104308 140150 104348
rect 140190 104308 140232 104348
rect 140272 104308 148320 104348
rect 75648 104284 148320 104308
rect 75648 103592 148320 103616
rect 75648 103552 78184 103592
rect 78224 103552 78266 103592
rect 78306 103552 78348 103592
rect 78388 103552 78430 103592
rect 78470 103552 78512 103592
rect 78552 103552 93304 103592
rect 93344 103552 93386 103592
rect 93426 103552 93468 103592
rect 93508 103552 93550 103592
rect 93590 103552 93632 103592
rect 93672 103552 108424 103592
rect 108464 103552 108506 103592
rect 108546 103552 108588 103592
rect 108628 103552 108670 103592
rect 108710 103552 108752 103592
rect 108792 103552 123544 103592
rect 123584 103552 123626 103592
rect 123666 103552 123708 103592
rect 123748 103552 123790 103592
rect 123830 103552 123872 103592
rect 123912 103552 138664 103592
rect 138704 103552 138746 103592
rect 138786 103552 138828 103592
rect 138868 103552 138910 103592
rect 138950 103552 138992 103592
rect 139032 103552 148320 103592
rect 75648 103528 148320 103552
rect 75648 102836 148320 102860
rect 75648 102796 79424 102836
rect 79464 102796 79506 102836
rect 79546 102796 79588 102836
rect 79628 102796 79670 102836
rect 79710 102796 79752 102836
rect 79792 102796 94544 102836
rect 94584 102796 94626 102836
rect 94666 102796 94708 102836
rect 94748 102796 94790 102836
rect 94830 102796 94872 102836
rect 94912 102796 109664 102836
rect 109704 102796 109746 102836
rect 109786 102796 109828 102836
rect 109868 102796 109910 102836
rect 109950 102796 109992 102836
rect 110032 102796 124784 102836
rect 124824 102796 124866 102836
rect 124906 102796 124948 102836
rect 124988 102796 125030 102836
rect 125070 102796 125112 102836
rect 125152 102796 139904 102836
rect 139944 102796 139986 102836
rect 140026 102796 140068 102836
rect 140108 102796 140150 102836
rect 140190 102796 140232 102836
rect 140272 102796 148320 102836
rect 75648 102772 148320 102796
rect 75648 102080 148320 102104
rect 75648 102040 78184 102080
rect 78224 102040 78266 102080
rect 78306 102040 78348 102080
rect 78388 102040 78430 102080
rect 78470 102040 78512 102080
rect 78552 102040 93304 102080
rect 93344 102040 93386 102080
rect 93426 102040 93468 102080
rect 93508 102040 93550 102080
rect 93590 102040 93632 102080
rect 93672 102040 108424 102080
rect 108464 102040 108506 102080
rect 108546 102040 108588 102080
rect 108628 102040 108670 102080
rect 108710 102040 108752 102080
rect 108792 102040 123544 102080
rect 123584 102040 123626 102080
rect 123666 102040 123708 102080
rect 123748 102040 123790 102080
rect 123830 102040 123872 102080
rect 123912 102040 138664 102080
rect 138704 102040 138746 102080
rect 138786 102040 138828 102080
rect 138868 102040 138910 102080
rect 138950 102040 138992 102080
rect 139032 102040 148320 102080
rect 75648 102016 148320 102040
rect 75648 101324 148320 101348
rect 75648 101284 79424 101324
rect 79464 101284 79506 101324
rect 79546 101284 79588 101324
rect 79628 101284 79670 101324
rect 79710 101284 79752 101324
rect 79792 101284 94544 101324
rect 94584 101284 94626 101324
rect 94666 101284 94708 101324
rect 94748 101284 94790 101324
rect 94830 101284 94872 101324
rect 94912 101284 109664 101324
rect 109704 101284 109746 101324
rect 109786 101284 109828 101324
rect 109868 101284 109910 101324
rect 109950 101284 109992 101324
rect 110032 101284 124784 101324
rect 124824 101284 124866 101324
rect 124906 101284 124948 101324
rect 124988 101284 125030 101324
rect 125070 101284 125112 101324
rect 125152 101284 139904 101324
rect 139944 101284 139986 101324
rect 140026 101284 140068 101324
rect 140108 101284 140150 101324
rect 140190 101284 140232 101324
rect 140272 101284 148320 101324
rect 75648 101260 148320 101284
rect 75648 100568 148320 100592
rect 75648 100528 78184 100568
rect 78224 100528 78266 100568
rect 78306 100528 78348 100568
rect 78388 100528 78430 100568
rect 78470 100528 78512 100568
rect 78552 100528 93304 100568
rect 93344 100528 93386 100568
rect 93426 100528 93468 100568
rect 93508 100528 93550 100568
rect 93590 100528 93632 100568
rect 93672 100528 108424 100568
rect 108464 100528 108506 100568
rect 108546 100528 108588 100568
rect 108628 100528 108670 100568
rect 108710 100528 108752 100568
rect 108792 100528 123544 100568
rect 123584 100528 123626 100568
rect 123666 100528 123708 100568
rect 123748 100528 123790 100568
rect 123830 100528 123872 100568
rect 123912 100528 138664 100568
rect 138704 100528 138746 100568
rect 138786 100528 138828 100568
rect 138868 100528 138910 100568
rect 138950 100528 138992 100568
rect 139032 100528 148320 100568
rect 75648 100504 148320 100528
rect 75648 99812 148320 99836
rect 75648 99772 79424 99812
rect 79464 99772 79506 99812
rect 79546 99772 79588 99812
rect 79628 99772 79670 99812
rect 79710 99772 79752 99812
rect 79792 99772 94544 99812
rect 94584 99772 94626 99812
rect 94666 99772 94708 99812
rect 94748 99772 94790 99812
rect 94830 99772 94872 99812
rect 94912 99772 109664 99812
rect 109704 99772 109746 99812
rect 109786 99772 109828 99812
rect 109868 99772 109910 99812
rect 109950 99772 109992 99812
rect 110032 99772 124784 99812
rect 124824 99772 124866 99812
rect 124906 99772 124948 99812
rect 124988 99772 125030 99812
rect 125070 99772 125112 99812
rect 125152 99772 139904 99812
rect 139944 99772 139986 99812
rect 140026 99772 140068 99812
rect 140108 99772 140150 99812
rect 140190 99772 140232 99812
rect 140272 99772 148320 99812
rect 75648 99748 148320 99772
rect 75648 99056 148320 99080
rect 75648 99016 78184 99056
rect 78224 99016 78266 99056
rect 78306 99016 78348 99056
rect 78388 99016 78430 99056
rect 78470 99016 78512 99056
rect 78552 99016 93304 99056
rect 93344 99016 93386 99056
rect 93426 99016 93468 99056
rect 93508 99016 93550 99056
rect 93590 99016 93632 99056
rect 93672 99016 108424 99056
rect 108464 99016 108506 99056
rect 108546 99016 108588 99056
rect 108628 99016 108670 99056
rect 108710 99016 108752 99056
rect 108792 99016 123544 99056
rect 123584 99016 123626 99056
rect 123666 99016 123708 99056
rect 123748 99016 123790 99056
rect 123830 99016 123872 99056
rect 123912 99016 138664 99056
rect 138704 99016 138746 99056
rect 138786 99016 138828 99056
rect 138868 99016 138910 99056
rect 138950 99016 138992 99056
rect 139032 99016 148320 99056
rect 75648 98992 148320 99016
rect 75648 98300 148320 98324
rect 75648 98260 79424 98300
rect 79464 98260 79506 98300
rect 79546 98260 79588 98300
rect 79628 98260 79670 98300
rect 79710 98260 79752 98300
rect 79792 98260 94544 98300
rect 94584 98260 94626 98300
rect 94666 98260 94708 98300
rect 94748 98260 94790 98300
rect 94830 98260 94872 98300
rect 94912 98260 109664 98300
rect 109704 98260 109746 98300
rect 109786 98260 109828 98300
rect 109868 98260 109910 98300
rect 109950 98260 109992 98300
rect 110032 98260 124784 98300
rect 124824 98260 124866 98300
rect 124906 98260 124948 98300
rect 124988 98260 125030 98300
rect 125070 98260 125112 98300
rect 125152 98260 139904 98300
rect 139944 98260 139986 98300
rect 140026 98260 140068 98300
rect 140108 98260 140150 98300
rect 140190 98260 140232 98300
rect 140272 98260 148320 98300
rect 75648 98236 148320 98260
rect 75648 97544 148320 97568
rect 75648 97504 78184 97544
rect 78224 97504 78266 97544
rect 78306 97504 78348 97544
rect 78388 97504 78430 97544
rect 78470 97504 78512 97544
rect 78552 97504 93304 97544
rect 93344 97504 93386 97544
rect 93426 97504 93468 97544
rect 93508 97504 93550 97544
rect 93590 97504 93632 97544
rect 93672 97504 108424 97544
rect 108464 97504 108506 97544
rect 108546 97504 108588 97544
rect 108628 97504 108670 97544
rect 108710 97504 108752 97544
rect 108792 97504 123544 97544
rect 123584 97504 123626 97544
rect 123666 97504 123708 97544
rect 123748 97504 123790 97544
rect 123830 97504 123872 97544
rect 123912 97504 138664 97544
rect 138704 97504 138746 97544
rect 138786 97504 138828 97544
rect 138868 97504 138910 97544
rect 138950 97504 138992 97544
rect 139032 97504 148320 97544
rect 75648 97480 148320 97504
rect 75648 96788 148320 96812
rect 75648 96748 79424 96788
rect 79464 96748 79506 96788
rect 79546 96748 79588 96788
rect 79628 96748 79670 96788
rect 79710 96748 79752 96788
rect 79792 96748 94544 96788
rect 94584 96748 94626 96788
rect 94666 96748 94708 96788
rect 94748 96748 94790 96788
rect 94830 96748 94872 96788
rect 94912 96748 109664 96788
rect 109704 96748 109746 96788
rect 109786 96748 109828 96788
rect 109868 96748 109910 96788
rect 109950 96748 109992 96788
rect 110032 96748 124784 96788
rect 124824 96748 124866 96788
rect 124906 96748 124948 96788
rect 124988 96748 125030 96788
rect 125070 96748 125112 96788
rect 125152 96748 139904 96788
rect 139944 96748 139986 96788
rect 140026 96748 140068 96788
rect 140108 96748 140150 96788
rect 140190 96748 140232 96788
rect 140272 96748 148320 96788
rect 75648 96724 148320 96748
rect 75648 96032 148320 96056
rect 75648 95992 78184 96032
rect 78224 95992 78266 96032
rect 78306 95992 78348 96032
rect 78388 95992 78430 96032
rect 78470 95992 78512 96032
rect 78552 95992 93304 96032
rect 93344 95992 93386 96032
rect 93426 95992 93468 96032
rect 93508 95992 93550 96032
rect 93590 95992 93632 96032
rect 93672 95992 108424 96032
rect 108464 95992 108506 96032
rect 108546 95992 108588 96032
rect 108628 95992 108670 96032
rect 108710 95992 108752 96032
rect 108792 95992 123544 96032
rect 123584 95992 123626 96032
rect 123666 95992 123708 96032
rect 123748 95992 123790 96032
rect 123830 95992 123872 96032
rect 123912 95992 138664 96032
rect 138704 95992 138746 96032
rect 138786 95992 138828 96032
rect 138868 95992 138910 96032
rect 138950 95992 138992 96032
rect 139032 95992 148320 96032
rect 75648 95968 148320 95992
rect 104323 95864 104381 95865
rect 104323 95824 104332 95864
rect 104372 95824 104381 95864
rect 104323 95823 104381 95824
rect 103651 95612 103709 95613
rect 103651 95572 103660 95612
rect 103700 95572 103709 95612
rect 103651 95571 103709 95572
rect 75648 95276 148320 95300
rect 75648 95236 79424 95276
rect 79464 95236 79506 95276
rect 79546 95236 79588 95276
rect 79628 95236 79670 95276
rect 79710 95236 79752 95276
rect 79792 95236 94544 95276
rect 94584 95236 94626 95276
rect 94666 95236 94708 95276
rect 94748 95236 94790 95276
rect 94830 95236 94872 95276
rect 94912 95236 109664 95276
rect 109704 95236 109746 95276
rect 109786 95236 109828 95276
rect 109868 95236 109910 95276
rect 109950 95236 109992 95276
rect 110032 95236 124784 95276
rect 124824 95236 124866 95276
rect 124906 95236 124948 95276
rect 124988 95236 125030 95276
rect 125070 95236 125112 95276
rect 125152 95236 139904 95276
rect 139944 95236 139986 95276
rect 140026 95236 140068 95276
rect 140108 95236 140150 95276
rect 140190 95236 140232 95276
rect 140272 95236 148320 95276
rect 75648 95212 148320 95236
rect 75648 94520 148320 94544
rect 75648 94480 78184 94520
rect 78224 94480 78266 94520
rect 78306 94480 78348 94520
rect 78388 94480 78430 94520
rect 78470 94480 78512 94520
rect 78552 94480 93304 94520
rect 93344 94480 93386 94520
rect 93426 94480 93468 94520
rect 93508 94480 93550 94520
rect 93590 94480 93632 94520
rect 93672 94480 108424 94520
rect 108464 94480 108506 94520
rect 108546 94480 108588 94520
rect 108628 94480 108670 94520
rect 108710 94480 108752 94520
rect 108792 94480 123544 94520
rect 123584 94480 123626 94520
rect 123666 94480 123708 94520
rect 123748 94480 123790 94520
rect 123830 94480 123872 94520
rect 123912 94480 138664 94520
rect 138704 94480 138746 94520
rect 138786 94480 138828 94520
rect 138868 94480 138910 94520
rect 138950 94480 138992 94520
rect 139032 94480 148320 94520
rect 75648 94456 148320 94480
rect 75648 93764 148320 93788
rect 75648 93724 79424 93764
rect 79464 93724 79506 93764
rect 79546 93724 79588 93764
rect 79628 93724 79670 93764
rect 79710 93724 79752 93764
rect 79792 93724 94544 93764
rect 94584 93724 94626 93764
rect 94666 93724 94708 93764
rect 94748 93724 94790 93764
rect 94830 93724 94872 93764
rect 94912 93724 109664 93764
rect 109704 93724 109746 93764
rect 109786 93724 109828 93764
rect 109868 93724 109910 93764
rect 109950 93724 109992 93764
rect 110032 93724 124784 93764
rect 124824 93724 124866 93764
rect 124906 93724 124948 93764
rect 124988 93724 125030 93764
rect 125070 93724 125112 93764
rect 125152 93724 139904 93764
rect 139944 93724 139986 93764
rect 140026 93724 140068 93764
rect 140108 93724 140150 93764
rect 140190 93724 140232 93764
rect 140272 93724 148320 93764
rect 75648 93700 148320 93724
rect 75648 93008 148320 93032
rect 75648 92968 78184 93008
rect 78224 92968 78266 93008
rect 78306 92968 78348 93008
rect 78388 92968 78430 93008
rect 78470 92968 78512 93008
rect 78552 92968 93304 93008
rect 93344 92968 93386 93008
rect 93426 92968 93468 93008
rect 93508 92968 93550 93008
rect 93590 92968 93632 93008
rect 93672 92968 108424 93008
rect 108464 92968 108506 93008
rect 108546 92968 108588 93008
rect 108628 92968 108670 93008
rect 108710 92968 108752 93008
rect 108792 92968 123544 93008
rect 123584 92968 123626 93008
rect 123666 92968 123708 93008
rect 123748 92968 123790 93008
rect 123830 92968 123872 93008
rect 123912 92968 138664 93008
rect 138704 92968 138746 93008
rect 138786 92968 138828 93008
rect 138868 92968 138910 93008
rect 138950 92968 138992 93008
rect 139032 92968 148320 93008
rect 75648 92944 148320 92968
rect 75648 92252 148320 92276
rect 75648 92212 79424 92252
rect 79464 92212 79506 92252
rect 79546 92212 79588 92252
rect 79628 92212 79670 92252
rect 79710 92212 79752 92252
rect 79792 92212 94544 92252
rect 94584 92212 94626 92252
rect 94666 92212 94708 92252
rect 94748 92212 94790 92252
rect 94830 92212 94872 92252
rect 94912 92212 109664 92252
rect 109704 92212 109746 92252
rect 109786 92212 109828 92252
rect 109868 92212 109910 92252
rect 109950 92212 109992 92252
rect 110032 92212 124784 92252
rect 124824 92212 124866 92252
rect 124906 92212 124948 92252
rect 124988 92212 125030 92252
rect 125070 92212 125112 92252
rect 125152 92212 139904 92252
rect 139944 92212 139986 92252
rect 140026 92212 140068 92252
rect 140108 92212 140150 92252
rect 140190 92212 140232 92252
rect 140272 92212 148320 92252
rect 75648 92188 148320 92212
rect 75648 91496 148320 91520
rect 75648 91456 78184 91496
rect 78224 91456 78266 91496
rect 78306 91456 78348 91496
rect 78388 91456 78430 91496
rect 78470 91456 78512 91496
rect 78552 91456 93304 91496
rect 93344 91456 93386 91496
rect 93426 91456 93468 91496
rect 93508 91456 93550 91496
rect 93590 91456 93632 91496
rect 93672 91456 108424 91496
rect 108464 91456 108506 91496
rect 108546 91456 108588 91496
rect 108628 91456 108670 91496
rect 108710 91456 108752 91496
rect 108792 91456 123544 91496
rect 123584 91456 123626 91496
rect 123666 91456 123708 91496
rect 123748 91456 123790 91496
rect 123830 91456 123872 91496
rect 123912 91456 138664 91496
rect 138704 91456 138746 91496
rect 138786 91456 138828 91496
rect 138868 91456 138910 91496
rect 138950 91456 138992 91496
rect 139032 91456 148320 91496
rect 75648 91432 148320 91456
rect 75648 90740 148320 90764
rect 75648 90700 79424 90740
rect 79464 90700 79506 90740
rect 79546 90700 79588 90740
rect 79628 90700 79670 90740
rect 79710 90700 79752 90740
rect 79792 90700 94544 90740
rect 94584 90700 94626 90740
rect 94666 90700 94708 90740
rect 94748 90700 94790 90740
rect 94830 90700 94872 90740
rect 94912 90700 109664 90740
rect 109704 90700 109746 90740
rect 109786 90700 109828 90740
rect 109868 90700 109910 90740
rect 109950 90700 109992 90740
rect 110032 90700 124784 90740
rect 124824 90700 124866 90740
rect 124906 90700 124948 90740
rect 124988 90700 125030 90740
rect 125070 90700 125112 90740
rect 125152 90700 139904 90740
rect 139944 90700 139986 90740
rect 140026 90700 140068 90740
rect 140108 90700 140150 90740
rect 140190 90700 140232 90740
rect 140272 90700 148320 90740
rect 75648 90676 148320 90700
rect 75648 89984 148320 90008
rect 75648 89944 78184 89984
rect 78224 89944 78266 89984
rect 78306 89944 78348 89984
rect 78388 89944 78430 89984
rect 78470 89944 78512 89984
rect 78552 89944 93304 89984
rect 93344 89944 93386 89984
rect 93426 89944 93468 89984
rect 93508 89944 93550 89984
rect 93590 89944 93632 89984
rect 93672 89944 108424 89984
rect 108464 89944 108506 89984
rect 108546 89944 108588 89984
rect 108628 89944 108670 89984
rect 108710 89944 108752 89984
rect 108792 89944 123544 89984
rect 123584 89944 123626 89984
rect 123666 89944 123708 89984
rect 123748 89944 123790 89984
rect 123830 89944 123872 89984
rect 123912 89944 138664 89984
rect 138704 89944 138746 89984
rect 138786 89944 138828 89984
rect 138868 89944 138910 89984
rect 138950 89944 138992 89984
rect 139032 89944 148320 89984
rect 75648 89920 148320 89944
rect 75648 89228 148320 89252
rect 75648 89188 79424 89228
rect 79464 89188 79506 89228
rect 79546 89188 79588 89228
rect 79628 89188 79670 89228
rect 79710 89188 79752 89228
rect 79792 89188 94544 89228
rect 94584 89188 94626 89228
rect 94666 89188 94708 89228
rect 94748 89188 94790 89228
rect 94830 89188 94872 89228
rect 94912 89188 109664 89228
rect 109704 89188 109746 89228
rect 109786 89188 109828 89228
rect 109868 89188 109910 89228
rect 109950 89188 109992 89228
rect 110032 89188 124784 89228
rect 124824 89188 124866 89228
rect 124906 89188 124948 89228
rect 124988 89188 125030 89228
rect 125070 89188 125112 89228
rect 125152 89188 139904 89228
rect 139944 89188 139986 89228
rect 140026 89188 140068 89228
rect 140108 89188 140150 89228
rect 140190 89188 140232 89228
rect 140272 89188 148320 89228
rect 75648 89164 148320 89188
rect 75648 88472 148320 88496
rect 75648 88432 78184 88472
rect 78224 88432 78266 88472
rect 78306 88432 78348 88472
rect 78388 88432 78430 88472
rect 78470 88432 78512 88472
rect 78552 88432 93304 88472
rect 93344 88432 93386 88472
rect 93426 88432 93468 88472
rect 93508 88432 93550 88472
rect 93590 88432 93632 88472
rect 93672 88432 108424 88472
rect 108464 88432 108506 88472
rect 108546 88432 108588 88472
rect 108628 88432 108670 88472
rect 108710 88432 108752 88472
rect 108792 88432 123544 88472
rect 123584 88432 123626 88472
rect 123666 88432 123708 88472
rect 123748 88432 123790 88472
rect 123830 88432 123872 88472
rect 123912 88432 138664 88472
rect 138704 88432 138746 88472
rect 138786 88432 138828 88472
rect 138868 88432 138910 88472
rect 138950 88432 138992 88472
rect 139032 88432 148320 88472
rect 75648 88408 148320 88432
rect 148195 87884 148253 87885
rect 148195 87844 148204 87884
rect 148244 87844 148253 87884
rect 148195 87843 148253 87844
rect 75648 87716 148320 87740
rect 75648 87676 79424 87716
rect 79464 87676 79506 87716
rect 79546 87676 79588 87716
rect 79628 87676 79670 87716
rect 79710 87676 79752 87716
rect 79792 87676 94544 87716
rect 94584 87676 94626 87716
rect 94666 87676 94708 87716
rect 94748 87676 94790 87716
rect 94830 87676 94872 87716
rect 94912 87676 109664 87716
rect 109704 87676 109746 87716
rect 109786 87676 109828 87716
rect 109868 87676 109910 87716
rect 109950 87676 109992 87716
rect 110032 87676 124784 87716
rect 124824 87676 124866 87716
rect 124906 87676 124948 87716
rect 124988 87676 125030 87716
rect 125070 87676 125112 87716
rect 125152 87676 139904 87716
rect 139944 87676 139986 87716
rect 140026 87676 140068 87716
rect 140108 87676 140150 87716
rect 140190 87676 140232 87716
rect 140272 87676 148320 87716
rect 75648 87652 148320 87676
rect 75648 86960 148320 86984
rect 75648 86920 78184 86960
rect 78224 86920 78266 86960
rect 78306 86920 78348 86960
rect 78388 86920 78430 86960
rect 78470 86920 78512 86960
rect 78552 86920 93304 86960
rect 93344 86920 93386 86960
rect 93426 86920 93468 86960
rect 93508 86920 93550 86960
rect 93590 86920 93632 86960
rect 93672 86920 108424 86960
rect 108464 86920 108506 86960
rect 108546 86920 108588 86960
rect 108628 86920 108670 86960
rect 108710 86920 108752 86960
rect 108792 86920 123544 86960
rect 123584 86920 123626 86960
rect 123666 86920 123708 86960
rect 123748 86920 123790 86960
rect 123830 86920 123872 86960
rect 123912 86920 138664 86960
rect 138704 86920 138746 86960
rect 138786 86920 138828 86960
rect 138868 86920 138910 86960
rect 138950 86920 138992 86960
rect 139032 86920 148320 86960
rect 75648 86896 148320 86920
rect 75648 86204 148320 86228
rect 75648 86164 79424 86204
rect 79464 86164 79506 86204
rect 79546 86164 79588 86204
rect 79628 86164 79670 86204
rect 79710 86164 79752 86204
rect 79792 86164 94544 86204
rect 94584 86164 94626 86204
rect 94666 86164 94708 86204
rect 94748 86164 94790 86204
rect 94830 86164 94872 86204
rect 94912 86164 109664 86204
rect 109704 86164 109746 86204
rect 109786 86164 109828 86204
rect 109868 86164 109910 86204
rect 109950 86164 109992 86204
rect 110032 86164 124784 86204
rect 124824 86164 124866 86204
rect 124906 86164 124948 86204
rect 124988 86164 125030 86204
rect 125070 86164 125112 86204
rect 125152 86164 139904 86204
rect 139944 86164 139986 86204
rect 140026 86164 140068 86204
rect 140108 86164 140150 86204
rect 140190 86164 140232 86204
rect 140272 86164 148320 86204
rect 75648 86140 148320 86164
rect 75648 85448 148320 85472
rect 75648 85408 78184 85448
rect 78224 85408 78266 85448
rect 78306 85408 78348 85448
rect 78388 85408 78430 85448
rect 78470 85408 78512 85448
rect 78552 85408 93304 85448
rect 93344 85408 93386 85448
rect 93426 85408 93468 85448
rect 93508 85408 93550 85448
rect 93590 85408 93632 85448
rect 93672 85408 108424 85448
rect 108464 85408 108506 85448
rect 108546 85408 108588 85448
rect 108628 85408 108670 85448
rect 108710 85408 108752 85448
rect 108792 85408 123544 85448
rect 123584 85408 123626 85448
rect 123666 85408 123708 85448
rect 123748 85408 123790 85448
rect 123830 85408 123872 85448
rect 123912 85408 138664 85448
rect 138704 85408 138746 85448
rect 138786 85408 138828 85448
rect 138868 85408 138910 85448
rect 138950 85408 138992 85448
rect 139032 85408 148320 85448
rect 75648 85384 148320 85408
rect 75648 84692 148320 84716
rect 75648 84652 79424 84692
rect 79464 84652 79506 84692
rect 79546 84652 79588 84692
rect 79628 84652 79670 84692
rect 79710 84652 79752 84692
rect 79792 84652 94544 84692
rect 94584 84652 94626 84692
rect 94666 84652 94708 84692
rect 94748 84652 94790 84692
rect 94830 84652 94872 84692
rect 94912 84652 109664 84692
rect 109704 84652 109746 84692
rect 109786 84652 109828 84692
rect 109868 84652 109910 84692
rect 109950 84652 109992 84692
rect 110032 84652 124784 84692
rect 124824 84652 124866 84692
rect 124906 84652 124948 84692
rect 124988 84652 125030 84692
rect 125070 84652 125112 84692
rect 125152 84652 139904 84692
rect 139944 84652 139986 84692
rect 140026 84652 140068 84692
rect 140108 84652 140150 84692
rect 140190 84652 140232 84692
rect 140272 84652 148320 84692
rect 75648 84628 148320 84652
rect 75648 83936 148320 83960
rect 75648 83896 78184 83936
rect 78224 83896 78266 83936
rect 78306 83896 78348 83936
rect 78388 83896 78430 83936
rect 78470 83896 78512 83936
rect 78552 83896 93304 83936
rect 93344 83896 93386 83936
rect 93426 83896 93468 83936
rect 93508 83896 93550 83936
rect 93590 83896 93632 83936
rect 93672 83896 108424 83936
rect 108464 83896 108506 83936
rect 108546 83896 108588 83936
rect 108628 83896 108670 83936
rect 108710 83896 108752 83936
rect 108792 83896 123544 83936
rect 123584 83896 123626 83936
rect 123666 83896 123708 83936
rect 123748 83896 123790 83936
rect 123830 83896 123872 83936
rect 123912 83896 138664 83936
rect 138704 83896 138746 83936
rect 138786 83896 138828 83936
rect 138868 83896 138910 83936
rect 138950 83896 138992 83936
rect 139032 83896 148320 83936
rect 75648 83872 148320 83896
rect 75648 83180 148320 83204
rect 75648 83140 79424 83180
rect 79464 83140 79506 83180
rect 79546 83140 79588 83180
rect 79628 83140 79670 83180
rect 79710 83140 79752 83180
rect 79792 83140 94544 83180
rect 94584 83140 94626 83180
rect 94666 83140 94708 83180
rect 94748 83140 94790 83180
rect 94830 83140 94872 83180
rect 94912 83140 109664 83180
rect 109704 83140 109746 83180
rect 109786 83140 109828 83180
rect 109868 83140 109910 83180
rect 109950 83140 109992 83180
rect 110032 83140 124784 83180
rect 124824 83140 124866 83180
rect 124906 83140 124948 83180
rect 124988 83140 125030 83180
rect 125070 83140 125112 83180
rect 125152 83140 139904 83180
rect 139944 83140 139986 83180
rect 140026 83140 140068 83180
rect 140108 83140 140150 83180
rect 140190 83140 140232 83180
rect 140272 83140 148320 83180
rect 75648 83116 148320 83140
rect 75648 82424 148320 82448
rect 75648 82384 78184 82424
rect 78224 82384 78266 82424
rect 78306 82384 78348 82424
rect 78388 82384 78430 82424
rect 78470 82384 78512 82424
rect 78552 82384 93304 82424
rect 93344 82384 93386 82424
rect 93426 82384 93468 82424
rect 93508 82384 93550 82424
rect 93590 82384 93632 82424
rect 93672 82384 108424 82424
rect 108464 82384 108506 82424
rect 108546 82384 108588 82424
rect 108628 82384 108670 82424
rect 108710 82384 108752 82424
rect 108792 82384 123544 82424
rect 123584 82384 123626 82424
rect 123666 82384 123708 82424
rect 123748 82384 123790 82424
rect 123830 82384 123872 82424
rect 123912 82384 138664 82424
rect 138704 82384 138746 82424
rect 138786 82384 138828 82424
rect 138868 82384 138910 82424
rect 138950 82384 138992 82424
rect 139032 82384 148320 82424
rect 75648 82360 148320 82384
rect 75648 81668 148320 81692
rect 75648 81628 79424 81668
rect 79464 81628 79506 81668
rect 79546 81628 79588 81668
rect 79628 81628 79670 81668
rect 79710 81628 79752 81668
rect 79792 81628 94544 81668
rect 94584 81628 94626 81668
rect 94666 81628 94708 81668
rect 94748 81628 94790 81668
rect 94830 81628 94872 81668
rect 94912 81628 109664 81668
rect 109704 81628 109746 81668
rect 109786 81628 109828 81668
rect 109868 81628 109910 81668
rect 109950 81628 109992 81668
rect 110032 81628 124784 81668
rect 124824 81628 124866 81668
rect 124906 81628 124948 81668
rect 124988 81628 125030 81668
rect 125070 81628 125112 81668
rect 125152 81628 139904 81668
rect 139944 81628 139986 81668
rect 140026 81628 140068 81668
rect 140108 81628 140150 81668
rect 140190 81628 140232 81668
rect 140272 81628 148320 81668
rect 75648 81604 148320 81628
rect 75648 80912 148320 80936
rect 75648 80872 78184 80912
rect 78224 80872 78266 80912
rect 78306 80872 78348 80912
rect 78388 80872 78430 80912
rect 78470 80872 78512 80912
rect 78552 80872 93304 80912
rect 93344 80872 93386 80912
rect 93426 80872 93468 80912
rect 93508 80872 93550 80912
rect 93590 80872 93632 80912
rect 93672 80872 108424 80912
rect 108464 80872 108506 80912
rect 108546 80872 108588 80912
rect 108628 80872 108670 80912
rect 108710 80872 108752 80912
rect 108792 80872 123544 80912
rect 123584 80872 123626 80912
rect 123666 80872 123708 80912
rect 123748 80872 123790 80912
rect 123830 80872 123872 80912
rect 123912 80872 138664 80912
rect 138704 80872 138746 80912
rect 138786 80872 138828 80912
rect 138868 80872 138910 80912
rect 138950 80872 138992 80912
rect 139032 80872 148320 80912
rect 75648 80848 148320 80872
rect 75648 80156 148320 80180
rect 75648 80116 79424 80156
rect 79464 80116 79506 80156
rect 79546 80116 79588 80156
rect 79628 80116 79670 80156
rect 79710 80116 79752 80156
rect 79792 80116 94544 80156
rect 94584 80116 94626 80156
rect 94666 80116 94708 80156
rect 94748 80116 94790 80156
rect 94830 80116 94872 80156
rect 94912 80116 109664 80156
rect 109704 80116 109746 80156
rect 109786 80116 109828 80156
rect 109868 80116 109910 80156
rect 109950 80116 109992 80156
rect 110032 80116 124784 80156
rect 124824 80116 124866 80156
rect 124906 80116 124948 80156
rect 124988 80116 125030 80156
rect 125070 80116 125112 80156
rect 125152 80116 139904 80156
rect 139944 80116 139986 80156
rect 140026 80116 140068 80156
rect 140108 80116 140150 80156
rect 140190 80116 140232 80156
rect 140272 80116 148320 80156
rect 75648 80092 148320 80116
rect 75648 79400 148320 79424
rect 75648 79360 78184 79400
rect 78224 79360 78266 79400
rect 78306 79360 78348 79400
rect 78388 79360 78430 79400
rect 78470 79360 78512 79400
rect 78552 79360 93304 79400
rect 93344 79360 93386 79400
rect 93426 79360 93468 79400
rect 93508 79360 93550 79400
rect 93590 79360 93632 79400
rect 93672 79360 108424 79400
rect 108464 79360 108506 79400
rect 108546 79360 108588 79400
rect 108628 79360 108670 79400
rect 108710 79360 108752 79400
rect 108792 79360 123544 79400
rect 123584 79360 123626 79400
rect 123666 79360 123708 79400
rect 123748 79360 123790 79400
rect 123830 79360 123872 79400
rect 123912 79360 138664 79400
rect 138704 79360 138746 79400
rect 138786 79360 138828 79400
rect 138868 79360 138910 79400
rect 138950 79360 138992 79400
rect 139032 79360 148320 79400
rect 75648 79336 148320 79360
rect 75648 78644 148320 78668
rect 75648 78604 79424 78644
rect 79464 78604 79506 78644
rect 79546 78604 79588 78644
rect 79628 78604 79670 78644
rect 79710 78604 79752 78644
rect 79792 78604 94544 78644
rect 94584 78604 94626 78644
rect 94666 78604 94708 78644
rect 94748 78604 94790 78644
rect 94830 78604 94872 78644
rect 94912 78604 109664 78644
rect 109704 78604 109746 78644
rect 109786 78604 109828 78644
rect 109868 78604 109910 78644
rect 109950 78604 109992 78644
rect 110032 78604 124784 78644
rect 124824 78604 124866 78644
rect 124906 78604 124948 78644
rect 124988 78604 125030 78644
rect 125070 78604 125112 78644
rect 125152 78604 139904 78644
rect 139944 78604 139986 78644
rect 140026 78604 140068 78644
rect 140108 78604 140150 78644
rect 140190 78604 140232 78644
rect 140272 78604 148320 78644
rect 75648 78580 148320 78604
rect 75648 77888 148320 77912
rect 75648 77848 78184 77888
rect 78224 77848 78266 77888
rect 78306 77848 78348 77888
rect 78388 77848 78430 77888
rect 78470 77848 78512 77888
rect 78552 77848 93304 77888
rect 93344 77848 93386 77888
rect 93426 77848 93468 77888
rect 93508 77848 93550 77888
rect 93590 77848 93632 77888
rect 93672 77848 108424 77888
rect 108464 77848 108506 77888
rect 108546 77848 108588 77888
rect 108628 77848 108670 77888
rect 108710 77848 108752 77888
rect 108792 77848 123544 77888
rect 123584 77848 123626 77888
rect 123666 77848 123708 77888
rect 123748 77848 123790 77888
rect 123830 77848 123872 77888
rect 123912 77848 138664 77888
rect 138704 77848 138746 77888
rect 138786 77848 138828 77888
rect 138868 77848 138910 77888
rect 138950 77848 138992 77888
rect 139032 77848 148320 77888
rect 75648 77824 148320 77848
rect 75648 77132 148320 77156
rect 75648 77092 79424 77132
rect 79464 77092 79506 77132
rect 79546 77092 79588 77132
rect 79628 77092 79670 77132
rect 79710 77092 79752 77132
rect 79792 77092 94544 77132
rect 94584 77092 94626 77132
rect 94666 77092 94708 77132
rect 94748 77092 94790 77132
rect 94830 77092 94872 77132
rect 94912 77092 109664 77132
rect 109704 77092 109746 77132
rect 109786 77092 109828 77132
rect 109868 77092 109910 77132
rect 109950 77092 109992 77132
rect 110032 77092 124784 77132
rect 124824 77092 124866 77132
rect 124906 77092 124948 77132
rect 124988 77092 125030 77132
rect 125070 77092 125112 77132
rect 125152 77092 139904 77132
rect 139944 77092 139986 77132
rect 140026 77092 140068 77132
rect 140108 77092 140150 77132
rect 140190 77092 140232 77132
rect 140272 77092 148320 77132
rect 75648 77068 148320 77092
rect 75648 76376 148320 76400
rect 75648 76336 78184 76376
rect 78224 76336 78266 76376
rect 78306 76336 78348 76376
rect 78388 76336 78430 76376
rect 78470 76336 78512 76376
rect 78552 76336 93304 76376
rect 93344 76336 93386 76376
rect 93426 76336 93468 76376
rect 93508 76336 93550 76376
rect 93590 76336 93632 76376
rect 93672 76336 108424 76376
rect 108464 76336 108506 76376
rect 108546 76336 108588 76376
rect 108628 76336 108670 76376
rect 108710 76336 108752 76376
rect 108792 76336 123544 76376
rect 123584 76336 123626 76376
rect 123666 76336 123708 76376
rect 123748 76336 123790 76376
rect 123830 76336 123872 76376
rect 123912 76336 138664 76376
rect 138704 76336 138746 76376
rect 138786 76336 138828 76376
rect 138868 76336 138910 76376
rect 138950 76336 138992 76376
rect 139032 76336 148320 76376
rect 75648 76312 148320 76336
rect 148195 75788 148253 75789
rect 148195 75748 148204 75788
rect 148244 75748 148253 75788
rect 148195 75747 148253 75748
rect 75648 75620 148320 75644
rect 75648 75580 79424 75620
rect 79464 75580 79506 75620
rect 79546 75580 79588 75620
rect 79628 75580 79670 75620
rect 79710 75580 79752 75620
rect 79792 75580 94544 75620
rect 94584 75580 94626 75620
rect 94666 75580 94708 75620
rect 94748 75580 94790 75620
rect 94830 75580 94872 75620
rect 94912 75580 109664 75620
rect 109704 75580 109746 75620
rect 109786 75580 109828 75620
rect 109868 75580 109910 75620
rect 109950 75580 109992 75620
rect 110032 75580 124784 75620
rect 124824 75580 124866 75620
rect 124906 75580 124948 75620
rect 124988 75580 125030 75620
rect 125070 75580 125112 75620
rect 125152 75580 139904 75620
rect 139944 75580 139986 75620
rect 140026 75580 140068 75620
rect 140108 75580 140150 75620
rect 140190 75580 140232 75620
rect 140272 75580 148320 75620
rect 75648 75556 148320 75580
<< via1 >>
rect 79424 148156 79464 148196
rect 79506 148156 79546 148196
rect 79588 148156 79628 148196
rect 79670 148156 79710 148196
rect 79752 148156 79792 148196
rect 94544 148156 94584 148196
rect 94626 148156 94666 148196
rect 94708 148156 94748 148196
rect 94790 148156 94830 148196
rect 94872 148156 94912 148196
rect 109664 148156 109704 148196
rect 109746 148156 109786 148196
rect 109828 148156 109868 148196
rect 109910 148156 109950 148196
rect 109992 148156 110032 148196
rect 124784 148156 124824 148196
rect 124866 148156 124906 148196
rect 124948 148156 124988 148196
rect 125030 148156 125070 148196
rect 125112 148156 125152 148196
rect 139904 148156 139944 148196
rect 139986 148156 140026 148196
rect 140068 148156 140108 148196
rect 140150 148156 140190 148196
rect 140232 148156 140272 148196
rect 78184 147400 78224 147440
rect 78266 147400 78306 147440
rect 78348 147400 78388 147440
rect 78430 147400 78470 147440
rect 78512 147400 78552 147440
rect 93304 147400 93344 147440
rect 93386 147400 93426 147440
rect 93468 147400 93508 147440
rect 93550 147400 93590 147440
rect 93632 147400 93672 147440
rect 108424 147400 108464 147440
rect 108506 147400 108546 147440
rect 108588 147400 108628 147440
rect 108670 147400 108710 147440
rect 108752 147400 108792 147440
rect 123544 147400 123584 147440
rect 123626 147400 123666 147440
rect 123708 147400 123748 147440
rect 123790 147400 123830 147440
rect 123872 147400 123912 147440
rect 138664 147400 138704 147440
rect 138746 147400 138786 147440
rect 138828 147400 138868 147440
rect 138910 147400 138950 147440
rect 138992 147400 139032 147440
rect 79424 146644 79464 146684
rect 79506 146644 79546 146684
rect 79588 146644 79628 146684
rect 79670 146644 79710 146684
rect 79752 146644 79792 146684
rect 94544 146644 94584 146684
rect 94626 146644 94666 146684
rect 94708 146644 94748 146684
rect 94790 146644 94830 146684
rect 94872 146644 94912 146684
rect 109664 146644 109704 146684
rect 109746 146644 109786 146684
rect 109828 146644 109868 146684
rect 109910 146644 109950 146684
rect 109992 146644 110032 146684
rect 124784 146644 124824 146684
rect 124866 146644 124906 146684
rect 124948 146644 124988 146684
rect 125030 146644 125070 146684
rect 125112 146644 125152 146684
rect 139904 146644 139944 146684
rect 139986 146644 140026 146684
rect 140068 146644 140108 146684
rect 140150 146644 140190 146684
rect 140232 146644 140272 146684
rect 78184 145888 78224 145928
rect 78266 145888 78306 145928
rect 78348 145888 78388 145928
rect 78430 145888 78470 145928
rect 78512 145888 78552 145928
rect 93304 145888 93344 145928
rect 93386 145888 93426 145928
rect 93468 145888 93508 145928
rect 93550 145888 93590 145928
rect 93632 145888 93672 145928
rect 108424 145888 108464 145928
rect 108506 145888 108546 145928
rect 108588 145888 108628 145928
rect 108670 145888 108710 145928
rect 108752 145888 108792 145928
rect 123544 145888 123584 145928
rect 123626 145888 123666 145928
rect 123708 145888 123748 145928
rect 123790 145888 123830 145928
rect 123872 145888 123912 145928
rect 138664 145888 138704 145928
rect 138746 145888 138786 145928
rect 138828 145888 138868 145928
rect 138910 145888 138950 145928
rect 138992 145888 139032 145928
rect 79424 145132 79464 145172
rect 79506 145132 79546 145172
rect 79588 145132 79628 145172
rect 79670 145132 79710 145172
rect 79752 145132 79792 145172
rect 94544 145132 94584 145172
rect 94626 145132 94666 145172
rect 94708 145132 94748 145172
rect 94790 145132 94830 145172
rect 94872 145132 94912 145172
rect 109664 145132 109704 145172
rect 109746 145132 109786 145172
rect 109828 145132 109868 145172
rect 109910 145132 109950 145172
rect 109992 145132 110032 145172
rect 124784 145132 124824 145172
rect 124866 145132 124906 145172
rect 124948 145132 124988 145172
rect 125030 145132 125070 145172
rect 125112 145132 125152 145172
rect 139904 145132 139944 145172
rect 139986 145132 140026 145172
rect 140068 145132 140108 145172
rect 140150 145132 140190 145172
rect 140232 145132 140272 145172
rect 78184 144376 78224 144416
rect 78266 144376 78306 144416
rect 78348 144376 78388 144416
rect 78430 144376 78470 144416
rect 78512 144376 78552 144416
rect 93304 144376 93344 144416
rect 93386 144376 93426 144416
rect 93468 144376 93508 144416
rect 93550 144376 93590 144416
rect 93632 144376 93672 144416
rect 108424 144376 108464 144416
rect 108506 144376 108546 144416
rect 108588 144376 108628 144416
rect 108670 144376 108710 144416
rect 108752 144376 108792 144416
rect 123544 144376 123584 144416
rect 123626 144376 123666 144416
rect 123708 144376 123748 144416
rect 123790 144376 123830 144416
rect 123872 144376 123912 144416
rect 138664 144376 138704 144416
rect 138746 144376 138786 144416
rect 138828 144376 138868 144416
rect 138910 144376 138950 144416
rect 138992 144376 139032 144416
rect 79424 143620 79464 143660
rect 79506 143620 79546 143660
rect 79588 143620 79628 143660
rect 79670 143620 79710 143660
rect 79752 143620 79792 143660
rect 94544 143620 94584 143660
rect 94626 143620 94666 143660
rect 94708 143620 94748 143660
rect 94790 143620 94830 143660
rect 94872 143620 94912 143660
rect 109664 143620 109704 143660
rect 109746 143620 109786 143660
rect 109828 143620 109868 143660
rect 109910 143620 109950 143660
rect 109992 143620 110032 143660
rect 124784 143620 124824 143660
rect 124866 143620 124906 143660
rect 124948 143620 124988 143660
rect 125030 143620 125070 143660
rect 125112 143620 125152 143660
rect 139904 143620 139944 143660
rect 139986 143620 140026 143660
rect 140068 143620 140108 143660
rect 140150 143620 140190 143660
rect 140232 143620 140272 143660
rect 78184 142864 78224 142904
rect 78266 142864 78306 142904
rect 78348 142864 78388 142904
rect 78430 142864 78470 142904
rect 78512 142864 78552 142904
rect 93304 142864 93344 142904
rect 93386 142864 93426 142904
rect 93468 142864 93508 142904
rect 93550 142864 93590 142904
rect 93632 142864 93672 142904
rect 108424 142864 108464 142904
rect 108506 142864 108546 142904
rect 108588 142864 108628 142904
rect 108670 142864 108710 142904
rect 108752 142864 108792 142904
rect 123544 142864 123584 142904
rect 123626 142864 123666 142904
rect 123708 142864 123748 142904
rect 123790 142864 123830 142904
rect 123872 142864 123912 142904
rect 138664 142864 138704 142904
rect 138746 142864 138786 142904
rect 138828 142864 138868 142904
rect 138910 142864 138950 142904
rect 138992 142864 139032 142904
rect 79424 142108 79464 142148
rect 79506 142108 79546 142148
rect 79588 142108 79628 142148
rect 79670 142108 79710 142148
rect 79752 142108 79792 142148
rect 94544 142108 94584 142148
rect 94626 142108 94666 142148
rect 94708 142108 94748 142148
rect 94790 142108 94830 142148
rect 94872 142108 94912 142148
rect 109664 142108 109704 142148
rect 109746 142108 109786 142148
rect 109828 142108 109868 142148
rect 109910 142108 109950 142148
rect 109992 142108 110032 142148
rect 124784 142108 124824 142148
rect 124866 142108 124906 142148
rect 124948 142108 124988 142148
rect 125030 142108 125070 142148
rect 125112 142108 125152 142148
rect 139904 142108 139944 142148
rect 139986 142108 140026 142148
rect 140068 142108 140108 142148
rect 140150 142108 140190 142148
rect 140232 142108 140272 142148
rect 78184 141352 78224 141392
rect 78266 141352 78306 141392
rect 78348 141352 78388 141392
rect 78430 141352 78470 141392
rect 78512 141352 78552 141392
rect 93304 141352 93344 141392
rect 93386 141352 93426 141392
rect 93468 141352 93508 141392
rect 93550 141352 93590 141392
rect 93632 141352 93672 141392
rect 108424 141352 108464 141392
rect 108506 141352 108546 141392
rect 108588 141352 108628 141392
rect 108670 141352 108710 141392
rect 108752 141352 108792 141392
rect 123544 141352 123584 141392
rect 123626 141352 123666 141392
rect 123708 141352 123748 141392
rect 123790 141352 123830 141392
rect 123872 141352 123912 141392
rect 138664 141352 138704 141392
rect 138746 141352 138786 141392
rect 138828 141352 138868 141392
rect 138910 141352 138950 141392
rect 138992 141352 139032 141392
rect 79424 140596 79464 140636
rect 79506 140596 79546 140636
rect 79588 140596 79628 140636
rect 79670 140596 79710 140636
rect 79752 140596 79792 140636
rect 94544 140596 94584 140636
rect 94626 140596 94666 140636
rect 94708 140596 94748 140636
rect 94790 140596 94830 140636
rect 94872 140596 94912 140636
rect 109664 140596 109704 140636
rect 109746 140596 109786 140636
rect 109828 140596 109868 140636
rect 109910 140596 109950 140636
rect 109992 140596 110032 140636
rect 124784 140596 124824 140636
rect 124866 140596 124906 140636
rect 124948 140596 124988 140636
rect 125030 140596 125070 140636
rect 125112 140596 125152 140636
rect 139904 140596 139944 140636
rect 139986 140596 140026 140636
rect 140068 140596 140108 140636
rect 140150 140596 140190 140636
rect 140232 140596 140272 140636
rect 78184 139840 78224 139880
rect 78266 139840 78306 139880
rect 78348 139840 78388 139880
rect 78430 139840 78470 139880
rect 78512 139840 78552 139880
rect 93304 139840 93344 139880
rect 93386 139840 93426 139880
rect 93468 139840 93508 139880
rect 93550 139840 93590 139880
rect 93632 139840 93672 139880
rect 108424 139840 108464 139880
rect 108506 139840 108546 139880
rect 108588 139840 108628 139880
rect 108670 139840 108710 139880
rect 108752 139840 108792 139880
rect 123544 139840 123584 139880
rect 123626 139840 123666 139880
rect 123708 139840 123748 139880
rect 123790 139840 123830 139880
rect 123872 139840 123912 139880
rect 138664 139840 138704 139880
rect 138746 139840 138786 139880
rect 138828 139840 138868 139880
rect 138910 139840 138950 139880
rect 138992 139840 139032 139880
rect 79424 139084 79464 139124
rect 79506 139084 79546 139124
rect 79588 139084 79628 139124
rect 79670 139084 79710 139124
rect 79752 139084 79792 139124
rect 94544 139084 94584 139124
rect 94626 139084 94666 139124
rect 94708 139084 94748 139124
rect 94790 139084 94830 139124
rect 94872 139084 94912 139124
rect 109664 139084 109704 139124
rect 109746 139084 109786 139124
rect 109828 139084 109868 139124
rect 109910 139084 109950 139124
rect 109992 139084 110032 139124
rect 124784 139084 124824 139124
rect 124866 139084 124906 139124
rect 124948 139084 124988 139124
rect 125030 139084 125070 139124
rect 125112 139084 125152 139124
rect 139904 139084 139944 139124
rect 139986 139084 140026 139124
rect 140068 139084 140108 139124
rect 140150 139084 140190 139124
rect 140232 139084 140272 139124
rect 78184 138328 78224 138368
rect 78266 138328 78306 138368
rect 78348 138328 78388 138368
rect 78430 138328 78470 138368
rect 78512 138328 78552 138368
rect 93304 138328 93344 138368
rect 93386 138328 93426 138368
rect 93468 138328 93508 138368
rect 93550 138328 93590 138368
rect 93632 138328 93672 138368
rect 108424 138328 108464 138368
rect 108506 138328 108546 138368
rect 108588 138328 108628 138368
rect 108670 138328 108710 138368
rect 108752 138328 108792 138368
rect 123544 138328 123584 138368
rect 123626 138328 123666 138368
rect 123708 138328 123748 138368
rect 123790 138328 123830 138368
rect 123872 138328 123912 138368
rect 138664 138328 138704 138368
rect 138746 138328 138786 138368
rect 138828 138328 138868 138368
rect 138910 138328 138950 138368
rect 138992 138328 139032 138368
rect 79424 137572 79464 137612
rect 79506 137572 79546 137612
rect 79588 137572 79628 137612
rect 79670 137572 79710 137612
rect 79752 137572 79792 137612
rect 94544 137572 94584 137612
rect 94626 137572 94666 137612
rect 94708 137572 94748 137612
rect 94790 137572 94830 137612
rect 94872 137572 94912 137612
rect 109664 137572 109704 137612
rect 109746 137572 109786 137612
rect 109828 137572 109868 137612
rect 109910 137572 109950 137612
rect 109992 137572 110032 137612
rect 124784 137572 124824 137612
rect 124866 137572 124906 137612
rect 124948 137572 124988 137612
rect 125030 137572 125070 137612
rect 125112 137572 125152 137612
rect 139904 137572 139944 137612
rect 139986 137572 140026 137612
rect 140068 137572 140108 137612
rect 140150 137572 140190 137612
rect 140232 137572 140272 137612
rect 78184 136816 78224 136856
rect 78266 136816 78306 136856
rect 78348 136816 78388 136856
rect 78430 136816 78470 136856
rect 78512 136816 78552 136856
rect 93304 136816 93344 136856
rect 93386 136816 93426 136856
rect 93468 136816 93508 136856
rect 93550 136816 93590 136856
rect 93632 136816 93672 136856
rect 108424 136816 108464 136856
rect 108506 136816 108546 136856
rect 108588 136816 108628 136856
rect 108670 136816 108710 136856
rect 108752 136816 108792 136856
rect 123544 136816 123584 136856
rect 123626 136816 123666 136856
rect 123708 136816 123748 136856
rect 123790 136816 123830 136856
rect 123872 136816 123912 136856
rect 138664 136816 138704 136856
rect 138746 136816 138786 136856
rect 138828 136816 138868 136856
rect 138910 136816 138950 136856
rect 138992 136816 139032 136856
rect 79424 136060 79464 136100
rect 79506 136060 79546 136100
rect 79588 136060 79628 136100
rect 79670 136060 79710 136100
rect 79752 136060 79792 136100
rect 94544 136060 94584 136100
rect 94626 136060 94666 136100
rect 94708 136060 94748 136100
rect 94790 136060 94830 136100
rect 94872 136060 94912 136100
rect 109664 136060 109704 136100
rect 109746 136060 109786 136100
rect 109828 136060 109868 136100
rect 109910 136060 109950 136100
rect 109992 136060 110032 136100
rect 124784 136060 124824 136100
rect 124866 136060 124906 136100
rect 124948 136060 124988 136100
rect 125030 136060 125070 136100
rect 125112 136060 125152 136100
rect 139904 136060 139944 136100
rect 139986 136060 140026 136100
rect 140068 136060 140108 136100
rect 140150 136060 140190 136100
rect 140232 136060 140272 136100
rect 78184 135304 78224 135344
rect 78266 135304 78306 135344
rect 78348 135304 78388 135344
rect 78430 135304 78470 135344
rect 78512 135304 78552 135344
rect 93304 135304 93344 135344
rect 93386 135304 93426 135344
rect 93468 135304 93508 135344
rect 93550 135304 93590 135344
rect 93632 135304 93672 135344
rect 108424 135304 108464 135344
rect 108506 135304 108546 135344
rect 108588 135304 108628 135344
rect 108670 135304 108710 135344
rect 108752 135304 108792 135344
rect 123544 135304 123584 135344
rect 123626 135304 123666 135344
rect 123708 135304 123748 135344
rect 123790 135304 123830 135344
rect 123872 135304 123912 135344
rect 138664 135304 138704 135344
rect 138746 135304 138786 135344
rect 138828 135304 138868 135344
rect 138910 135304 138950 135344
rect 138992 135304 139032 135344
rect 79424 134548 79464 134588
rect 79506 134548 79546 134588
rect 79588 134548 79628 134588
rect 79670 134548 79710 134588
rect 79752 134548 79792 134588
rect 94544 134548 94584 134588
rect 94626 134548 94666 134588
rect 94708 134548 94748 134588
rect 94790 134548 94830 134588
rect 94872 134548 94912 134588
rect 109664 134548 109704 134588
rect 109746 134548 109786 134588
rect 109828 134548 109868 134588
rect 109910 134548 109950 134588
rect 109992 134548 110032 134588
rect 124784 134548 124824 134588
rect 124866 134548 124906 134588
rect 124948 134548 124988 134588
rect 125030 134548 125070 134588
rect 125112 134548 125152 134588
rect 139904 134548 139944 134588
rect 139986 134548 140026 134588
rect 140068 134548 140108 134588
rect 140150 134548 140190 134588
rect 140232 134548 140272 134588
rect 115948 134380 115988 134420
rect 97420 134212 97460 134252
rect 97804 134212 97844 134252
rect 98668 134212 98708 134252
rect 113548 134212 113588 134252
rect 113932 134212 113972 134252
rect 114796 134212 114836 134252
rect 99820 134044 99860 134084
rect 119884 134044 119924 134084
rect 115948 133960 115988 134000
rect 78184 133792 78224 133832
rect 78266 133792 78306 133832
rect 78348 133792 78388 133832
rect 78430 133792 78470 133832
rect 78512 133792 78552 133832
rect 93304 133792 93344 133832
rect 93386 133792 93426 133832
rect 93468 133792 93508 133832
rect 93550 133792 93590 133832
rect 93632 133792 93672 133832
rect 108424 133792 108464 133832
rect 108506 133792 108546 133832
rect 108588 133792 108628 133832
rect 108670 133792 108710 133832
rect 108752 133792 108792 133832
rect 123544 133792 123584 133832
rect 123626 133792 123666 133832
rect 123708 133792 123748 133832
rect 123790 133792 123830 133832
rect 123872 133792 123912 133832
rect 138664 133792 138704 133832
rect 138746 133792 138786 133832
rect 138828 133792 138868 133832
rect 138910 133792 138950 133832
rect 138992 133792 139032 133832
rect 98188 133624 98228 133664
rect 121804 133624 121844 133664
rect 97804 133540 97844 133580
rect 114028 133540 114068 133580
rect 98860 133372 98900 133412
rect 115084 133372 115124 133412
rect 119788 133372 119828 133412
rect 120652 133372 120692 133412
rect 119404 133288 119444 133328
rect 114412 133204 114452 133244
rect 121804 133204 121844 133244
rect 79424 133036 79464 133076
rect 79506 133036 79546 133076
rect 79588 133036 79628 133076
rect 79670 133036 79710 133076
rect 79752 133036 79792 133076
rect 94544 133036 94584 133076
rect 94626 133036 94666 133076
rect 94708 133036 94748 133076
rect 94790 133036 94830 133076
rect 94872 133036 94912 133076
rect 109664 133036 109704 133076
rect 109746 133036 109786 133076
rect 109828 133036 109868 133076
rect 109910 133036 109950 133076
rect 109992 133036 110032 133076
rect 124784 133036 124824 133076
rect 124866 133036 124906 133076
rect 124948 133036 124988 133076
rect 125030 133036 125070 133076
rect 125112 133036 125152 133076
rect 139904 133036 139944 133076
rect 139986 133036 140026 133076
rect 140068 133036 140108 133076
rect 140150 133036 140190 133076
rect 140232 133036 140272 133076
rect 98668 132868 98708 132908
rect 119404 132868 119444 132908
rect 78604 132700 78644 132740
rect 98572 132700 98612 132740
rect 98764 132700 98804 132740
rect 98860 132700 98900 132740
rect 102988 132700 103028 132740
rect 103660 132700 103700 132740
rect 103852 132700 103892 132740
rect 104236 132700 104276 132740
rect 105100 132700 105140 132740
rect 120076 132700 120116 132740
rect 120940 132700 120980 132740
rect 106252 132616 106292 132656
rect 79276 132532 79316 132572
rect 109900 132532 109940 132572
rect 120268 132532 120308 132572
rect 78184 132280 78224 132320
rect 78266 132280 78306 132320
rect 78348 132280 78388 132320
rect 78430 132280 78470 132320
rect 78512 132280 78552 132320
rect 93304 132280 93344 132320
rect 93386 132280 93426 132320
rect 93468 132280 93508 132320
rect 93550 132280 93590 132320
rect 93632 132280 93672 132320
rect 108424 132280 108464 132320
rect 108506 132280 108546 132320
rect 108588 132280 108628 132320
rect 108670 132280 108710 132320
rect 108752 132280 108792 132320
rect 123544 132280 123584 132320
rect 123626 132280 123666 132320
rect 123708 132280 123748 132320
rect 123790 132280 123830 132320
rect 123872 132280 123912 132320
rect 138664 132280 138704 132320
rect 138746 132280 138786 132320
rect 138828 132280 138868 132320
rect 138910 132280 138950 132320
rect 138992 132280 139032 132320
rect 99052 132028 99092 132068
rect 104332 132028 104372 132068
rect 98380 131860 98420 131900
rect 99244 131860 99284 131900
rect 99340 131860 99380 131900
rect 99436 131860 99476 131900
rect 99532 131860 99572 131900
rect 100012 131860 100052 131900
rect 100204 131860 100244 131900
rect 101068 131860 101108 131900
rect 101164 131860 101204 131900
rect 101356 131860 101396 131900
rect 101644 131860 101684 131900
rect 109804 131860 109844 131900
rect 110668 131860 110708 131900
rect 112204 131860 112244 131900
rect 112300 131860 112340 131900
rect 112780 131860 112820 131900
rect 118540 131860 118580 131900
rect 100108 131776 100148 131816
rect 109420 131776 109460 131816
rect 112404 131776 112444 131816
rect 101260 131692 101300 131732
rect 101548 131692 101588 131732
rect 111820 131692 111860 131732
rect 112492 131692 112532 131732
rect 112588 131692 112628 131732
rect 113452 131692 113492 131732
rect 118444 131692 118484 131732
rect 79424 131524 79464 131564
rect 79506 131524 79546 131564
rect 79588 131524 79628 131564
rect 79670 131524 79710 131564
rect 79752 131524 79792 131564
rect 94544 131524 94584 131564
rect 94626 131524 94666 131564
rect 94708 131524 94748 131564
rect 94790 131524 94830 131564
rect 94872 131524 94912 131564
rect 109664 131524 109704 131564
rect 109746 131524 109786 131564
rect 109828 131524 109868 131564
rect 109910 131524 109950 131564
rect 109992 131524 110032 131564
rect 124784 131524 124824 131564
rect 124866 131524 124906 131564
rect 124948 131524 124988 131564
rect 125030 131524 125070 131564
rect 125112 131524 125152 131564
rect 139904 131524 139944 131564
rect 139986 131524 140026 131564
rect 140068 131524 140108 131564
rect 140150 131524 140190 131564
rect 140232 131524 140272 131564
rect 102220 131356 102260 131396
rect 108844 131356 108884 131396
rect 109804 131356 109844 131396
rect 110764 131356 110804 131396
rect 112300 131356 112340 131396
rect 113068 131356 113108 131396
rect 115180 131356 115220 131396
rect 119308 131356 119348 131396
rect 113356 131272 113396 131312
rect 115084 131272 115124 131312
rect 99916 131188 99956 131228
rect 100588 131188 100628 131228
rect 102028 131188 102068 131228
rect 102124 131188 102164 131228
rect 102316 131188 102356 131228
rect 103180 131188 103220 131228
rect 103372 131188 103412 131228
rect 108940 131188 108980 131228
rect 109036 131188 109076 131228
rect 109132 131188 109172 131228
rect 109324 131188 109364 131228
rect 109420 131188 109460 131228
rect 109612 131188 109652 131228
rect 110476 131188 110516 131228
rect 111436 131188 111476 131228
rect 112492 131188 112532 131228
rect 112588 131188 112628 131228
rect 113068 131188 113108 131228
rect 113164 131188 113204 131228
rect 114892 131188 114932 131228
rect 114988 131188 115028 131228
rect 119116 131188 119156 131228
rect 119212 131188 119252 131228
rect 119404 131188 119444 131228
rect 104044 131020 104084 131060
rect 102508 130936 102548 130976
rect 115180 130936 115220 130976
rect 78184 130768 78224 130808
rect 78266 130768 78306 130808
rect 78348 130768 78388 130808
rect 78430 130768 78470 130808
rect 78512 130768 78552 130808
rect 93304 130768 93344 130808
rect 93386 130768 93426 130808
rect 93468 130768 93508 130808
rect 93550 130768 93590 130808
rect 93632 130768 93672 130808
rect 108424 130768 108464 130808
rect 108506 130768 108546 130808
rect 108588 130768 108628 130808
rect 108670 130768 108710 130808
rect 108752 130768 108792 130808
rect 123544 130768 123584 130808
rect 123626 130768 123666 130808
rect 123708 130768 123748 130808
rect 123790 130768 123830 130808
rect 123872 130768 123912 130808
rect 138664 130768 138704 130808
rect 138746 130768 138786 130808
rect 138828 130768 138868 130808
rect 138910 130768 138950 130808
rect 138992 130768 139032 130808
rect 98092 130600 98132 130640
rect 102604 130600 102644 130640
rect 110476 130600 110516 130640
rect 117580 130600 117620 130640
rect 103084 130516 103124 130556
rect 108748 130432 108788 130472
rect 97911 130337 97951 130377
rect 98092 130348 98132 130388
rect 102508 130348 102548 130388
rect 102796 130348 102836 130388
rect 102988 130348 103028 130388
rect 103084 130348 103124 130388
rect 105388 130348 105428 130388
rect 110188 130348 110228 130388
rect 110476 130348 110516 130388
rect 110668 130348 110708 130388
rect 110764 130348 110804 130388
rect 117484 130348 117524 130388
rect 117676 130348 117716 130388
rect 104716 130180 104756 130220
rect 79424 130012 79464 130052
rect 79506 130012 79546 130052
rect 79588 130012 79628 130052
rect 79670 130012 79710 130052
rect 79752 130012 79792 130052
rect 94544 130012 94584 130052
rect 94626 130012 94666 130052
rect 94708 130012 94748 130052
rect 94790 130012 94830 130052
rect 94872 130012 94912 130052
rect 109664 130012 109704 130052
rect 109746 130012 109786 130052
rect 109828 130012 109868 130052
rect 109910 130012 109950 130052
rect 109992 130012 110032 130052
rect 124784 130012 124824 130052
rect 124866 130012 124906 130052
rect 124948 130012 124988 130052
rect 125030 130012 125070 130052
rect 125112 130012 125152 130052
rect 139904 130012 139944 130052
rect 139986 130012 140026 130052
rect 140068 130012 140108 130052
rect 140150 130012 140190 130052
rect 140232 130012 140272 130052
rect 96844 129844 96884 129884
rect 97228 129844 97268 129884
rect 103180 129844 103220 129884
rect 105964 129844 106004 129884
rect 103564 129760 103604 129800
rect 96172 129676 96212 129716
rect 97132 129676 97172 129716
rect 97324 129676 97364 129716
rect 97420 129676 97460 129716
rect 103084 129676 103124 129716
rect 103276 129676 103316 129716
rect 103948 129676 103988 129716
rect 104812 129676 104852 129716
rect 110572 129676 110612 129716
rect 112012 129676 112052 129716
rect 113932 129676 113972 129716
rect 115372 129676 115412 129716
rect 78184 129256 78224 129296
rect 78266 129256 78306 129296
rect 78348 129256 78388 129296
rect 78430 129256 78470 129296
rect 78512 129256 78552 129296
rect 93304 129256 93344 129296
rect 93386 129256 93426 129296
rect 93468 129256 93508 129296
rect 93550 129256 93590 129296
rect 93632 129256 93672 129296
rect 108424 129256 108464 129296
rect 108506 129256 108546 129296
rect 108588 129256 108628 129296
rect 108670 129256 108710 129296
rect 108752 129256 108792 129296
rect 123544 129256 123584 129296
rect 123626 129256 123666 129296
rect 123708 129256 123748 129296
rect 123790 129256 123830 129296
rect 123872 129256 123912 129296
rect 138664 129256 138704 129296
rect 138746 129256 138786 129296
rect 138828 129256 138868 129296
rect 138910 129256 138950 129296
rect 138992 129256 139032 129296
rect 94156 129088 94196 129128
rect 96748 129088 96788 129128
rect 104044 129004 104084 129044
rect 121228 129004 121268 129044
rect 93868 128836 93908 128876
rect 93964 128836 94004 128876
rect 96076 128836 96116 128876
rect 119500 128836 119540 128876
rect 120364 128836 120404 128876
rect 121996 128836 122036 128876
rect 94060 128752 94100 128792
rect 94156 128668 94196 128708
rect 120172 128668 120212 128708
rect 121036 128668 121076 128708
rect 121900 128668 121940 128708
rect 79424 128500 79464 128540
rect 79506 128500 79546 128540
rect 79588 128500 79628 128540
rect 79670 128500 79710 128540
rect 79752 128500 79792 128540
rect 94544 128500 94584 128540
rect 94626 128500 94666 128540
rect 94708 128500 94748 128540
rect 94790 128500 94830 128540
rect 94872 128500 94912 128540
rect 109664 128500 109704 128540
rect 109746 128500 109786 128540
rect 109828 128500 109868 128540
rect 109910 128500 109950 128540
rect 109992 128500 110032 128540
rect 124784 128500 124824 128540
rect 124866 128500 124906 128540
rect 124948 128500 124988 128540
rect 125030 128500 125070 128540
rect 125112 128500 125152 128540
rect 139904 128500 139944 128540
rect 139986 128500 140026 128540
rect 140068 128500 140108 128540
rect 140150 128500 140190 128540
rect 140232 128500 140272 128540
rect 99148 128332 99188 128372
rect 119308 128332 119348 128372
rect 119788 128332 119828 128372
rect 123148 128332 123188 128372
rect 120748 128248 120788 128288
rect 99148 128164 99188 128204
rect 99244 128164 99284 128204
rect 118252 128164 118292 128204
rect 118444 128162 118484 128202
rect 118540 128164 118580 128204
rect 118636 128164 118676 128204
rect 119020 128164 119060 128204
rect 119116 128164 119156 128204
rect 119212 128164 119252 128204
rect 119596 128164 119636 128204
rect 119692 128164 119732 128204
rect 119884 128164 119924 128204
rect 121132 128164 121172 128204
rect 121996 128164 122036 128204
rect 99052 128080 99092 128120
rect 98956 127996 98996 128036
rect 118828 127912 118868 127952
rect 123148 127912 123188 127952
rect 78184 127744 78224 127784
rect 78266 127744 78306 127784
rect 78348 127744 78388 127784
rect 78430 127744 78470 127784
rect 78512 127744 78552 127784
rect 93304 127744 93344 127784
rect 93386 127744 93426 127784
rect 93468 127744 93508 127784
rect 93550 127744 93590 127784
rect 93632 127744 93672 127784
rect 108424 127744 108464 127784
rect 108506 127744 108546 127784
rect 108588 127744 108628 127784
rect 108670 127744 108710 127784
rect 108752 127744 108792 127784
rect 123544 127744 123584 127784
rect 123626 127744 123666 127784
rect 123708 127744 123748 127784
rect 123790 127744 123830 127784
rect 123872 127744 123912 127784
rect 138664 127744 138704 127784
rect 138746 127744 138786 127784
rect 138828 127744 138868 127784
rect 138910 127744 138950 127784
rect 138992 127744 139032 127784
rect 94828 127576 94868 127616
rect 94599 127324 94639 127364
rect 94712 127324 94752 127364
rect 94828 127324 94868 127364
rect 94924 127324 94964 127364
rect 118828 127324 118868 127364
rect 118924 127324 118964 127364
rect 119020 127324 119060 127364
rect 119116 127156 119156 127196
rect 79424 126988 79464 127028
rect 79506 126988 79546 127028
rect 79588 126988 79628 127028
rect 79670 126988 79710 127028
rect 79752 126988 79792 127028
rect 94544 126988 94584 127028
rect 94626 126988 94666 127028
rect 94708 126988 94748 127028
rect 94790 126988 94830 127028
rect 94872 126988 94912 127028
rect 109664 126988 109704 127028
rect 109746 126988 109786 127028
rect 109828 126988 109868 127028
rect 109910 126988 109950 127028
rect 109992 126988 110032 127028
rect 124784 126988 124824 127028
rect 124866 126988 124906 127028
rect 124948 126988 124988 127028
rect 125030 126988 125070 127028
rect 125112 126988 125152 127028
rect 139904 126988 139944 127028
rect 139986 126988 140026 127028
rect 140068 126988 140108 127028
rect 140150 126988 140190 127028
rect 140232 126988 140272 127028
rect 94636 126820 94676 126860
rect 95500 126820 95540 126860
rect 94732 126736 94772 126776
rect 94828 126652 94868 126692
rect 94924 126652 94964 126692
rect 95559 126652 95599 126692
rect 95672 126652 95712 126692
rect 95788 126652 95828 126692
rect 95884 126652 95924 126692
rect 94828 126400 94868 126440
rect 78184 126232 78224 126272
rect 78266 126232 78306 126272
rect 78348 126232 78388 126272
rect 78430 126232 78470 126272
rect 78512 126232 78552 126272
rect 93304 126232 93344 126272
rect 93386 126232 93426 126272
rect 93468 126232 93508 126272
rect 93550 126232 93590 126272
rect 93632 126232 93672 126272
rect 108424 126232 108464 126272
rect 108506 126232 108546 126272
rect 108588 126232 108628 126272
rect 108670 126232 108710 126272
rect 108752 126232 108792 126272
rect 123544 126232 123584 126272
rect 123626 126232 123666 126272
rect 123708 126232 123748 126272
rect 123790 126232 123830 126272
rect 123872 126232 123912 126272
rect 138664 126232 138704 126272
rect 138746 126232 138786 126272
rect 138828 126232 138868 126272
rect 138910 126232 138950 126272
rect 138992 126232 139032 126272
rect 119116 125812 119156 125852
rect 119212 125837 119252 125877
rect 119404 125728 119444 125768
rect 119116 125644 119156 125684
rect 79424 125476 79464 125516
rect 79506 125476 79546 125516
rect 79588 125476 79628 125516
rect 79670 125476 79710 125516
rect 79752 125476 79792 125516
rect 94544 125476 94584 125516
rect 94626 125476 94666 125516
rect 94708 125476 94748 125516
rect 94790 125476 94830 125516
rect 94872 125476 94912 125516
rect 109664 125476 109704 125516
rect 109746 125476 109786 125516
rect 109828 125476 109868 125516
rect 109910 125476 109950 125516
rect 109992 125476 110032 125516
rect 124784 125476 124824 125516
rect 124866 125476 124906 125516
rect 124948 125476 124988 125516
rect 125030 125476 125070 125516
rect 125112 125476 125152 125516
rect 139904 125476 139944 125516
rect 139986 125476 140026 125516
rect 140068 125476 140108 125516
rect 140150 125476 140190 125516
rect 140232 125476 140272 125516
rect 121036 125308 121076 125348
rect 121132 125140 121172 125180
rect 121516 125140 121556 125180
rect 122188 125140 122228 125180
rect 78184 124720 78224 124760
rect 78266 124720 78306 124760
rect 78348 124720 78388 124760
rect 78430 124720 78470 124760
rect 78512 124720 78552 124760
rect 93304 124720 93344 124760
rect 93386 124720 93426 124760
rect 93468 124720 93508 124760
rect 93550 124720 93590 124760
rect 93632 124720 93672 124760
rect 108424 124720 108464 124760
rect 108506 124720 108546 124760
rect 108588 124720 108628 124760
rect 108670 124720 108710 124760
rect 108752 124720 108792 124760
rect 123544 124720 123584 124760
rect 123626 124720 123666 124760
rect 123708 124720 123748 124760
rect 123790 124720 123830 124760
rect 123872 124720 123912 124760
rect 138664 124720 138704 124760
rect 138746 124720 138786 124760
rect 138828 124720 138868 124760
rect 138910 124720 138950 124760
rect 138992 124720 139032 124760
rect 79564 124552 79604 124592
rect 78892 124300 78932 124340
rect 79424 123964 79464 124004
rect 79506 123964 79546 124004
rect 79588 123964 79628 124004
rect 79670 123964 79710 124004
rect 79752 123964 79792 124004
rect 94544 123964 94584 124004
rect 94626 123964 94666 124004
rect 94708 123964 94748 124004
rect 94790 123964 94830 124004
rect 94872 123964 94912 124004
rect 109664 123964 109704 124004
rect 109746 123964 109786 124004
rect 109828 123964 109868 124004
rect 109910 123964 109950 124004
rect 109992 123964 110032 124004
rect 124784 123964 124824 124004
rect 124866 123964 124906 124004
rect 124948 123964 124988 124004
rect 125030 123964 125070 124004
rect 125112 123964 125152 124004
rect 139904 123964 139944 124004
rect 139986 123964 140026 124004
rect 140068 123964 140108 124004
rect 140150 123964 140190 124004
rect 140232 123964 140272 124004
rect 121612 123796 121652 123836
rect 119212 123712 119252 123752
rect 119596 123628 119636 123668
rect 120460 123628 120500 123668
rect 121612 123376 121652 123416
rect 78184 123208 78224 123248
rect 78266 123208 78306 123248
rect 78348 123208 78388 123248
rect 78430 123208 78470 123248
rect 78512 123208 78552 123248
rect 93304 123208 93344 123248
rect 93386 123208 93426 123248
rect 93468 123208 93508 123248
rect 93550 123208 93590 123248
rect 93632 123208 93672 123248
rect 108424 123208 108464 123248
rect 108506 123208 108546 123248
rect 108588 123208 108628 123248
rect 108670 123208 108710 123248
rect 108752 123208 108792 123248
rect 123544 123208 123584 123248
rect 123626 123208 123666 123248
rect 123708 123208 123748 123248
rect 123790 123208 123830 123248
rect 123872 123208 123912 123248
rect 138664 123208 138704 123248
rect 138746 123208 138786 123248
rect 138828 123208 138868 123248
rect 138910 123208 138950 123248
rect 138992 123208 139032 123248
rect 119692 122956 119732 122996
rect 79424 122452 79464 122492
rect 79506 122452 79546 122492
rect 79588 122452 79628 122492
rect 79670 122452 79710 122492
rect 79752 122452 79792 122492
rect 94544 122452 94584 122492
rect 94626 122452 94666 122492
rect 94708 122452 94748 122492
rect 94790 122452 94830 122492
rect 94872 122452 94912 122492
rect 109664 122452 109704 122492
rect 109746 122452 109786 122492
rect 109828 122452 109868 122492
rect 109910 122452 109950 122492
rect 109992 122452 110032 122492
rect 124784 122452 124824 122492
rect 124866 122452 124906 122492
rect 124948 122452 124988 122492
rect 125030 122452 125070 122492
rect 125112 122452 125152 122492
rect 139904 122452 139944 122492
rect 139986 122452 140026 122492
rect 140068 122452 140108 122492
rect 140150 122452 140190 122492
rect 140232 122452 140272 122492
rect 78184 121696 78224 121736
rect 78266 121696 78306 121736
rect 78348 121696 78388 121736
rect 78430 121696 78470 121736
rect 78512 121696 78552 121736
rect 93304 121696 93344 121736
rect 93386 121696 93426 121736
rect 93468 121696 93508 121736
rect 93550 121696 93590 121736
rect 93632 121696 93672 121736
rect 108424 121696 108464 121736
rect 108506 121696 108546 121736
rect 108588 121696 108628 121736
rect 108670 121696 108710 121736
rect 108752 121696 108792 121736
rect 123544 121696 123584 121736
rect 123626 121696 123666 121736
rect 123708 121696 123748 121736
rect 123790 121696 123830 121736
rect 123872 121696 123912 121736
rect 138664 121696 138704 121736
rect 138746 121696 138786 121736
rect 138828 121696 138868 121736
rect 138910 121696 138950 121736
rect 138992 121696 139032 121736
rect 79424 120940 79464 120980
rect 79506 120940 79546 120980
rect 79588 120940 79628 120980
rect 79670 120940 79710 120980
rect 79752 120940 79792 120980
rect 94544 120940 94584 120980
rect 94626 120940 94666 120980
rect 94708 120940 94748 120980
rect 94790 120940 94830 120980
rect 94872 120940 94912 120980
rect 109664 120940 109704 120980
rect 109746 120940 109786 120980
rect 109828 120940 109868 120980
rect 109910 120940 109950 120980
rect 109992 120940 110032 120980
rect 124784 120940 124824 120980
rect 124866 120940 124906 120980
rect 124948 120940 124988 120980
rect 125030 120940 125070 120980
rect 125112 120940 125152 120980
rect 139904 120940 139944 120980
rect 139986 120940 140026 120980
rect 140068 120940 140108 120980
rect 140150 120940 140190 120980
rect 140232 120940 140272 120980
rect 78184 120184 78224 120224
rect 78266 120184 78306 120224
rect 78348 120184 78388 120224
rect 78430 120184 78470 120224
rect 78512 120184 78552 120224
rect 93304 120184 93344 120224
rect 93386 120184 93426 120224
rect 93468 120184 93508 120224
rect 93550 120184 93590 120224
rect 93632 120184 93672 120224
rect 108424 120184 108464 120224
rect 108506 120184 108546 120224
rect 108588 120184 108628 120224
rect 108670 120184 108710 120224
rect 108752 120184 108792 120224
rect 123544 120184 123584 120224
rect 123626 120184 123666 120224
rect 123708 120184 123748 120224
rect 123790 120184 123830 120224
rect 123872 120184 123912 120224
rect 138664 120184 138704 120224
rect 138746 120184 138786 120224
rect 138828 120184 138868 120224
rect 138910 120184 138950 120224
rect 138992 120184 139032 120224
rect 79424 119428 79464 119468
rect 79506 119428 79546 119468
rect 79588 119428 79628 119468
rect 79670 119428 79710 119468
rect 79752 119428 79792 119468
rect 94544 119428 94584 119468
rect 94626 119428 94666 119468
rect 94708 119428 94748 119468
rect 94790 119428 94830 119468
rect 94872 119428 94912 119468
rect 109664 119428 109704 119468
rect 109746 119428 109786 119468
rect 109828 119428 109868 119468
rect 109910 119428 109950 119468
rect 109992 119428 110032 119468
rect 124784 119428 124824 119468
rect 124866 119428 124906 119468
rect 124948 119428 124988 119468
rect 125030 119428 125070 119468
rect 125112 119428 125152 119468
rect 139904 119428 139944 119468
rect 139986 119428 140026 119468
rect 140068 119428 140108 119468
rect 140150 119428 140190 119468
rect 140232 119428 140272 119468
rect 78184 118672 78224 118712
rect 78266 118672 78306 118712
rect 78348 118672 78388 118712
rect 78430 118672 78470 118712
rect 78512 118672 78552 118712
rect 93304 118672 93344 118712
rect 93386 118672 93426 118712
rect 93468 118672 93508 118712
rect 93550 118672 93590 118712
rect 93632 118672 93672 118712
rect 108424 118672 108464 118712
rect 108506 118672 108546 118712
rect 108588 118672 108628 118712
rect 108670 118672 108710 118712
rect 108752 118672 108792 118712
rect 123544 118672 123584 118712
rect 123626 118672 123666 118712
rect 123708 118672 123748 118712
rect 123790 118672 123830 118712
rect 123872 118672 123912 118712
rect 138664 118672 138704 118712
rect 138746 118672 138786 118712
rect 138828 118672 138868 118712
rect 138910 118672 138950 118712
rect 138992 118672 139032 118712
rect 79424 117916 79464 117956
rect 79506 117916 79546 117956
rect 79588 117916 79628 117956
rect 79670 117916 79710 117956
rect 79752 117916 79792 117956
rect 94544 117916 94584 117956
rect 94626 117916 94666 117956
rect 94708 117916 94748 117956
rect 94790 117916 94830 117956
rect 94872 117916 94912 117956
rect 109664 117916 109704 117956
rect 109746 117916 109786 117956
rect 109828 117916 109868 117956
rect 109910 117916 109950 117956
rect 109992 117916 110032 117956
rect 124784 117916 124824 117956
rect 124866 117916 124906 117956
rect 124948 117916 124988 117956
rect 125030 117916 125070 117956
rect 125112 117916 125152 117956
rect 139904 117916 139944 117956
rect 139986 117916 140026 117956
rect 140068 117916 140108 117956
rect 140150 117916 140190 117956
rect 140232 117916 140272 117956
rect 78184 117160 78224 117200
rect 78266 117160 78306 117200
rect 78348 117160 78388 117200
rect 78430 117160 78470 117200
rect 78512 117160 78552 117200
rect 93304 117160 93344 117200
rect 93386 117160 93426 117200
rect 93468 117160 93508 117200
rect 93550 117160 93590 117200
rect 93632 117160 93672 117200
rect 108424 117160 108464 117200
rect 108506 117160 108546 117200
rect 108588 117160 108628 117200
rect 108670 117160 108710 117200
rect 108752 117160 108792 117200
rect 123544 117160 123584 117200
rect 123626 117160 123666 117200
rect 123708 117160 123748 117200
rect 123790 117160 123830 117200
rect 123872 117160 123912 117200
rect 138664 117160 138704 117200
rect 138746 117160 138786 117200
rect 138828 117160 138868 117200
rect 138910 117160 138950 117200
rect 138992 117160 139032 117200
rect 79424 116404 79464 116444
rect 79506 116404 79546 116444
rect 79588 116404 79628 116444
rect 79670 116404 79710 116444
rect 79752 116404 79792 116444
rect 94544 116404 94584 116444
rect 94626 116404 94666 116444
rect 94708 116404 94748 116444
rect 94790 116404 94830 116444
rect 94872 116404 94912 116444
rect 109664 116404 109704 116444
rect 109746 116404 109786 116444
rect 109828 116404 109868 116444
rect 109910 116404 109950 116444
rect 109992 116404 110032 116444
rect 124784 116404 124824 116444
rect 124866 116404 124906 116444
rect 124948 116404 124988 116444
rect 125030 116404 125070 116444
rect 125112 116404 125152 116444
rect 139904 116404 139944 116444
rect 139986 116404 140026 116444
rect 140068 116404 140108 116444
rect 140150 116404 140190 116444
rect 140232 116404 140272 116444
rect 78184 115648 78224 115688
rect 78266 115648 78306 115688
rect 78348 115648 78388 115688
rect 78430 115648 78470 115688
rect 78512 115648 78552 115688
rect 93304 115648 93344 115688
rect 93386 115648 93426 115688
rect 93468 115648 93508 115688
rect 93550 115648 93590 115688
rect 93632 115648 93672 115688
rect 108424 115648 108464 115688
rect 108506 115648 108546 115688
rect 108588 115648 108628 115688
rect 108670 115648 108710 115688
rect 108752 115648 108792 115688
rect 123544 115648 123584 115688
rect 123626 115648 123666 115688
rect 123708 115648 123748 115688
rect 123790 115648 123830 115688
rect 123872 115648 123912 115688
rect 138664 115648 138704 115688
rect 138746 115648 138786 115688
rect 138828 115648 138868 115688
rect 138910 115648 138950 115688
rect 138992 115648 139032 115688
rect 79424 114892 79464 114932
rect 79506 114892 79546 114932
rect 79588 114892 79628 114932
rect 79670 114892 79710 114932
rect 79752 114892 79792 114932
rect 94544 114892 94584 114932
rect 94626 114892 94666 114932
rect 94708 114892 94748 114932
rect 94790 114892 94830 114932
rect 94872 114892 94912 114932
rect 109664 114892 109704 114932
rect 109746 114892 109786 114932
rect 109828 114892 109868 114932
rect 109910 114892 109950 114932
rect 109992 114892 110032 114932
rect 124784 114892 124824 114932
rect 124866 114892 124906 114932
rect 124948 114892 124988 114932
rect 125030 114892 125070 114932
rect 125112 114892 125152 114932
rect 139904 114892 139944 114932
rect 139986 114892 140026 114932
rect 140068 114892 140108 114932
rect 140150 114892 140190 114932
rect 140232 114892 140272 114932
rect 78184 114136 78224 114176
rect 78266 114136 78306 114176
rect 78348 114136 78388 114176
rect 78430 114136 78470 114176
rect 78512 114136 78552 114176
rect 93304 114136 93344 114176
rect 93386 114136 93426 114176
rect 93468 114136 93508 114176
rect 93550 114136 93590 114176
rect 93632 114136 93672 114176
rect 108424 114136 108464 114176
rect 108506 114136 108546 114176
rect 108588 114136 108628 114176
rect 108670 114136 108710 114176
rect 108752 114136 108792 114176
rect 123544 114136 123584 114176
rect 123626 114136 123666 114176
rect 123708 114136 123748 114176
rect 123790 114136 123830 114176
rect 123872 114136 123912 114176
rect 138664 114136 138704 114176
rect 138746 114136 138786 114176
rect 138828 114136 138868 114176
rect 138910 114136 138950 114176
rect 138992 114136 139032 114176
rect 79424 113380 79464 113420
rect 79506 113380 79546 113420
rect 79588 113380 79628 113420
rect 79670 113380 79710 113420
rect 79752 113380 79792 113420
rect 94544 113380 94584 113420
rect 94626 113380 94666 113420
rect 94708 113380 94748 113420
rect 94790 113380 94830 113420
rect 94872 113380 94912 113420
rect 109664 113380 109704 113420
rect 109746 113380 109786 113420
rect 109828 113380 109868 113420
rect 109910 113380 109950 113420
rect 109992 113380 110032 113420
rect 124784 113380 124824 113420
rect 124866 113380 124906 113420
rect 124948 113380 124988 113420
rect 125030 113380 125070 113420
rect 125112 113380 125152 113420
rect 139904 113380 139944 113420
rect 139986 113380 140026 113420
rect 140068 113380 140108 113420
rect 140150 113380 140190 113420
rect 140232 113380 140272 113420
rect 78184 112624 78224 112664
rect 78266 112624 78306 112664
rect 78348 112624 78388 112664
rect 78430 112624 78470 112664
rect 78512 112624 78552 112664
rect 93304 112624 93344 112664
rect 93386 112624 93426 112664
rect 93468 112624 93508 112664
rect 93550 112624 93590 112664
rect 93632 112624 93672 112664
rect 108424 112624 108464 112664
rect 108506 112624 108546 112664
rect 108588 112624 108628 112664
rect 108670 112624 108710 112664
rect 108752 112624 108792 112664
rect 123544 112624 123584 112664
rect 123626 112624 123666 112664
rect 123708 112624 123748 112664
rect 123790 112624 123830 112664
rect 123872 112624 123912 112664
rect 138664 112624 138704 112664
rect 138746 112624 138786 112664
rect 138828 112624 138868 112664
rect 138910 112624 138950 112664
rect 138992 112624 139032 112664
rect 79424 111868 79464 111908
rect 79506 111868 79546 111908
rect 79588 111868 79628 111908
rect 79670 111868 79710 111908
rect 79752 111868 79792 111908
rect 94544 111868 94584 111908
rect 94626 111868 94666 111908
rect 94708 111868 94748 111908
rect 94790 111868 94830 111908
rect 94872 111868 94912 111908
rect 109664 111868 109704 111908
rect 109746 111868 109786 111908
rect 109828 111868 109868 111908
rect 109910 111868 109950 111908
rect 109992 111868 110032 111908
rect 124784 111868 124824 111908
rect 124866 111868 124906 111908
rect 124948 111868 124988 111908
rect 125030 111868 125070 111908
rect 125112 111868 125152 111908
rect 139904 111868 139944 111908
rect 139986 111868 140026 111908
rect 140068 111868 140108 111908
rect 140150 111868 140190 111908
rect 140232 111868 140272 111908
rect 78184 111112 78224 111152
rect 78266 111112 78306 111152
rect 78348 111112 78388 111152
rect 78430 111112 78470 111152
rect 78512 111112 78552 111152
rect 93304 111112 93344 111152
rect 93386 111112 93426 111152
rect 93468 111112 93508 111152
rect 93550 111112 93590 111152
rect 93632 111112 93672 111152
rect 108424 111112 108464 111152
rect 108506 111112 108546 111152
rect 108588 111112 108628 111152
rect 108670 111112 108710 111152
rect 108752 111112 108792 111152
rect 123544 111112 123584 111152
rect 123626 111112 123666 111152
rect 123708 111112 123748 111152
rect 123790 111112 123830 111152
rect 123872 111112 123912 111152
rect 138664 111112 138704 111152
rect 138746 111112 138786 111152
rect 138828 111112 138868 111152
rect 138910 111112 138950 111152
rect 138992 111112 139032 111152
rect 79424 110356 79464 110396
rect 79506 110356 79546 110396
rect 79588 110356 79628 110396
rect 79670 110356 79710 110396
rect 79752 110356 79792 110396
rect 94544 110356 94584 110396
rect 94626 110356 94666 110396
rect 94708 110356 94748 110396
rect 94790 110356 94830 110396
rect 94872 110356 94912 110396
rect 109664 110356 109704 110396
rect 109746 110356 109786 110396
rect 109828 110356 109868 110396
rect 109910 110356 109950 110396
rect 109992 110356 110032 110396
rect 124784 110356 124824 110396
rect 124866 110356 124906 110396
rect 124948 110356 124988 110396
rect 125030 110356 125070 110396
rect 125112 110356 125152 110396
rect 139904 110356 139944 110396
rect 139986 110356 140026 110396
rect 140068 110356 140108 110396
rect 140150 110356 140190 110396
rect 140232 110356 140272 110396
rect 78184 109600 78224 109640
rect 78266 109600 78306 109640
rect 78348 109600 78388 109640
rect 78430 109600 78470 109640
rect 78512 109600 78552 109640
rect 93304 109600 93344 109640
rect 93386 109600 93426 109640
rect 93468 109600 93508 109640
rect 93550 109600 93590 109640
rect 93632 109600 93672 109640
rect 108424 109600 108464 109640
rect 108506 109600 108546 109640
rect 108588 109600 108628 109640
rect 108670 109600 108710 109640
rect 108752 109600 108792 109640
rect 123544 109600 123584 109640
rect 123626 109600 123666 109640
rect 123708 109600 123748 109640
rect 123790 109600 123830 109640
rect 123872 109600 123912 109640
rect 138664 109600 138704 109640
rect 138746 109600 138786 109640
rect 138828 109600 138868 109640
rect 138910 109600 138950 109640
rect 138992 109600 139032 109640
rect 79424 108844 79464 108884
rect 79506 108844 79546 108884
rect 79588 108844 79628 108884
rect 79670 108844 79710 108884
rect 79752 108844 79792 108884
rect 94544 108844 94584 108884
rect 94626 108844 94666 108884
rect 94708 108844 94748 108884
rect 94790 108844 94830 108884
rect 94872 108844 94912 108884
rect 109664 108844 109704 108884
rect 109746 108844 109786 108884
rect 109828 108844 109868 108884
rect 109910 108844 109950 108884
rect 109992 108844 110032 108884
rect 124784 108844 124824 108884
rect 124866 108844 124906 108884
rect 124948 108844 124988 108884
rect 125030 108844 125070 108884
rect 125112 108844 125152 108884
rect 139904 108844 139944 108884
rect 139986 108844 140026 108884
rect 140068 108844 140108 108884
rect 140150 108844 140190 108884
rect 140232 108844 140272 108884
rect 78184 108088 78224 108128
rect 78266 108088 78306 108128
rect 78348 108088 78388 108128
rect 78430 108088 78470 108128
rect 78512 108088 78552 108128
rect 93304 108088 93344 108128
rect 93386 108088 93426 108128
rect 93468 108088 93508 108128
rect 93550 108088 93590 108128
rect 93632 108088 93672 108128
rect 108424 108088 108464 108128
rect 108506 108088 108546 108128
rect 108588 108088 108628 108128
rect 108670 108088 108710 108128
rect 108752 108088 108792 108128
rect 123544 108088 123584 108128
rect 123626 108088 123666 108128
rect 123708 108088 123748 108128
rect 123790 108088 123830 108128
rect 123872 108088 123912 108128
rect 138664 108088 138704 108128
rect 138746 108088 138786 108128
rect 138828 108088 138868 108128
rect 138910 108088 138950 108128
rect 138992 108088 139032 108128
rect 79424 107332 79464 107372
rect 79506 107332 79546 107372
rect 79588 107332 79628 107372
rect 79670 107332 79710 107372
rect 79752 107332 79792 107372
rect 94544 107332 94584 107372
rect 94626 107332 94666 107372
rect 94708 107332 94748 107372
rect 94790 107332 94830 107372
rect 94872 107332 94912 107372
rect 109664 107332 109704 107372
rect 109746 107332 109786 107372
rect 109828 107332 109868 107372
rect 109910 107332 109950 107372
rect 109992 107332 110032 107372
rect 124784 107332 124824 107372
rect 124866 107332 124906 107372
rect 124948 107332 124988 107372
rect 125030 107332 125070 107372
rect 125112 107332 125152 107372
rect 139904 107332 139944 107372
rect 139986 107332 140026 107372
rect 140068 107332 140108 107372
rect 140150 107332 140190 107372
rect 140232 107332 140272 107372
rect 78184 106576 78224 106616
rect 78266 106576 78306 106616
rect 78348 106576 78388 106616
rect 78430 106576 78470 106616
rect 78512 106576 78552 106616
rect 93304 106576 93344 106616
rect 93386 106576 93426 106616
rect 93468 106576 93508 106616
rect 93550 106576 93590 106616
rect 93632 106576 93672 106616
rect 108424 106576 108464 106616
rect 108506 106576 108546 106616
rect 108588 106576 108628 106616
rect 108670 106576 108710 106616
rect 108752 106576 108792 106616
rect 123544 106576 123584 106616
rect 123626 106576 123666 106616
rect 123708 106576 123748 106616
rect 123790 106576 123830 106616
rect 123872 106576 123912 106616
rect 138664 106576 138704 106616
rect 138746 106576 138786 106616
rect 138828 106576 138868 106616
rect 138910 106576 138950 106616
rect 138992 106576 139032 106616
rect 79424 105820 79464 105860
rect 79506 105820 79546 105860
rect 79588 105820 79628 105860
rect 79670 105820 79710 105860
rect 79752 105820 79792 105860
rect 94544 105820 94584 105860
rect 94626 105820 94666 105860
rect 94708 105820 94748 105860
rect 94790 105820 94830 105860
rect 94872 105820 94912 105860
rect 109664 105820 109704 105860
rect 109746 105820 109786 105860
rect 109828 105820 109868 105860
rect 109910 105820 109950 105860
rect 109992 105820 110032 105860
rect 124784 105820 124824 105860
rect 124866 105820 124906 105860
rect 124948 105820 124988 105860
rect 125030 105820 125070 105860
rect 125112 105820 125152 105860
rect 139904 105820 139944 105860
rect 139986 105820 140026 105860
rect 140068 105820 140108 105860
rect 140150 105820 140190 105860
rect 140232 105820 140272 105860
rect 78184 105064 78224 105104
rect 78266 105064 78306 105104
rect 78348 105064 78388 105104
rect 78430 105064 78470 105104
rect 78512 105064 78552 105104
rect 93304 105064 93344 105104
rect 93386 105064 93426 105104
rect 93468 105064 93508 105104
rect 93550 105064 93590 105104
rect 93632 105064 93672 105104
rect 108424 105064 108464 105104
rect 108506 105064 108546 105104
rect 108588 105064 108628 105104
rect 108670 105064 108710 105104
rect 108752 105064 108792 105104
rect 123544 105064 123584 105104
rect 123626 105064 123666 105104
rect 123708 105064 123748 105104
rect 123790 105064 123830 105104
rect 123872 105064 123912 105104
rect 138664 105064 138704 105104
rect 138746 105064 138786 105104
rect 138828 105064 138868 105104
rect 138910 105064 138950 105104
rect 138992 105064 139032 105104
rect 79424 104308 79464 104348
rect 79506 104308 79546 104348
rect 79588 104308 79628 104348
rect 79670 104308 79710 104348
rect 79752 104308 79792 104348
rect 94544 104308 94584 104348
rect 94626 104308 94666 104348
rect 94708 104308 94748 104348
rect 94790 104308 94830 104348
rect 94872 104308 94912 104348
rect 109664 104308 109704 104348
rect 109746 104308 109786 104348
rect 109828 104308 109868 104348
rect 109910 104308 109950 104348
rect 109992 104308 110032 104348
rect 124784 104308 124824 104348
rect 124866 104308 124906 104348
rect 124948 104308 124988 104348
rect 125030 104308 125070 104348
rect 125112 104308 125152 104348
rect 139904 104308 139944 104348
rect 139986 104308 140026 104348
rect 140068 104308 140108 104348
rect 140150 104308 140190 104348
rect 140232 104308 140272 104348
rect 78184 103552 78224 103592
rect 78266 103552 78306 103592
rect 78348 103552 78388 103592
rect 78430 103552 78470 103592
rect 78512 103552 78552 103592
rect 93304 103552 93344 103592
rect 93386 103552 93426 103592
rect 93468 103552 93508 103592
rect 93550 103552 93590 103592
rect 93632 103552 93672 103592
rect 108424 103552 108464 103592
rect 108506 103552 108546 103592
rect 108588 103552 108628 103592
rect 108670 103552 108710 103592
rect 108752 103552 108792 103592
rect 123544 103552 123584 103592
rect 123626 103552 123666 103592
rect 123708 103552 123748 103592
rect 123790 103552 123830 103592
rect 123872 103552 123912 103592
rect 138664 103552 138704 103592
rect 138746 103552 138786 103592
rect 138828 103552 138868 103592
rect 138910 103552 138950 103592
rect 138992 103552 139032 103592
rect 79424 102796 79464 102836
rect 79506 102796 79546 102836
rect 79588 102796 79628 102836
rect 79670 102796 79710 102836
rect 79752 102796 79792 102836
rect 94544 102796 94584 102836
rect 94626 102796 94666 102836
rect 94708 102796 94748 102836
rect 94790 102796 94830 102836
rect 94872 102796 94912 102836
rect 109664 102796 109704 102836
rect 109746 102796 109786 102836
rect 109828 102796 109868 102836
rect 109910 102796 109950 102836
rect 109992 102796 110032 102836
rect 124784 102796 124824 102836
rect 124866 102796 124906 102836
rect 124948 102796 124988 102836
rect 125030 102796 125070 102836
rect 125112 102796 125152 102836
rect 139904 102796 139944 102836
rect 139986 102796 140026 102836
rect 140068 102796 140108 102836
rect 140150 102796 140190 102836
rect 140232 102796 140272 102836
rect 78184 102040 78224 102080
rect 78266 102040 78306 102080
rect 78348 102040 78388 102080
rect 78430 102040 78470 102080
rect 78512 102040 78552 102080
rect 93304 102040 93344 102080
rect 93386 102040 93426 102080
rect 93468 102040 93508 102080
rect 93550 102040 93590 102080
rect 93632 102040 93672 102080
rect 108424 102040 108464 102080
rect 108506 102040 108546 102080
rect 108588 102040 108628 102080
rect 108670 102040 108710 102080
rect 108752 102040 108792 102080
rect 123544 102040 123584 102080
rect 123626 102040 123666 102080
rect 123708 102040 123748 102080
rect 123790 102040 123830 102080
rect 123872 102040 123912 102080
rect 138664 102040 138704 102080
rect 138746 102040 138786 102080
rect 138828 102040 138868 102080
rect 138910 102040 138950 102080
rect 138992 102040 139032 102080
rect 79424 101284 79464 101324
rect 79506 101284 79546 101324
rect 79588 101284 79628 101324
rect 79670 101284 79710 101324
rect 79752 101284 79792 101324
rect 94544 101284 94584 101324
rect 94626 101284 94666 101324
rect 94708 101284 94748 101324
rect 94790 101284 94830 101324
rect 94872 101284 94912 101324
rect 109664 101284 109704 101324
rect 109746 101284 109786 101324
rect 109828 101284 109868 101324
rect 109910 101284 109950 101324
rect 109992 101284 110032 101324
rect 124784 101284 124824 101324
rect 124866 101284 124906 101324
rect 124948 101284 124988 101324
rect 125030 101284 125070 101324
rect 125112 101284 125152 101324
rect 139904 101284 139944 101324
rect 139986 101284 140026 101324
rect 140068 101284 140108 101324
rect 140150 101284 140190 101324
rect 140232 101284 140272 101324
rect 78184 100528 78224 100568
rect 78266 100528 78306 100568
rect 78348 100528 78388 100568
rect 78430 100528 78470 100568
rect 78512 100528 78552 100568
rect 93304 100528 93344 100568
rect 93386 100528 93426 100568
rect 93468 100528 93508 100568
rect 93550 100528 93590 100568
rect 93632 100528 93672 100568
rect 108424 100528 108464 100568
rect 108506 100528 108546 100568
rect 108588 100528 108628 100568
rect 108670 100528 108710 100568
rect 108752 100528 108792 100568
rect 123544 100528 123584 100568
rect 123626 100528 123666 100568
rect 123708 100528 123748 100568
rect 123790 100528 123830 100568
rect 123872 100528 123912 100568
rect 138664 100528 138704 100568
rect 138746 100528 138786 100568
rect 138828 100528 138868 100568
rect 138910 100528 138950 100568
rect 138992 100528 139032 100568
rect 79424 99772 79464 99812
rect 79506 99772 79546 99812
rect 79588 99772 79628 99812
rect 79670 99772 79710 99812
rect 79752 99772 79792 99812
rect 94544 99772 94584 99812
rect 94626 99772 94666 99812
rect 94708 99772 94748 99812
rect 94790 99772 94830 99812
rect 94872 99772 94912 99812
rect 109664 99772 109704 99812
rect 109746 99772 109786 99812
rect 109828 99772 109868 99812
rect 109910 99772 109950 99812
rect 109992 99772 110032 99812
rect 124784 99772 124824 99812
rect 124866 99772 124906 99812
rect 124948 99772 124988 99812
rect 125030 99772 125070 99812
rect 125112 99772 125152 99812
rect 139904 99772 139944 99812
rect 139986 99772 140026 99812
rect 140068 99772 140108 99812
rect 140150 99772 140190 99812
rect 140232 99772 140272 99812
rect 78184 99016 78224 99056
rect 78266 99016 78306 99056
rect 78348 99016 78388 99056
rect 78430 99016 78470 99056
rect 78512 99016 78552 99056
rect 93304 99016 93344 99056
rect 93386 99016 93426 99056
rect 93468 99016 93508 99056
rect 93550 99016 93590 99056
rect 93632 99016 93672 99056
rect 108424 99016 108464 99056
rect 108506 99016 108546 99056
rect 108588 99016 108628 99056
rect 108670 99016 108710 99056
rect 108752 99016 108792 99056
rect 123544 99016 123584 99056
rect 123626 99016 123666 99056
rect 123708 99016 123748 99056
rect 123790 99016 123830 99056
rect 123872 99016 123912 99056
rect 138664 99016 138704 99056
rect 138746 99016 138786 99056
rect 138828 99016 138868 99056
rect 138910 99016 138950 99056
rect 138992 99016 139032 99056
rect 79424 98260 79464 98300
rect 79506 98260 79546 98300
rect 79588 98260 79628 98300
rect 79670 98260 79710 98300
rect 79752 98260 79792 98300
rect 94544 98260 94584 98300
rect 94626 98260 94666 98300
rect 94708 98260 94748 98300
rect 94790 98260 94830 98300
rect 94872 98260 94912 98300
rect 109664 98260 109704 98300
rect 109746 98260 109786 98300
rect 109828 98260 109868 98300
rect 109910 98260 109950 98300
rect 109992 98260 110032 98300
rect 124784 98260 124824 98300
rect 124866 98260 124906 98300
rect 124948 98260 124988 98300
rect 125030 98260 125070 98300
rect 125112 98260 125152 98300
rect 139904 98260 139944 98300
rect 139986 98260 140026 98300
rect 140068 98260 140108 98300
rect 140150 98260 140190 98300
rect 140232 98260 140272 98300
rect 78184 97504 78224 97544
rect 78266 97504 78306 97544
rect 78348 97504 78388 97544
rect 78430 97504 78470 97544
rect 78512 97504 78552 97544
rect 93304 97504 93344 97544
rect 93386 97504 93426 97544
rect 93468 97504 93508 97544
rect 93550 97504 93590 97544
rect 93632 97504 93672 97544
rect 108424 97504 108464 97544
rect 108506 97504 108546 97544
rect 108588 97504 108628 97544
rect 108670 97504 108710 97544
rect 108752 97504 108792 97544
rect 123544 97504 123584 97544
rect 123626 97504 123666 97544
rect 123708 97504 123748 97544
rect 123790 97504 123830 97544
rect 123872 97504 123912 97544
rect 138664 97504 138704 97544
rect 138746 97504 138786 97544
rect 138828 97504 138868 97544
rect 138910 97504 138950 97544
rect 138992 97504 139032 97544
rect 79424 96748 79464 96788
rect 79506 96748 79546 96788
rect 79588 96748 79628 96788
rect 79670 96748 79710 96788
rect 79752 96748 79792 96788
rect 94544 96748 94584 96788
rect 94626 96748 94666 96788
rect 94708 96748 94748 96788
rect 94790 96748 94830 96788
rect 94872 96748 94912 96788
rect 109664 96748 109704 96788
rect 109746 96748 109786 96788
rect 109828 96748 109868 96788
rect 109910 96748 109950 96788
rect 109992 96748 110032 96788
rect 124784 96748 124824 96788
rect 124866 96748 124906 96788
rect 124948 96748 124988 96788
rect 125030 96748 125070 96788
rect 125112 96748 125152 96788
rect 139904 96748 139944 96788
rect 139986 96748 140026 96788
rect 140068 96748 140108 96788
rect 140150 96748 140190 96788
rect 140232 96748 140272 96788
rect 78184 95992 78224 96032
rect 78266 95992 78306 96032
rect 78348 95992 78388 96032
rect 78430 95992 78470 96032
rect 78512 95992 78552 96032
rect 93304 95992 93344 96032
rect 93386 95992 93426 96032
rect 93468 95992 93508 96032
rect 93550 95992 93590 96032
rect 93632 95992 93672 96032
rect 108424 95992 108464 96032
rect 108506 95992 108546 96032
rect 108588 95992 108628 96032
rect 108670 95992 108710 96032
rect 108752 95992 108792 96032
rect 123544 95992 123584 96032
rect 123626 95992 123666 96032
rect 123708 95992 123748 96032
rect 123790 95992 123830 96032
rect 123872 95992 123912 96032
rect 138664 95992 138704 96032
rect 138746 95992 138786 96032
rect 138828 95992 138868 96032
rect 138910 95992 138950 96032
rect 138992 95992 139032 96032
rect 104332 95824 104372 95864
rect 103660 95572 103700 95612
rect 79424 95236 79464 95276
rect 79506 95236 79546 95276
rect 79588 95236 79628 95276
rect 79670 95236 79710 95276
rect 79752 95236 79792 95276
rect 94544 95236 94584 95276
rect 94626 95236 94666 95276
rect 94708 95236 94748 95276
rect 94790 95236 94830 95276
rect 94872 95236 94912 95276
rect 109664 95236 109704 95276
rect 109746 95236 109786 95276
rect 109828 95236 109868 95276
rect 109910 95236 109950 95276
rect 109992 95236 110032 95276
rect 124784 95236 124824 95276
rect 124866 95236 124906 95276
rect 124948 95236 124988 95276
rect 125030 95236 125070 95276
rect 125112 95236 125152 95276
rect 139904 95236 139944 95276
rect 139986 95236 140026 95276
rect 140068 95236 140108 95276
rect 140150 95236 140190 95276
rect 140232 95236 140272 95276
rect 78184 94480 78224 94520
rect 78266 94480 78306 94520
rect 78348 94480 78388 94520
rect 78430 94480 78470 94520
rect 78512 94480 78552 94520
rect 93304 94480 93344 94520
rect 93386 94480 93426 94520
rect 93468 94480 93508 94520
rect 93550 94480 93590 94520
rect 93632 94480 93672 94520
rect 108424 94480 108464 94520
rect 108506 94480 108546 94520
rect 108588 94480 108628 94520
rect 108670 94480 108710 94520
rect 108752 94480 108792 94520
rect 123544 94480 123584 94520
rect 123626 94480 123666 94520
rect 123708 94480 123748 94520
rect 123790 94480 123830 94520
rect 123872 94480 123912 94520
rect 138664 94480 138704 94520
rect 138746 94480 138786 94520
rect 138828 94480 138868 94520
rect 138910 94480 138950 94520
rect 138992 94480 139032 94520
rect 79424 93724 79464 93764
rect 79506 93724 79546 93764
rect 79588 93724 79628 93764
rect 79670 93724 79710 93764
rect 79752 93724 79792 93764
rect 94544 93724 94584 93764
rect 94626 93724 94666 93764
rect 94708 93724 94748 93764
rect 94790 93724 94830 93764
rect 94872 93724 94912 93764
rect 109664 93724 109704 93764
rect 109746 93724 109786 93764
rect 109828 93724 109868 93764
rect 109910 93724 109950 93764
rect 109992 93724 110032 93764
rect 124784 93724 124824 93764
rect 124866 93724 124906 93764
rect 124948 93724 124988 93764
rect 125030 93724 125070 93764
rect 125112 93724 125152 93764
rect 139904 93724 139944 93764
rect 139986 93724 140026 93764
rect 140068 93724 140108 93764
rect 140150 93724 140190 93764
rect 140232 93724 140272 93764
rect 78184 92968 78224 93008
rect 78266 92968 78306 93008
rect 78348 92968 78388 93008
rect 78430 92968 78470 93008
rect 78512 92968 78552 93008
rect 93304 92968 93344 93008
rect 93386 92968 93426 93008
rect 93468 92968 93508 93008
rect 93550 92968 93590 93008
rect 93632 92968 93672 93008
rect 108424 92968 108464 93008
rect 108506 92968 108546 93008
rect 108588 92968 108628 93008
rect 108670 92968 108710 93008
rect 108752 92968 108792 93008
rect 123544 92968 123584 93008
rect 123626 92968 123666 93008
rect 123708 92968 123748 93008
rect 123790 92968 123830 93008
rect 123872 92968 123912 93008
rect 138664 92968 138704 93008
rect 138746 92968 138786 93008
rect 138828 92968 138868 93008
rect 138910 92968 138950 93008
rect 138992 92968 139032 93008
rect 79424 92212 79464 92252
rect 79506 92212 79546 92252
rect 79588 92212 79628 92252
rect 79670 92212 79710 92252
rect 79752 92212 79792 92252
rect 94544 92212 94584 92252
rect 94626 92212 94666 92252
rect 94708 92212 94748 92252
rect 94790 92212 94830 92252
rect 94872 92212 94912 92252
rect 109664 92212 109704 92252
rect 109746 92212 109786 92252
rect 109828 92212 109868 92252
rect 109910 92212 109950 92252
rect 109992 92212 110032 92252
rect 124784 92212 124824 92252
rect 124866 92212 124906 92252
rect 124948 92212 124988 92252
rect 125030 92212 125070 92252
rect 125112 92212 125152 92252
rect 139904 92212 139944 92252
rect 139986 92212 140026 92252
rect 140068 92212 140108 92252
rect 140150 92212 140190 92252
rect 140232 92212 140272 92252
rect 78184 91456 78224 91496
rect 78266 91456 78306 91496
rect 78348 91456 78388 91496
rect 78430 91456 78470 91496
rect 78512 91456 78552 91496
rect 93304 91456 93344 91496
rect 93386 91456 93426 91496
rect 93468 91456 93508 91496
rect 93550 91456 93590 91496
rect 93632 91456 93672 91496
rect 108424 91456 108464 91496
rect 108506 91456 108546 91496
rect 108588 91456 108628 91496
rect 108670 91456 108710 91496
rect 108752 91456 108792 91496
rect 123544 91456 123584 91496
rect 123626 91456 123666 91496
rect 123708 91456 123748 91496
rect 123790 91456 123830 91496
rect 123872 91456 123912 91496
rect 138664 91456 138704 91496
rect 138746 91456 138786 91496
rect 138828 91456 138868 91496
rect 138910 91456 138950 91496
rect 138992 91456 139032 91496
rect 79424 90700 79464 90740
rect 79506 90700 79546 90740
rect 79588 90700 79628 90740
rect 79670 90700 79710 90740
rect 79752 90700 79792 90740
rect 94544 90700 94584 90740
rect 94626 90700 94666 90740
rect 94708 90700 94748 90740
rect 94790 90700 94830 90740
rect 94872 90700 94912 90740
rect 109664 90700 109704 90740
rect 109746 90700 109786 90740
rect 109828 90700 109868 90740
rect 109910 90700 109950 90740
rect 109992 90700 110032 90740
rect 124784 90700 124824 90740
rect 124866 90700 124906 90740
rect 124948 90700 124988 90740
rect 125030 90700 125070 90740
rect 125112 90700 125152 90740
rect 139904 90700 139944 90740
rect 139986 90700 140026 90740
rect 140068 90700 140108 90740
rect 140150 90700 140190 90740
rect 140232 90700 140272 90740
rect 78184 89944 78224 89984
rect 78266 89944 78306 89984
rect 78348 89944 78388 89984
rect 78430 89944 78470 89984
rect 78512 89944 78552 89984
rect 93304 89944 93344 89984
rect 93386 89944 93426 89984
rect 93468 89944 93508 89984
rect 93550 89944 93590 89984
rect 93632 89944 93672 89984
rect 108424 89944 108464 89984
rect 108506 89944 108546 89984
rect 108588 89944 108628 89984
rect 108670 89944 108710 89984
rect 108752 89944 108792 89984
rect 123544 89944 123584 89984
rect 123626 89944 123666 89984
rect 123708 89944 123748 89984
rect 123790 89944 123830 89984
rect 123872 89944 123912 89984
rect 138664 89944 138704 89984
rect 138746 89944 138786 89984
rect 138828 89944 138868 89984
rect 138910 89944 138950 89984
rect 138992 89944 139032 89984
rect 79424 89188 79464 89228
rect 79506 89188 79546 89228
rect 79588 89188 79628 89228
rect 79670 89188 79710 89228
rect 79752 89188 79792 89228
rect 94544 89188 94584 89228
rect 94626 89188 94666 89228
rect 94708 89188 94748 89228
rect 94790 89188 94830 89228
rect 94872 89188 94912 89228
rect 109664 89188 109704 89228
rect 109746 89188 109786 89228
rect 109828 89188 109868 89228
rect 109910 89188 109950 89228
rect 109992 89188 110032 89228
rect 124784 89188 124824 89228
rect 124866 89188 124906 89228
rect 124948 89188 124988 89228
rect 125030 89188 125070 89228
rect 125112 89188 125152 89228
rect 139904 89188 139944 89228
rect 139986 89188 140026 89228
rect 140068 89188 140108 89228
rect 140150 89188 140190 89228
rect 140232 89188 140272 89228
rect 78184 88432 78224 88472
rect 78266 88432 78306 88472
rect 78348 88432 78388 88472
rect 78430 88432 78470 88472
rect 78512 88432 78552 88472
rect 93304 88432 93344 88472
rect 93386 88432 93426 88472
rect 93468 88432 93508 88472
rect 93550 88432 93590 88472
rect 93632 88432 93672 88472
rect 108424 88432 108464 88472
rect 108506 88432 108546 88472
rect 108588 88432 108628 88472
rect 108670 88432 108710 88472
rect 108752 88432 108792 88472
rect 123544 88432 123584 88472
rect 123626 88432 123666 88472
rect 123708 88432 123748 88472
rect 123790 88432 123830 88472
rect 123872 88432 123912 88472
rect 138664 88432 138704 88472
rect 138746 88432 138786 88472
rect 138828 88432 138868 88472
rect 138910 88432 138950 88472
rect 138992 88432 139032 88472
rect 148204 87844 148244 87884
rect 79424 87676 79464 87716
rect 79506 87676 79546 87716
rect 79588 87676 79628 87716
rect 79670 87676 79710 87716
rect 79752 87676 79792 87716
rect 94544 87676 94584 87716
rect 94626 87676 94666 87716
rect 94708 87676 94748 87716
rect 94790 87676 94830 87716
rect 94872 87676 94912 87716
rect 109664 87676 109704 87716
rect 109746 87676 109786 87716
rect 109828 87676 109868 87716
rect 109910 87676 109950 87716
rect 109992 87676 110032 87716
rect 124784 87676 124824 87716
rect 124866 87676 124906 87716
rect 124948 87676 124988 87716
rect 125030 87676 125070 87716
rect 125112 87676 125152 87716
rect 139904 87676 139944 87716
rect 139986 87676 140026 87716
rect 140068 87676 140108 87716
rect 140150 87676 140190 87716
rect 140232 87676 140272 87716
rect 78184 86920 78224 86960
rect 78266 86920 78306 86960
rect 78348 86920 78388 86960
rect 78430 86920 78470 86960
rect 78512 86920 78552 86960
rect 93304 86920 93344 86960
rect 93386 86920 93426 86960
rect 93468 86920 93508 86960
rect 93550 86920 93590 86960
rect 93632 86920 93672 86960
rect 108424 86920 108464 86960
rect 108506 86920 108546 86960
rect 108588 86920 108628 86960
rect 108670 86920 108710 86960
rect 108752 86920 108792 86960
rect 123544 86920 123584 86960
rect 123626 86920 123666 86960
rect 123708 86920 123748 86960
rect 123790 86920 123830 86960
rect 123872 86920 123912 86960
rect 138664 86920 138704 86960
rect 138746 86920 138786 86960
rect 138828 86920 138868 86960
rect 138910 86920 138950 86960
rect 138992 86920 139032 86960
rect 79424 86164 79464 86204
rect 79506 86164 79546 86204
rect 79588 86164 79628 86204
rect 79670 86164 79710 86204
rect 79752 86164 79792 86204
rect 94544 86164 94584 86204
rect 94626 86164 94666 86204
rect 94708 86164 94748 86204
rect 94790 86164 94830 86204
rect 94872 86164 94912 86204
rect 109664 86164 109704 86204
rect 109746 86164 109786 86204
rect 109828 86164 109868 86204
rect 109910 86164 109950 86204
rect 109992 86164 110032 86204
rect 124784 86164 124824 86204
rect 124866 86164 124906 86204
rect 124948 86164 124988 86204
rect 125030 86164 125070 86204
rect 125112 86164 125152 86204
rect 139904 86164 139944 86204
rect 139986 86164 140026 86204
rect 140068 86164 140108 86204
rect 140150 86164 140190 86204
rect 140232 86164 140272 86204
rect 78184 85408 78224 85448
rect 78266 85408 78306 85448
rect 78348 85408 78388 85448
rect 78430 85408 78470 85448
rect 78512 85408 78552 85448
rect 93304 85408 93344 85448
rect 93386 85408 93426 85448
rect 93468 85408 93508 85448
rect 93550 85408 93590 85448
rect 93632 85408 93672 85448
rect 108424 85408 108464 85448
rect 108506 85408 108546 85448
rect 108588 85408 108628 85448
rect 108670 85408 108710 85448
rect 108752 85408 108792 85448
rect 123544 85408 123584 85448
rect 123626 85408 123666 85448
rect 123708 85408 123748 85448
rect 123790 85408 123830 85448
rect 123872 85408 123912 85448
rect 138664 85408 138704 85448
rect 138746 85408 138786 85448
rect 138828 85408 138868 85448
rect 138910 85408 138950 85448
rect 138992 85408 139032 85448
rect 79424 84652 79464 84692
rect 79506 84652 79546 84692
rect 79588 84652 79628 84692
rect 79670 84652 79710 84692
rect 79752 84652 79792 84692
rect 94544 84652 94584 84692
rect 94626 84652 94666 84692
rect 94708 84652 94748 84692
rect 94790 84652 94830 84692
rect 94872 84652 94912 84692
rect 109664 84652 109704 84692
rect 109746 84652 109786 84692
rect 109828 84652 109868 84692
rect 109910 84652 109950 84692
rect 109992 84652 110032 84692
rect 124784 84652 124824 84692
rect 124866 84652 124906 84692
rect 124948 84652 124988 84692
rect 125030 84652 125070 84692
rect 125112 84652 125152 84692
rect 139904 84652 139944 84692
rect 139986 84652 140026 84692
rect 140068 84652 140108 84692
rect 140150 84652 140190 84692
rect 140232 84652 140272 84692
rect 78184 83896 78224 83936
rect 78266 83896 78306 83936
rect 78348 83896 78388 83936
rect 78430 83896 78470 83936
rect 78512 83896 78552 83936
rect 93304 83896 93344 83936
rect 93386 83896 93426 83936
rect 93468 83896 93508 83936
rect 93550 83896 93590 83936
rect 93632 83896 93672 83936
rect 108424 83896 108464 83936
rect 108506 83896 108546 83936
rect 108588 83896 108628 83936
rect 108670 83896 108710 83936
rect 108752 83896 108792 83936
rect 123544 83896 123584 83936
rect 123626 83896 123666 83936
rect 123708 83896 123748 83936
rect 123790 83896 123830 83936
rect 123872 83896 123912 83936
rect 138664 83896 138704 83936
rect 138746 83896 138786 83936
rect 138828 83896 138868 83936
rect 138910 83896 138950 83936
rect 138992 83896 139032 83936
rect 79424 83140 79464 83180
rect 79506 83140 79546 83180
rect 79588 83140 79628 83180
rect 79670 83140 79710 83180
rect 79752 83140 79792 83180
rect 94544 83140 94584 83180
rect 94626 83140 94666 83180
rect 94708 83140 94748 83180
rect 94790 83140 94830 83180
rect 94872 83140 94912 83180
rect 109664 83140 109704 83180
rect 109746 83140 109786 83180
rect 109828 83140 109868 83180
rect 109910 83140 109950 83180
rect 109992 83140 110032 83180
rect 124784 83140 124824 83180
rect 124866 83140 124906 83180
rect 124948 83140 124988 83180
rect 125030 83140 125070 83180
rect 125112 83140 125152 83180
rect 139904 83140 139944 83180
rect 139986 83140 140026 83180
rect 140068 83140 140108 83180
rect 140150 83140 140190 83180
rect 140232 83140 140272 83180
rect 78184 82384 78224 82424
rect 78266 82384 78306 82424
rect 78348 82384 78388 82424
rect 78430 82384 78470 82424
rect 78512 82384 78552 82424
rect 93304 82384 93344 82424
rect 93386 82384 93426 82424
rect 93468 82384 93508 82424
rect 93550 82384 93590 82424
rect 93632 82384 93672 82424
rect 108424 82384 108464 82424
rect 108506 82384 108546 82424
rect 108588 82384 108628 82424
rect 108670 82384 108710 82424
rect 108752 82384 108792 82424
rect 123544 82384 123584 82424
rect 123626 82384 123666 82424
rect 123708 82384 123748 82424
rect 123790 82384 123830 82424
rect 123872 82384 123912 82424
rect 138664 82384 138704 82424
rect 138746 82384 138786 82424
rect 138828 82384 138868 82424
rect 138910 82384 138950 82424
rect 138992 82384 139032 82424
rect 79424 81628 79464 81668
rect 79506 81628 79546 81668
rect 79588 81628 79628 81668
rect 79670 81628 79710 81668
rect 79752 81628 79792 81668
rect 94544 81628 94584 81668
rect 94626 81628 94666 81668
rect 94708 81628 94748 81668
rect 94790 81628 94830 81668
rect 94872 81628 94912 81668
rect 109664 81628 109704 81668
rect 109746 81628 109786 81668
rect 109828 81628 109868 81668
rect 109910 81628 109950 81668
rect 109992 81628 110032 81668
rect 124784 81628 124824 81668
rect 124866 81628 124906 81668
rect 124948 81628 124988 81668
rect 125030 81628 125070 81668
rect 125112 81628 125152 81668
rect 139904 81628 139944 81668
rect 139986 81628 140026 81668
rect 140068 81628 140108 81668
rect 140150 81628 140190 81668
rect 140232 81628 140272 81668
rect 78184 80872 78224 80912
rect 78266 80872 78306 80912
rect 78348 80872 78388 80912
rect 78430 80872 78470 80912
rect 78512 80872 78552 80912
rect 93304 80872 93344 80912
rect 93386 80872 93426 80912
rect 93468 80872 93508 80912
rect 93550 80872 93590 80912
rect 93632 80872 93672 80912
rect 108424 80872 108464 80912
rect 108506 80872 108546 80912
rect 108588 80872 108628 80912
rect 108670 80872 108710 80912
rect 108752 80872 108792 80912
rect 123544 80872 123584 80912
rect 123626 80872 123666 80912
rect 123708 80872 123748 80912
rect 123790 80872 123830 80912
rect 123872 80872 123912 80912
rect 138664 80872 138704 80912
rect 138746 80872 138786 80912
rect 138828 80872 138868 80912
rect 138910 80872 138950 80912
rect 138992 80872 139032 80912
rect 79424 80116 79464 80156
rect 79506 80116 79546 80156
rect 79588 80116 79628 80156
rect 79670 80116 79710 80156
rect 79752 80116 79792 80156
rect 94544 80116 94584 80156
rect 94626 80116 94666 80156
rect 94708 80116 94748 80156
rect 94790 80116 94830 80156
rect 94872 80116 94912 80156
rect 109664 80116 109704 80156
rect 109746 80116 109786 80156
rect 109828 80116 109868 80156
rect 109910 80116 109950 80156
rect 109992 80116 110032 80156
rect 124784 80116 124824 80156
rect 124866 80116 124906 80156
rect 124948 80116 124988 80156
rect 125030 80116 125070 80156
rect 125112 80116 125152 80156
rect 139904 80116 139944 80156
rect 139986 80116 140026 80156
rect 140068 80116 140108 80156
rect 140150 80116 140190 80156
rect 140232 80116 140272 80156
rect 78184 79360 78224 79400
rect 78266 79360 78306 79400
rect 78348 79360 78388 79400
rect 78430 79360 78470 79400
rect 78512 79360 78552 79400
rect 93304 79360 93344 79400
rect 93386 79360 93426 79400
rect 93468 79360 93508 79400
rect 93550 79360 93590 79400
rect 93632 79360 93672 79400
rect 108424 79360 108464 79400
rect 108506 79360 108546 79400
rect 108588 79360 108628 79400
rect 108670 79360 108710 79400
rect 108752 79360 108792 79400
rect 123544 79360 123584 79400
rect 123626 79360 123666 79400
rect 123708 79360 123748 79400
rect 123790 79360 123830 79400
rect 123872 79360 123912 79400
rect 138664 79360 138704 79400
rect 138746 79360 138786 79400
rect 138828 79360 138868 79400
rect 138910 79360 138950 79400
rect 138992 79360 139032 79400
rect 79424 78604 79464 78644
rect 79506 78604 79546 78644
rect 79588 78604 79628 78644
rect 79670 78604 79710 78644
rect 79752 78604 79792 78644
rect 94544 78604 94584 78644
rect 94626 78604 94666 78644
rect 94708 78604 94748 78644
rect 94790 78604 94830 78644
rect 94872 78604 94912 78644
rect 109664 78604 109704 78644
rect 109746 78604 109786 78644
rect 109828 78604 109868 78644
rect 109910 78604 109950 78644
rect 109992 78604 110032 78644
rect 124784 78604 124824 78644
rect 124866 78604 124906 78644
rect 124948 78604 124988 78644
rect 125030 78604 125070 78644
rect 125112 78604 125152 78644
rect 139904 78604 139944 78644
rect 139986 78604 140026 78644
rect 140068 78604 140108 78644
rect 140150 78604 140190 78644
rect 140232 78604 140272 78644
rect 78184 77848 78224 77888
rect 78266 77848 78306 77888
rect 78348 77848 78388 77888
rect 78430 77848 78470 77888
rect 78512 77848 78552 77888
rect 93304 77848 93344 77888
rect 93386 77848 93426 77888
rect 93468 77848 93508 77888
rect 93550 77848 93590 77888
rect 93632 77848 93672 77888
rect 108424 77848 108464 77888
rect 108506 77848 108546 77888
rect 108588 77848 108628 77888
rect 108670 77848 108710 77888
rect 108752 77848 108792 77888
rect 123544 77848 123584 77888
rect 123626 77848 123666 77888
rect 123708 77848 123748 77888
rect 123790 77848 123830 77888
rect 123872 77848 123912 77888
rect 138664 77848 138704 77888
rect 138746 77848 138786 77888
rect 138828 77848 138868 77888
rect 138910 77848 138950 77888
rect 138992 77848 139032 77888
rect 79424 77092 79464 77132
rect 79506 77092 79546 77132
rect 79588 77092 79628 77132
rect 79670 77092 79710 77132
rect 79752 77092 79792 77132
rect 94544 77092 94584 77132
rect 94626 77092 94666 77132
rect 94708 77092 94748 77132
rect 94790 77092 94830 77132
rect 94872 77092 94912 77132
rect 109664 77092 109704 77132
rect 109746 77092 109786 77132
rect 109828 77092 109868 77132
rect 109910 77092 109950 77132
rect 109992 77092 110032 77132
rect 124784 77092 124824 77132
rect 124866 77092 124906 77132
rect 124948 77092 124988 77132
rect 125030 77092 125070 77132
rect 125112 77092 125152 77132
rect 139904 77092 139944 77132
rect 139986 77092 140026 77132
rect 140068 77092 140108 77132
rect 140150 77092 140190 77132
rect 140232 77092 140272 77132
rect 78184 76336 78224 76376
rect 78266 76336 78306 76376
rect 78348 76336 78388 76376
rect 78430 76336 78470 76376
rect 78512 76336 78552 76376
rect 93304 76336 93344 76376
rect 93386 76336 93426 76376
rect 93468 76336 93508 76376
rect 93550 76336 93590 76376
rect 93632 76336 93672 76376
rect 108424 76336 108464 76376
rect 108506 76336 108546 76376
rect 108588 76336 108628 76376
rect 108670 76336 108710 76376
rect 108752 76336 108792 76376
rect 123544 76336 123584 76376
rect 123626 76336 123666 76376
rect 123708 76336 123748 76376
rect 123790 76336 123830 76376
rect 123872 76336 123912 76376
rect 138664 76336 138704 76376
rect 138746 76336 138786 76376
rect 138828 76336 138868 76376
rect 138910 76336 138950 76376
rect 138992 76336 139032 76376
rect 148204 75748 148244 75788
rect 79424 75580 79464 75620
rect 79506 75580 79546 75620
rect 79588 75580 79628 75620
rect 79670 75580 79710 75620
rect 79752 75580 79792 75620
rect 94544 75580 94584 75620
rect 94626 75580 94666 75620
rect 94708 75580 94748 75620
rect 94790 75580 94830 75620
rect 94872 75580 94912 75620
rect 109664 75580 109704 75620
rect 109746 75580 109786 75620
rect 109828 75580 109868 75620
rect 109910 75580 109950 75620
rect 109992 75580 110032 75620
rect 124784 75580 124824 75620
rect 124866 75580 124906 75620
rect 124948 75580 124988 75620
rect 125030 75580 125070 75620
rect 125112 75580 125152 75620
rect 139904 75580 139944 75620
rect 139986 75580 140026 75620
rect 140068 75580 140108 75620
rect 140150 75580 140190 75620
rect 140232 75580 140272 75620
<< metal2 >>
rect 103660 158420 103700 160020
rect 112299 159704 112341 159713
rect 112299 159664 112300 159704
rect 112340 159664 112341 159704
rect 112299 159655 112341 159664
rect 103660 158380 103988 158420
rect 64107 152060 64149 152069
rect 64107 152020 64108 152060
rect 64148 152020 64149 152060
rect 64107 152018 64149 152020
rect 63984 152011 64149 152018
rect 94059 152060 94101 152069
rect 94059 152020 94060 152060
rect 94100 152020 94101 152060
rect 94059 152011 94101 152020
rect 63984 151978 64148 152011
rect 79424 148196 79792 148205
rect 79464 148156 79506 148196
rect 79546 148156 79588 148196
rect 79628 148156 79670 148196
rect 79710 148156 79752 148196
rect 79424 148147 79792 148156
rect 78184 147440 78552 147449
rect 78224 147400 78266 147440
rect 78306 147400 78348 147440
rect 78388 147400 78430 147440
rect 78470 147400 78512 147440
rect 78184 147391 78552 147400
rect 93304 147440 93672 147449
rect 93344 147400 93386 147440
rect 93426 147400 93468 147440
rect 93508 147400 93550 147440
rect 93590 147400 93632 147440
rect 93304 147391 93672 147400
rect 79424 146684 79792 146693
rect 79464 146644 79506 146684
rect 79546 146644 79588 146684
rect 79628 146644 79670 146684
rect 79710 146644 79752 146684
rect 79424 146635 79792 146644
rect 78184 145928 78552 145937
rect 78224 145888 78266 145928
rect 78306 145888 78348 145928
rect 78388 145888 78430 145928
rect 78470 145888 78512 145928
rect 78184 145879 78552 145888
rect 93304 145928 93672 145937
rect 93344 145888 93386 145928
rect 93426 145888 93468 145928
rect 93508 145888 93550 145928
rect 93590 145888 93632 145928
rect 93304 145879 93672 145888
rect 79424 145172 79792 145181
rect 79464 145132 79506 145172
rect 79546 145132 79588 145172
rect 79628 145132 79670 145172
rect 79710 145132 79752 145172
rect 79424 145123 79792 145132
rect 78184 144416 78552 144425
rect 78224 144376 78266 144416
rect 78306 144376 78348 144416
rect 78388 144376 78430 144416
rect 78470 144376 78512 144416
rect 78184 144367 78552 144376
rect 93304 144416 93672 144425
rect 93344 144376 93386 144416
rect 93426 144376 93468 144416
rect 93508 144376 93550 144416
rect 93590 144376 93632 144416
rect 93304 144367 93672 144376
rect 79424 143660 79792 143669
rect 79464 143620 79506 143660
rect 79546 143620 79588 143660
rect 79628 143620 79670 143660
rect 79710 143620 79752 143660
rect 79424 143611 79792 143620
rect 78184 142904 78552 142913
rect 78224 142864 78266 142904
rect 78306 142864 78348 142904
rect 78388 142864 78430 142904
rect 78470 142864 78512 142904
rect 78184 142855 78552 142864
rect 93304 142904 93672 142913
rect 93344 142864 93386 142904
rect 93426 142864 93468 142904
rect 93508 142864 93550 142904
rect 93590 142864 93632 142904
rect 93304 142855 93672 142864
rect 79424 142148 79792 142157
rect 79464 142108 79506 142148
rect 79546 142108 79588 142148
rect 79628 142108 79670 142148
rect 79710 142108 79752 142148
rect 79424 142099 79792 142108
rect 78184 141392 78552 141401
rect 78224 141352 78266 141392
rect 78306 141352 78348 141392
rect 78388 141352 78430 141392
rect 78470 141352 78512 141392
rect 78184 141343 78552 141352
rect 93304 141392 93672 141401
rect 93344 141352 93386 141392
rect 93426 141352 93468 141392
rect 93508 141352 93550 141392
rect 93590 141352 93632 141392
rect 93304 141343 93672 141352
rect 79424 140636 79792 140645
rect 79464 140596 79506 140636
rect 79546 140596 79588 140636
rect 79628 140596 79670 140636
rect 79710 140596 79752 140636
rect 79424 140587 79792 140596
rect 78184 139880 78552 139889
rect 78224 139840 78266 139880
rect 78306 139840 78348 139880
rect 78388 139840 78430 139880
rect 78470 139840 78512 139880
rect 78184 139831 78552 139840
rect 93304 139880 93672 139889
rect 93344 139840 93386 139880
rect 93426 139840 93468 139880
rect 93508 139840 93550 139880
rect 93590 139840 93632 139880
rect 93304 139831 93672 139840
rect 79424 139124 79792 139133
rect 79464 139084 79506 139124
rect 79546 139084 79588 139124
rect 79628 139084 79670 139124
rect 79710 139084 79752 139124
rect 79424 139075 79792 139084
rect 78184 138368 78552 138377
rect 78224 138328 78266 138368
rect 78306 138328 78348 138368
rect 78388 138328 78430 138368
rect 78470 138328 78512 138368
rect 78184 138319 78552 138328
rect 93304 138368 93672 138377
rect 93344 138328 93386 138368
rect 93426 138328 93468 138368
rect 93508 138328 93550 138368
rect 93590 138328 93632 138368
rect 93304 138319 93672 138328
rect 79424 137612 79792 137621
rect 79464 137572 79506 137612
rect 79546 137572 79588 137612
rect 79628 137572 79670 137612
rect 79710 137572 79752 137612
rect 79424 137563 79792 137572
rect 78184 136856 78552 136865
rect 78224 136816 78266 136856
rect 78306 136816 78348 136856
rect 78388 136816 78430 136856
rect 78470 136816 78512 136856
rect 78184 136807 78552 136816
rect 93304 136856 93672 136865
rect 93344 136816 93386 136856
rect 93426 136816 93468 136856
rect 93508 136816 93550 136856
rect 93590 136816 93632 136856
rect 93304 136807 93672 136816
rect 79424 136100 79792 136109
rect 79464 136060 79506 136100
rect 79546 136060 79588 136100
rect 79628 136060 79670 136100
rect 79710 136060 79752 136100
rect 79424 136051 79792 136060
rect 63984 135976 64148 136016
rect 64108 135437 64148 135976
rect 78603 135512 78645 135521
rect 78603 135472 78604 135512
rect 78644 135472 78645 135512
rect 78603 135463 78645 135472
rect 64107 135428 64149 135437
rect 64107 135388 64108 135428
rect 64148 135388 64149 135428
rect 64107 135379 64149 135388
rect 78184 135344 78552 135353
rect 78224 135304 78266 135344
rect 78306 135304 78348 135344
rect 78388 135304 78430 135344
rect 78470 135304 78512 135344
rect 78184 135295 78552 135304
rect 78184 133832 78552 133841
rect 78224 133792 78266 133832
rect 78306 133792 78348 133832
rect 78388 133792 78430 133832
rect 78470 133792 78512 133832
rect 78184 133783 78552 133792
rect 78604 132740 78644 135463
rect 93304 135344 93672 135353
rect 93344 135304 93386 135344
rect 93426 135304 93468 135344
rect 93508 135304 93550 135344
rect 93590 135304 93632 135344
rect 93304 135295 93672 135304
rect 79424 134588 79792 134597
rect 79464 134548 79506 134588
rect 79546 134548 79588 134588
rect 79628 134548 79670 134588
rect 79710 134548 79752 134588
rect 79424 134539 79792 134548
rect 93304 133832 93672 133841
rect 93344 133792 93386 133832
rect 93426 133792 93468 133832
rect 93508 133792 93550 133832
rect 93590 133792 93632 133832
rect 93304 133783 93672 133792
rect 79424 133076 79792 133085
rect 79464 133036 79506 133076
rect 79546 133036 79588 133076
rect 79628 133036 79670 133076
rect 79710 133036 79752 133076
rect 79424 133027 79792 133036
rect 78604 132691 78644 132700
rect 79275 132572 79317 132581
rect 79275 132532 79276 132572
rect 79316 132532 79317 132572
rect 79275 132523 79317 132532
rect 79276 132438 79316 132523
rect 78184 132320 78552 132329
rect 78224 132280 78266 132320
rect 78306 132280 78348 132320
rect 78388 132280 78430 132320
rect 78470 132280 78512 132320
rect 78184 132271 78552 132280
rect 93304 132320 93672 132329
rect 93344 132280 93386 132320
rect 93426 132280 93468 132320
rect 93508 132280 93550 132320
rect 93590 132280 93632 132320
rect 93304 132271 93672 132280
rect 79424 131564 79792 131573
rect 79464 131524 79506 131564
rect 79546 131524 79588 131564
rect 79628 131524 79670 131564
rect 79710 131524 79752 131564
rect 79424 131515 79792 131524
rect 78184 130808 78552 130817
rect 78224 130768 78266 130808
rect 78306 130768 78348 130808
rect 78388 130768 78430 130808
rect 78470 130768 78512 130808
rect 78184 130759 78552 130768
rect 93304 130808 93672 130817
rect 93344 130768 93386 130808
rect 93426 130768 93468 130808
rect 93508 130768 93550 130808
rect 93590 130768 93632 130808
rect 93304 130759 93672 130768
rect 79424 130052 79792 130061
rect 79464 130012 79506 130052
rect 79546 130012 79588 130052
rect 79628 130012 79670 130052
rect 79710 130012 79752 130052
rect 79424 130003 79792 130012
rect 73323 129716 73365 129725
rect 73323 129676 73324 129716
rect 73364 129676 73365 129716
rect 73323 129667 73365 129676
rect 64107 120896 64149 120905
rect 64107 120856 64108 120896
rect 64148 120856 64149 120896
rect 64107 120847 64149 120856
rect 64108 120014 64148 120847
rect 63984 119974 64148 120014
rect 64107 105020 64149 105029
rect 64107 104980 64108 105020
rect 64148 104980 64149 105020
rect 64107 104971 64149 104980
rect 64108 104012 64148 104971
rect 63984 103972 64148 104012
rect 64107 88010 64149 88019
rect 63984 87970 64108 88010
rect 64148 87970 64149 88010
rect 64107 87961 64149 87970
rect 64107 72008 64149 72017
rect 63984 71968 64108 72008
rect 64148 71968 64149 72008
rect 64107 71959 64149 71968
rect 73324 64205 73364 129667
rect 78184 129296 78552 129305
rect 78224 129256 78266 129296
rect 78306 129256 78348 129296
rect 78388 129256 78430 129296
rect 78470 129256 78512 129296
rect 78184 129247 78552 129256
rect 93304 129296 93672 129305
rect 93344 129256 93386 129296
rect 93426 129256 93468 129296
rect 93508 129256 93550 129296
rect 93590 129256 93632 129296
rect 93304 129247 93672 129256
rect 93868 128876 93908 128885
rect 79424 128540 79792 128549
rect 79464 128500 79506 128540
rect 79546 128500 79588 128540
rect 79628 128500 79670 128540
rect 79710 128500 79752 128540
rect 79424 128491 79792 128500
rect 78184 127784 78552 127793
rect 78224 127744 78266 127784
rect 78306 127744 78348 127784
rect 78388 127744 78430 127784
rect 78470 127744 78512 127784
rect 78184 127735 78552 127744
rect 93304 127784 93672 127793
rect 93344 127744 93386 127784
rect 93426 127744 93468 127784
rect 93508 127744 93550 127784
rect 93590 127744 93632 127784
rect 93304 127735 93672 127744
rect 79851 127280 79893 127289
rect 79851 127240 79852 127280
rect 79892 127240 79893 127280
rect 79851 127231 79893 127240
rect 79424 127028 79792 127037
rect 79464 126988 79506 127028
rect 79546 126988 79588 127028
rect 79628 126988 79670 127028
rect 79710 126988 79752 127028
rect 79424 126979 79792 126988
rect 78184 126272 78552 126281
rect 78224 126232 78266 126272
rect 78306 126232 78348 126272
rect 78388 126232 78430 126272
rect 78470 126232 78512 126272
rect 78184 126223 78552 126232
rect 79424 125516 79792 125525
rect 79464 125476 79506 125516
rect 79546 125476 79588 125516
rect 79628 125476 79670 125516
rect 79710 125476 79752 125516
rect 79424 125467 79792 125476
rect 78184 124760 78552 124769
rect 78224 124720 78266 124760
rect 78306 124720 78348 124760
rect 78388 124720 78430 124760
rect 78470 124720 78512 124760
rect 78184 124711 78552 124720
rect 79564 124592 79604 124601
rect 79852 124592 79892 127231
rect 93771 126608 93813 126617
rect 93771 126568 93772 126608
rect 93812 126568 93813 126608
rect 93771 126559 93813 126568
rect 93304 126272 93672 126281
rect 93344 126232 93386 126272
rect 93426 126232 93468 126272
rect 93508 126232 93550 126272
rect 93590 126232 93632 126272
rect 93304 126223 93672 126232
rect 93772 125273 93812 126559
rect 93771 125264 93813 125273
rect 93771 125224 93772 125264
rect 93812 125224 93813 125264
rect 93771 125215 93813 125224
rect 93304 124760 93672 124769
rect 93344 124720 93386 124760
rect 93426 124720 93468 124760
rect 93508 124720 93550 124760
rect 93590 124720 93632 124760
rect 93304 124711 93672 124720
rect 79604 124552 79892 124592
rect 79564 124543 79604 124552
rect 93868 124349 93908 128836
rect 93964 128876 94004 128885
rect 93964 126785 94004 128836
rect 94060 128792 94100 152011
rect 94544 148196 94912 148205
rect 94584 148156 94626 148196
rect 94666 148156 94708 148196
rect 94748 148156 94790 148196
rect 94830 148156 94872 148196
rect 94544 148147 94912 148156
rect 94544 146684 94912 146693
rect 94584 146644 94626 146684
rect 94666 146644 94708 146684
rect 94748 146644 94790 146684
rect 94830 146644 94872 146684
rect 94544 146635 94912 146644
rect 94544 145172 94912 145181
rect 94584 145132 94626 145172
rect 94666 145132 94708 145172
rect 94748 145132 94790 145172
rect 94830 145132 94872 145172
rect 94544 145123 94912 145132
rect 94544 143660 94912 143669
rect 94584 143620 94626 143660
rect 94666 143620 94708 143660
rect 94748 143620 94790 143660
rect 94830 143620 94872 143660
rect 94544 143611 94912 143620
rect 94544 142148 94912 142157
rect 94584 142108 94626 142148
rect 94666 142108 94708 142148
rect 94748 142108 94790 142148
rect 94830 142108 94872 142148
rect 94544 142099 94912 142108
rect 94544 140636 94912 140645
rect 94584 140596 94626 140636
rect 94666 140596 94708 140636
rect 94748 140596 94790 140636
rect 94830 140596 94872 140636
rect 94544 140587 94912 140596
rect 94544 139124 94912 139133
rect 94584 139084 94626 139124
rect 94666 139084 94708 139124
rect 94748 139084 94790 139124
rect 94830 139084 94872 139124
rect 94544 139075 94912 139084
rect 94544 137612 94912 137621
rect 94584 137572 94626 137612
rect 94666 137572 94708 137612
rect 94748 137572 94790 137612
rect 94830 137572 94872 137612
rect 94544 137563 94912 137572
rect 94544 136100 94912 136109
rect 94584 136060 94626 136100
rect 94666 136060 94708 136100
rect 94748 136060 94790 136100
rect 94830 136060 94872 136100
rect 94544 136051 94912 136060
rect 94544 134588 94912 134597
rect 94584 134548 94626 134588
rect 94666 134548 94708 134588
rect 94748 134548 94790 134588
rect 94830 134548 94872 134588
rect 94544 134539 94912 134548
rect 97419 134252 97461 134261
rect 97419 134212 97420 134252
rect 97460 134212 97461 134252
rect 97419 134203 97461 134212
rect 97804 134252 97844 134261
rect 97420 134118 97460 134203
rect 97804 133580 97844 134212
rect 98187 134252 98229 134261
rect 98187 134212 98188 134252
rect 98228 134212 98229 134252
rect 98187 134203 98229 134212
rect 98667 134252 98709 134261
rect 98667 134212 98668 134252
rect 98708 134212 98709 134252
rect 98667 134203 98709 134212
rect 98188 133664 98228 134203
rect 98668 134118 98708 134203
rect 99819 134084 99861 134093
rect 99819 134044 99820 134084
rect 99860 134044 99861 134084
rect 99819 134035 99861 134044
rect 100011 134084 100053 134093
rect 100011 134044 100012 134084
rect 100052 134044 100053 134084
rect 100011 134035 100053 134044
rect 99820 133950 99860 134035
rect 98188 133615 98228 133624
rect 97804 133531 97844 133540
rect 98860 133412 98900 133421
rect 94544 133076 94912 133085
rect 94584 133036 94626 133076
rect 94666 133036 94708 133076
rect 94748 133036 94790 133076
rect 94830 133036 94872 133076
rect 94544 133027 94912 133036
rect 98668 132908 98708 132917
rect 98860 132908 98900 133372
rect 98708 132868 98900 132908
rect 98668 132859 98708 132868
rect 100012 132749 100052 134035
rect 98572 132740 98612 132749
rect 94251 132572 94293 132581
rect 94251 132532 94252 132572
rect 94292 132532 94293 132572
rect 94251 132523 94293 132532
rect 94155 129884 94197 129893
rect 94155 129844 94156 129884
rect 94196 129844 94197 129884
rect 94155 129835 94197 129844
rect 94156 129128 94196 129835
rect 94156 129079 94196 129088
rect 94060 126869 94100 128752
rect 94156 128708 94196 128717
rect 94252 128708 94292 132523
rect 98380 131900 98420 131909
rect 98092 131860 98380 131900
rect 94544 131564 94912 131573
rect 94584 131524 94626 131564
rect 94666 131524 94708 131564
rect 94748 131524 94790 131564
rect 94830 131524 94872 131564
rect 94544 131515 94912 131524
rect 98092 130640 98132 131860
rect 98380 131851 98420 131860
rect 98572 131816 98612 132700
rect 98763 132740 98805 132749
rect 98763 132700 98764 132740
rect 98804 132700 98805 132740
rect 98763 132691 98805 132700
rect 98860 132740 98900 132749
rect 98764 132606 98804 132691
rect 98860 132077 98900 132700
rect 100011 132740 100053 132749
rect 100011 132700 100012 132740
rect 100052 132700 100053 132740
rect 100011 132691 100053 132700
rect 102219 132740 102261 132749
rect 102219 132700 102220 132740
rect 102260 132700 102261 132740
rect 102219 132691 102261 132700
rect 102987 132740 103029 132749
rect 102987 132700 102988 132740
rect 103028 132700 103029 132740
rect 102987 132691 103029 132700
rect 103660 132740 103700 132749
rect 103852 132740 103892 132749
rect 103700 132700 103852 132740
rect 103660 132691 103700 132700
rect 103852 132691 103892 132700
rect 98859 132068 98901 132077
rect 98859 132028 98860 132068
rect 98900 132028 98901 132068
rect 98859 132019 98901 132028
rect 99051 132068 99093 132077
rect 99051 132028 99052 132068
rect 99092 132028 99093 132068
rect 99051 132019 99093 132028
rect 99435 132068 99477 132077
rect 99435 132028 99436 132068
rect 99476 132028 99477 132068
rect 99435 132019 99477 132028
rect 99052 131934 99092 132019
rect 99244 131900 99284 131909
rect 99148 131860 99244 131900
rect 99148 131816 99188 131860
rect 99244 131851 99284 131860
rect 99340 131900 99380 131909
rect 98572 131776 99188 131816
rect 99243 131732 99285 131741
rect 99243 131692 99244 131732
rect 99284 131692 99285 131732
rect 99243 131683 99285 131692
rect 98092 130591 98132 130600
rect 96843 130388 96885 130397
rect 96843 130348 96844 130388
rect 96884 130348 96885 130388
rect 98091 130388 98133 130397
rect 96843 130339 96885 130348
rect 97911 130377 97951 130386
rect 94544 130052 94912 130061
rect 94584 130012 94626 130052
rect 94666 130012 94708 130052
rect 94748 130012 94790 130052
rect 94830 130012 94872 130052
rect 94544 130003 94912 130012
rect 95019 129968 95061 129977
rect 95019 129928 95020 129968
rect 95060 129928 95061 129968
rect 95019 129919 95061 129928
rect 94196 128668 94484 128708
rect 94156 128659 94196 128668
rect 94444 127448 94484 128668
rect 94544 128540 94912 128549
rect 94584 128500 94626 128540
rect 94666 128500 94708 128540
rect 94748 128500 94790 128540
rect 94830 128500 94872 128540
rect 94544 128491 94912 128500
rect 94827 128372 94869 128381
rect 94827 128332 94828 128372
rect 94868 128332 94869 128372
rect 94827 128323 94869 128332
rect 94828 127616 94868 128323
rect 94828 127567 94868 127576
rect 95020 127448 95060 129919
rect 96171 129884 96213 129893
rect 96171 129844 96172 129884
rect 96212 129844 96213 129884
rect 96171 129835 96213 129844
rect 96844 129884 96884 130339
rect 98091 130348 98092 130388
rect 98132 130348 98133 130388
rect 98091 130339 98133 130348
rect 99051 130388 99093 130397
rect 99051 130348 99052 130388
rect 99092 130348 99093 130388
rect 99051 130339 99093 130348
rect 97227 130136 97269 130145
rect 97227 130096 97228 130136
rect 97268 130096 97269 130136
rect 97227 130087 97269 130096
rect 97131 129968 97173 129977
rect 97131 129928 97132 129968
rect 97172 129928 97173 129968
rect 97131 129919 97173 129928
rect 96844 129835 96884 129844
rect 96172 129716 96212 129835
rect 96172 129667 96212 129676
rect 97132 129716 97172 129919
rect 97228 129884 97268 130087
rect 97911 129968 97951 130337
rect 98092 130254 98132 130339
rect 97911 129928 98036 129968
rect 97228 129835 97268 129844
rect 97419 129884 97461 129893
rect 97419 129844 97420 129884
rect 97460 129844 97461 129884
rect 97419 129835 97461 129844
rect 97132 129667 97172 129676
rect 97324 129716 97364 129725
rect 97324 129212 97364 129676
rect 97420 129716 97460 129835
rect 97420 129667 97460 129676
rect 96748 129172 97364 129212
rect 96748 129128 96788 129172
rect 96748 129079 96788 129088
rect 96076 128876 96116 128885
rect 96076 128381 96116 128836
rect 96075 128372 96117 128381
rect 96075 128332 96076 128372
rect 96116 128332 96117 128372
rect 96075 128323 96117 128332
rect 97996 128297 98036 129928
rect 98955 129884 98997 129893
rect 98955 129844 98956 129884
rect 98996 129844 98997 129884
rect 98955 129835 98997 129844
rect 95499 128288 95541 128297
rect 95499 128248 95500 128288
rect 95540 128248 95541 128288
rect 95499 128239 95541 128248
rect 97995 128288 98037 128297
rect 97995 128248 97996 128288
rect 98036 128248 98037 128288
rect 97995 128239 98037 128248
rect 94444 127408 94639 127448
rect 94599 127364 94639 127408
rect 94732 127373 94772 127439
rect 95020 127408 95156 127448
rect 94599 127315 94639 127324
rect 94712 127364 94773 127373
rect 94772 127324 94773 127364
rect 94712 127315 94773 127324
rect 94828 127364 94868 127373
rect 94828 127196 94868 127324
rect 94924 127364 94964 127373
rect 94964 127324 95060 127364
rect 94924 127315 94964 127324
rect 94252 127156 94868 127196
rect 94059 126860 94101 126869
rect 94059 126820 94060 126860
rect 94100 126820 94101 126860
rect 94059 126811 94101 126820
rect 93963 126776 94005 126785
rect 93963 126736 93964 126776
rect 94004 126736 94005 126776
rect 93963 126727 94005 126736
rect 94252 126449 94292 127156
rect 94544 127028 94912 127037
rect 94584 126988 94626 127028
rect 94666 126988 94708 127028
rect 94748 126988 94790 127028
rect 94830 126988 94872 127028
rect 94544 126979 94912 126988
rect 94635 126860 94677 126869
rect 94635 126820 94636 126860
rect 94676 126820 94677 126860
rect 94635 126811 94677 126820
rect 94636 126726 94676 126811
rect 94731 126776 94773 126785
rect 94731 126736 94732 126776
rect 94772 126736 94773 126776
rect 94731 126727 94773 126736
rect 94251 126440 94293 126449
rect 94251 126400 94252 126440
rect 94292 126400 94293 126440
rect 94251 126391 94293 126400
rect 78891 124340 78933 124349
rect 78891 124300 78892 124340
rect 78932 124300 78933 124340
rect 78891 124291 78933 124300
rect 93867 124340 93909 124349
rect 93867 124300 93868 124340
rect 93908 124300 93909 124340
rect 93867 124291 93909 124300
rect 78184 123248 78552 123257
rect 78224 123208 78266 123248
rect 78306 123208 78348 123248
rect 78388 123208 78430 123248
rect 78470 123208 78512 123248
rect 78184 123199 78552 123208
rect 78184 121736 78552 121745
rect 78224 121696 78266 121736
rect 78306 121696 78348 121736
rect 78388 121696 78430 121736
rect 78470 121696 78512 121736
rect 78184 121687 78552 121696
rect 78892 120905 78932 124291
rect 79424 124004 79792 124013
rect 79464 123964 79506 124004
rect 79546 123964 79588 124004
rect 79628 123964 79670 124004
rect 79710 123964 79752 124004
rect 79424 123955 79792 123964
rect 93304 123248 93672 123257
rect 93344 123208 93386 123248
rect 93426 123208 93468 123248
rect 93508 123208 93550 123248
rect 93590 123208 93632 123248
rect 93304 123199 93672 123208
rect 79424 122492 79792 122501
rect 79464 122452 79506 122492
rect 79546 122452 79588 122492
rect 79628 122452 79670 122492
rect 79710 122452 79752 122492
rect 79424 122443 79792 122452
rect 93771 122408 93813 122417
rect 93771 122368 93772 122408
rect 93812 122368 93813 122408
rect 93771 122359 93813 122368
rect 93304 121736 93672 121745
rect 93344 121696 93386 121736
rect 93426 121696 93468 121736
rect 93508 121696 93550 121736
rect 93590 121696 93632 121736
rect 93304 121687 93672 121696
rect 79424 120980 79792 120989
rect 79464 120940 79506 120980
rect 79546 120940 79588 120980
rect 79628 120940 79670 120980
rect 79710 120940 79752 120980
rect 79424 120931 79792 120940
rect 78891 120896 78933 120905
rect 78891 120856 78892 120896
rect 78932 120856 78933 120896
rect 78891 120847 78933 120856
rect 78184 120224 78552 120233
rect 78224 120184 78266 120224
rect 78306 120184 78348 120224
rect 78388 120184 78430 120224
rect 78470 120184 78512 120224
rect 78184 120175 78552 120184
rect 93304 120224 93672 120233
rect 93344 120184 93386 120224
rect 93426 120184 93468 120224
rect 93508 120184 93550 120224
rect 93590 120184 93632 120224
rect 93304 120175 93672 120184
rect 79424 119468 79792 119477
rect 79464 119428 79506 119468
rect 79546 119428 79588 119468
rect 79628 119428 79670 119468
rect 79710 119428 79752 119468
rect 79424 119419 79792 119428
rect 78184 118712 78552 118721
rect 78224 118672 78266 118712
rect 78306 118672 78348 118712
rect 78388 118672 78430 118712
rect 78470 118672 78512 118712
rect 78184 118663 78552 118672
rect 93304 118712 93672 118721
rect 93344 118672 93386 118712
rect 93426 118672 93468 118712
rect 93508 118672 93550 118712
rect 93590 118672 93632 118712
rect 93304 118663 93672 118672
rect 79424 117956 79792 117965
rect 79464 117916 79506 117956
rect 79546 117916 79588 117956
rect 79628 117916 79670 117956
rect 79710 117916 79752 117956
rect 79424 117907 79792 117916
rect 78184 117200 78552 117209
rect 78224 117160 78266 117200
rect 78306 117160 78348 117200
rect 78388 117160 78430 117200
rect 78470 117160 78512 117200
rect 78184 117151 78552 117160
rect 93304 117200 93672 117209
rect 93344 117160 93386 117200
rect 93426 117160 93468 117200
rect 93508 117160 93550 117200
rect 93590 117160 93632 117200
rect 93304 117151 93672 117160
rect 79424 116444 79792 116453
rect 79464 116404 79506 116444
rect 79546 116404 79588 116444
rect 79628 116404 79670 116444
rect 79710 116404 79752 116444
rect 79424 116395 79792 116404
rect 78184 115688 78552 115697
rect 78224 115648 78266 115688
rect 78306 115648 78348 115688
rect 78388 115648 78430 115688
rect 78470 115648 78512 115688
rect 78184 115639 78552 115648
rect 93304 115688 93672 115697
rect 93344 115648 93386 115688
rect 93426 115648 93468 115688
rect 93508 115648 93550 115688
rect 93590 115648 93632 115688
rect 93304 115639 93672 115648
rect 79424 114932 79792 114941
rect 79464 114892 79506 114932
rect 79546 114892 79588 114932
rect 79628 114892 79670 114932
rect 79710 114892 79752 114932
rect 79424 114883 79792 114892
rect 78184 114176 78552 114185
rect 78224 114136 78266 114176
rect 78306 114136 78348 114176
rect 78388 114136 78430 114176
rect 78470 114136 78512 114176
rect 78184 114127 78552 114136
rect 93304 114176 93672 114185
rect 93344 114136 93386 114176
rect 93426 114136 93468 114176
rect 93508 114136 93550 114176
rect 93590 114136 93632 114176
rect 93304 114127 93672 114136
rect 79424 113420 79792 113429
rect 79464 113380 79506 113420
rect 79546 113380 79588 113420
rect 79628 113380 79670 113420
rect 79710 113380 79752 113420
rect 79424 113371 79792 113380
rect 78184 112664 78552 112673
rect 78224 112624 78266 112664
rect 78306 112624 78348 112664
rect 78388 112624 78430 112664
rect 78470 112624 78512 112664
rect 78184 112615 78552 112624
rect 93304 112664 93672 112673
rect 93344 112624 93386 112664
rect 93426 112624 93468 112664
rect 93508 112624 93550 112664
rect 93590 112624 93632 112664
rect 93304 112615 93672 112624
rect 79424 111908 79792 111917
rect 79464 111868 79506 111908
rect 79546 111868 79588 111908
rect 79628 111868 79670 111908
rect 79710 111868 79752 111908
rect 79424 111859 79792 111868
rect 78184 111152 78552 111161
rect 78224 111112 78266 111152
rect 78306 111112 78348 111152
rect 78388 111112 78430 111152
rect 78470 111112 78512 111152
rect 78184 111103 78552 111112
rect 93304 111152 93672 111161
rect 93344 111112 93386 111152
rect 93426 111112 93468 111152
rect 93508 111112 93550 111152
rect 93590 111112 93632 111152
rect 93304 111103 93672 111112
rect 79424 110396 79792 110405
rect 79464 110356 79506 110396
rect 79546 110356 79588 110396
rect 79628 110356 79670 110396
rect 79710 110356 79752 110396
rect 79424 110347 79792 110356
rect 78184 109640 78552 109649
rect 78224 109600 78266 109640
rect 78306 109600 78348 109640
rect 78388 109600 78430 109640
rect 78470 109600 78512 109640
rect 78184 109591 78552 109600
rect 93304 109640 93672 109649
rect 93344 109600 93386 109640
rect 93426 109600 93468 109640
rect 93508 109600 93550 109640
rect 93590 109600 93632 109640
rect 93304 109591 93672 109600
rect 79424 108884 79792 108893
rect 79464 108844 79506 108884
rect 79546 108844 79588 108884
rect 79628 108844 79670 108884
rect 79710 108844 79752 108884
rect 79424 108835 79792 108844
rect 78184 108128 78552 108137
rect 78224 108088 78266 108128
rect 78306 108088 78348 108128
rect 78388 108088 78430 108128
rect 78470 108088 78512 108128
rect 78184 108079 78552 108088
rect 93304 108128 93672 108137
rect 93344 108088 93386 108128
rect 93426 108088 93468 108128
rect 93508 108088 93550 108128
rect 93590 108088 93632 108128
rect 93304 108079 93672 108088
rect 79424 107372 79792 107381
rect 79464 107332 79506 107372
rect 79546 107332 79588 107372
rect 79628 107332 79670 107372
rect 79710 107332 79752 107372
rect 79424 107323 79792 107332
rect 78184 106616 78552 106625
rect 78224 106576 78266 106616
rect 78306 106576 78348 106616
rect 78388 106576 78430 106616
rect 78470 106576 78512 106616
rect 78184 106567 78552 106576
rect 93304 106616 93672 106625
rect 93344 106576 93386 106616
rect 93426 106576 93468 106616
rect 93508 106576 93550 106616
rect 93590 106576 93632 106616
rect 93304 106567 93672 106576
rect 79424 105860 79792 105869
rect 79464 105820 79506 105860
rect 79546 105820 79588 105860
rect 79628 105820 79670 105860
rect 79710 105820 79752 105860
rect 79424 105811 79792 105820
rect 78184 105104 78552 105113
rect 78224 105064 78266 105104
rect 78306 105064 78348 105104
rect 78388 105064 78430 105104
rect 78470 105064 78512 105104
rect 78184 105055 78552 105064
rect 93304 105104 93672 105113
rect 93344 105064 93386 105104
rect 93426 105064 93468 105104
rect 93508 105064 93550 105104
rect 93590 105064 93632 105104
rect 93304 105055 93672 105064
rect 79424 104348 79792 104357
rect 79464 104308 79506 104348
rect 79546 104308 79588 104348
rect 79628 104308 79670 104348
rect 79710 104308 79752 104348
rect 79424 104299 79792 104308
rect 78184 103592 78552 103601
rect 78224 103552 78266 103592
rect 78306 103552 78348 103592
rect 78388 103552 78430 103592
rect 78470 103552 78512 103592
rect 78184 103543 78552 103552
rect 93304 103592 93672 103601
rect 93344 103552 93386 103592
rect 93426 103552 93468 103592
rect 93508 103552 93550 103592
rect 93590 103552 93632 103592
rect 93304 103543 93672 103552
rect 79424 102836 79792 102845
rect 79464 102796 79506 102836
rect 79546 102796 79588 102836
rect 79628 102796 79670 102836
rect 79710 102796 79752 102836
rect 79424 102787 79792 102796
rect 78184 102080 78552 102089
rect 78224 102040 78266 102080
rect 78306 102040 78348 102080
rect 78388 102040 78430 102080
rect 78470 102040 78512 102080
rect 78184 102031 78552 102040
rect 93304 102080 93672 102089
rect 93344 102040 93386 102080
rect 93426 102040 93468 102080
rect 93508 102040 93550 102080
rect 93590 102040 93632 102080
rect 93304 102031 93672 102040
rect 79424 101324 79792 101333
rect 79464 101284 79506 101324
rect 79546 101284 79588 101324
rect 79628 101284 79670 101324
rect 79710 101284 79752 101324
rect 79424 101275 79792 101284
rect 78184 100568 78552 100577
rect 78224 100528 78266 100568
rect 78306 100528 78348 100568
rect 78388 100528 78430 100568
rect 78470 100528 78512 100568
rect 78184 100519 78552 100528
rect 93304 100568 93672 100577
rect 93344 100528 93386 100568
rect 93426 100528 93468 100568
rect 93508 100528 93550 100568
rect 93590 100528 93632 100568
rect 93304 100519 93672 100528
rect 79424 99812 79792 99821
rect 79464 99772 79506 99812
rect 79546 99772 79588 99812
rect 79628 99772 79670 99812
rect 79710 99772 79752 99812
rect 79424 99763 79792 99772
rect 78184 99056 78552 99065
rect 78224 99016 78266 99056
rect 78306 99016 78348 99056
rect 78388 99016 78430 99056
rect 78470 99016 78512 99056
rect 78184 99007 78552 99016
rect 93304 99056 93672 99065
rect 93344 99016 93386 99056
rect 93426 99016 93468 99056
rect 93508 99016 93550 99056
rect 93590 99016 93632 99056
rect 93304 99007 93672 99016
rect 79424 98300 79792 98309
rect 79464 98260 79506 98300
rect 79546 98260 79588 98300
rect 79628 98260 79670 98300
rect 79710 98260 79752 98300
rect 79424 98251 79792 98260
rect 78184 97544 78552 97553
rect 78224 97504 78266 97544
rect 78306 97504 78348 97544
rect 78388 97504 78430 97544
rect 78470 97504 78512 97544
rect 78184 97495 78552 97504
rect 93304 97544 93672 97553
rect 93344 97504 93386 97544
rect 93426 97504 93468 97544
rect 93508 97504 93550 97544
rect 93590 97504 93632 97544
rect 93304 97495 93672 97504
rect 79424 96788 79792 96797
rect 79464 96748 79506 96788
rect 79546 96748 79588 96788
rect 79628 96748 79670 96788
rect 79710 96748 79752 96788
rect 79424 96739 79792 96748
rect 78184 96032 78552 96041
rect 78224 95992 78266 96032
rect 78306 95992 78348 96032
rect 78388 95992 78430 96032
rect 78470 95992 78512 96032
rect 78184 95983 78552 95992
rect 93304 96032 93672 96041
rect 93344 95992 93386 96032
rect 93426 95992 93468 96032
rect 93508 95992 93550 96032
rect 93590 95992 93632 96032
rect 93304 95983 93672 95992
rect 88011 95612 88053 95621
rect 88011 95572 88012 95612
rect 88052 95572 88053 95612
rect 88011 95563 88053 95572
rect 79424 95276 79792 95285
rect 79464 95236 79506 95276
rect 79546 95236 79588 95276
rect 79628 95236 79670 95276
rect 79710 95236 79752 95276
rect 79424 95227 79792 95236
rect 78184 94520 78552 94529
rect 78224 94480 78266 94520
rect 78306 94480 78348 94520
rect 78388 94480 78430 94520
rect 78470 94480 78512 94520
rect 78184 94471 78552 94480
rect 79424 93764 79792 93773
rect 79464 93724 79506 93764
rect 79546 93724 79588 93764
rect 79628 93724 79670 93764
rect 79710 93724 79752 93764
rect 79424 93715 79792 93724
rect 78184 93008 78552 93017
rect 78224 92968 78266 93008
rect 78306 92968 78348 93008
rect 78388 92968 78430 93008
rect 78470 92968 78512 93008
rect 78184 92959 78552 92968
rect 79424 92252 79792 92261
rect 79464 92212 79506 92252
rect 79546 92212 79588 92252
rect 79628 92212 79670 92252
rect 79710 92212 79752 92252
rect 79424 92203 79792 92212
rect 78184 91496 78552 91505
rect 78224 91456 78266 91496
rect 78306 91456 78348 91496
rect 78388 91456 78430 91496
rect 78470 91456 78512 91496
rect 78184 91447 78552 91456
rect 79424 90740 79792 90749
rect 79464 90700 79506 90740
rect 79546 90700 79588 90740
rect 79628 90700 79670 90740
rect 79710 90700 79752 90740
rect 79424 90691 79792 90700
rect 78184 89984 78552 89993
rect 78224 89944 78266 89984
rect 78306 89944 78348 89984
rect 78388 89944 78430 89984
rect 78470 89944 78512 89984
rect 78184 89935 78552 89944
rect 79424 89228 79792 89237
rect 79464 89188 79506 89228
rect 79546 89188 79588 89228
rect 79628 89188 79670 89228
rect 79710 89188 79752 89228
rect 79424 89179 79792 89188
rect 78184 88472 78552 88481
rect 78224 88432 78266 88472
rect 78306 88432 78348 88472
rect 78388 88432 78430 88472
rect 78470 88432 78512 88472
rect 78184 88423 78552 88432
rect 79424 87716 79792 87725
rect 79464 87676 79506 87716
rect 79546 87676 79588 87716
rect 79628 87676 79670 87716
rect 79710 87676 79752 87716
rect 79424 87667 79792 87676
rect 78184 86960 78552 86969
rect 78224 86920 78266 86960
rect 78306 86920 78348 86960
rect 78388 86920 78430 86960
rect 78470 86920 78512 86960
rect 78184 86911 78552 86920
rect 79424 86204 79792 86213
rect 79464 86164 79506 86204
rect 79546 86164 79588 86204
rect 79628 86164 79670 86204
rect 79710 86164 79752 86204
rect 79424 86155 79792 86164
rect 78184 85448 78552 85457
rect 78224 85408 78266 85448
rect 78306 85408 78348 85448
rect 78388 85408 78430 85448
rect 78470 85408 78512 85448
rect 78184 85399 78552 85408
rect 79424 84692 79792 84701
rect 79464 84652 79506 84692
rect 79546 84652 79588 84692
rect 79628 84652 79670 84692
rect 79710 84652 79752 84692
rect 79424 84643 79792 84652
rect 78184 83936 78552 83945
rect 78224 83896 78266 83936
rect 78306 83896 78348 83936
rect 78388 83896 78430 83936
rect 78470 83896 78512 83936
rect 78184 83887 78552 83896
rect 79424 83180 79792 83189
rect 79464 83140 79506 83180
rect 79546 83140 79588 83180
rect 79628 83140 79670 83180
rect 79710 83140 79752 83180
rect 79424 83131 79792 83140
rect 78184 82424 78552 82433
rect 78224 82384 78266 82424
rect 78306 82384 78348 82424
rect 78388 82384 78430 82424
rect 78470 82384 78512 82424
rect 78184 82375 78552 82384
rect 79424 81668 79792 81677
rect 79464 81628 79506 81668
rect 79546 81628 79588 81668
rect 79628 81628 79670 81668
rect 79710 81628 79752 81668
rect 79424 81619 79792 81628
rect 78184 80912 78552 80921
rect 78224 80872 78266 80912
rect 78306 80872 78348 80912
rect 78388 80872 78430 80912
rect 78470 80872 78512 80912
rect 78184 80863 78552 80872
rect 79424 80156 79792 80165
rect 79464 80116 79506 80156
rect 79546 80116 79588 80156
rect 79628 80116 79670 80156
rect 79710 80116 79752 80156
rect 79424 80107 79792 80116
rect 78184 79400 78552 79409
rect 78224 79360 78266 79400
rect 78306 79360 78348 79400
rect 78388 79360 78430 79400
rect 78470 79360 78512 79400
rect 78184 79351 78552 79360
rect 79424 78644 79792 78653
rect 79464 78604 79506 78644
rect 79546 78604 79588 78644
rect 79628 78604 79670 78644
rect 79710 78604 79752 78644
rect 79424 78595 79792 78604
rect 78184 77888 78552 77897
rect 78224 77848 78266 77888
rect 78306 77848 78348 77888
rect 78388 77848 78430 77888
rect 78470 77848 78512 77888
rect 78184 77839 78552 77848
rect 79424 77132 79792 77141
rect 79464 77092 79506 77132
rect 79546 77092 79588 77132
rect 79628 77092 79670 77132
rect 79710 77092 79752 77132
rect 79424 77083 79792 77092
rect 78184 76376 78552 76385
rect 78224 76336 78266 76376
rect 78306 76336 78348 76376
rect 78388 76336 78430 76376
rect 78470 76336 78512 76376
rect 78184 76327 78552 76336
rect 79424 75620 79792 75629
rect 79464 75580 79506 75620
rect 79546 75580 79588 75620
rect 79628 75580 79670 75620
rect 79710 75580 79752 75620
rect 79424 75571 79792 75580
rect 88012 64364 88052 95563
rect 93304 94520 93672 94529
rect 93344 94480 93386 94520
rect 93426 94480 93468 94520
rect 93508 94480 93550 94520
rect 93590 94480 93632 94520
rect 93304 94471 93672 94480
rect 93304 93008 93672 93017
rect 93344 92968 93386 93008
rect 93426 92968 93468 93008
rect 93508 92968 93550 93008
rect 93590 92968 93632 93008
rect 93304 92959 93672 92968
rect 93304 91496 93672 91505
rect 93344 91456 93386 91496
rect 93426 91456 93468 91496
rect 93508 91456 93550 91496
rect 93590 91456 93632 91496
rect 93304 91447 93672 91456
rect 93304 89984 93672 89993
rect 93344 89944 93386 89984
rect 93426 89944 93468 89984
rect 93508 89944 93550 89984
rect 93590 89944 93632 89984
rect 93304 89935 93672 89944
rect 93304 88472 93672 88481
rect 93344 88432 93386 88472
rect 93426 88432 93468 88472
rect 93508 88432 93550 88472
rect 93590 88432 93632 88472
rect 93304 88423 93672 88432
rect 93304 86960 93672 86969
rect 93344 86920 93386 86960
rect 93426 86920 93468 86960
rect 93508 86920 93550 86960
rect 93590 86920 93632 86960
rect 93304 86911 93672 86920
rect 93304 85448 93672 85457
rect 93344 85408 93386 85448
rect 93426 85408 93468 85448
rect 93508 85408 93550 85448
rect 93590 85408 93632 85448
rect 93304 85399 93672 85408
rect 93304 83936 93672 83945
rect 93344 83896 93386 83936
rect 93426 83896 93468 83936
rect 93508 83896 93550 83936
rect 93590 83896 93632 83936
rect 93304 83887 93672 83896
rect 93304 82424 93672 82433
rect 93344 82384 93386 82424
rect 93426 82384 93468 82424
rect 93508 82384 93550 82424
rect 93590 82384 93632 82424
rect 93304 82375 93672 82384
rect 93304 80912 93672 80921
rect 93344 80872 93386 80912
rect 93426 80872 93468 80912
rect 93508 80872 93550 80912
rect 93590 80872 93632 80912
rect 93304 80863 93672 80872
rect 93304 79400 93672 79409
rect 93344 79360 93386 79400
rect 93426 79360 93468 79400
rect 93508 79360 93550 79400
rect 93590 79360 93632 79400
rect 93304 79351 93672 79360
rect 93304 77888 93672 77897
rect 93344 77848 93386 77888
rect 93426 77848 93468 77888
rect 93508 77848 93550 77888
rect 93590 77848 93632 77888
rect 93304 77839 93672 77848
rect 93304 76376 93672 76385
rect 93344 76336 93386 76376
rect 93426 76336 93468 76376
rect 93508 76336 93550 76376
rect 93590 76336 93632 76376
rect 93304 76327 93672 76336
rect 93772 71261 93812 122359
rect 94252 89153 94292 126391
rect 94732 125684 94772 126727
rect 94828 126692 94868 126703
rect 94828 126617 94868 126652
rect 94923 126692 94965 126701
rect 94923 126652 94924 126692
rect 94964 126652 94965 126692
rect 94923 126643 94965 126652
rect 94827 126608 94869 126617
rect 94827 126568 94828 126608
rect 94868 126568 94869 126608
rect 94827 126559 94869 126568
rect 94924 126558 94964 126643
rect 95020 126617 95060 127324
rect 95019 126608 95061 126617
rect 95019 126568 95020 126608
rect 95060 126568 95061 126608
rect 95019 126559 95061 126568
rect 94828 126440 94868 126449
rect 95116 126440 95156 127408
rect 95500 126860 95540 128239
rect 98956 128036 98996 129835
rect 99052 128120 99092 130339
rect 99147 130304 99189 130313
rect 99147 130264 99148 130304
rect 99188 130264 99189 130304
rect 99147 130255 99189 130264
rect 99148 128372 99188 130255
rect 99148 128323 99188 128332
rect 99148 128204 99188 128275
rect 99147 128140 99148 128189
rect 99244 128204 99284 131683
rect 99340 131069 99380 131860
rect 99436 131900 99476 132019
rect 100012 131993 100052 132691
rect 101355 132656 101397 132665
rect 101355 132616 101356 132656
rect 101396 132616 101397 132656
rect 101355 132607 101397 132616
rect 101067 132068 101109 132077
rect 101067 132028 101068 132068
rect 101108 132028 101109 132068
rect 101067 132019 101109 132028
rect 99531 131984 99573 131993
rect 99531 131944 99532 131984
rect 99572 131944 99573 131984
rect 99531 131935 99573 131944
rect 100011 131984 100053 131993
rect 100011 131944 100012 131984
rect 100052 131944 100053 131984
rect 100011 131935 100053 131944
rect 99436 131851 99476 131860
rect 99532 131900 99572 131935
rect 99532 131849 99572 131860
rect 100012 131900 100052 131935
rect 100012 131850 100052 131860
rect 100203 131900 100245 131909
rect 100203 131860 100204 131900
rect 100244 131860 100245 131900
rect 100203 131851 100245 131860
rect 101068 131900 101108 132019
rect 101163 131984 101205 131993
rect 101163 131944 101164 131984
rect 101204 131944 101205 131984
rect 101163 131935 101205 131944
rect 101068 131851 101108 131860
rect 101164 131900 101204 131935
rect 101356 131909 101396 132607
rect 100108 131816 100148 131825
rect 99916 131228 99956 131237
rect 99339 131060 99381 131069
rect 99339 131020 99340 131060
rect 99380 131020 99381 131060
rect 99339 131011 99381 131020
rect 99916 130145 99956 131188
rect 99915 130136 99957 130145
rect 99915 130096 99916 130136
rect 99956 130096 99957 130136
rect 99915 130087 99957 130096
rect 99916 129977 99956 130087
rect 99915 129968 99957 129977
rect 99915 129928 99916 129968
rect 99956 129928 99957 129968
rect 99915 129919 99957 129928
rect 100108 129893 100148 131776
rect 100204 131766 100244 131851
rect 101164 131849 101204 131860
rect 101355 131900 101397 131909
rect 101355 131860 101356 131900
rect 101396 131860 101397 131900
rect 101355 131851 101397 131860
rect 101644 131900 101684 131909
rect 101260 131732 101300 131741
rect 101260 131321 101300 131692
rect 101547 131732 101589 131741
rect 101547 131692 101548 131732
rect 101588 131692 101589 131732
rect 101547 131683 101589 131692
rect 101548 131598 101588 131683
rect 101259 131312 101301 131321
rect 101259 131272 101260 131312
rect 101300 131272 101301 131312
rect 101259 131263 101301 131272
rect 100587 131228 100629 131237
rect 100587 131188 100588 131228
rect 100628 131188 100629 131228
rect 100587 131179 100629 131188
rect 100588 131094 100628 131179
rect 101644 130397 101684 131860
rect 102220 131396 102260 132691
rect 102988 132606 103028 132691
rect 103948 131489 103988 158380
rect 109664 148196 110032 148205
rect 109704 148156 109746 148196
rect 109786 148156 109828 148196
rect 109868 148156 109910 148196
rect 109950 148156 109992 148196
rect 109664 148147 110032 148156
rect 108424 147440 108792 147449
rect 108464 147400 108506 147440
rect 108546 147400 108588 147440
rect 108628 147400 108670 147440
rect 108710 147400 108752 147440
rect 108424 147391 108792 147400
rect 109664 146684 110032 146693
rect 109704 146644 109746 146684
rect 109786 146644 109828 146684
rect 109868 146644 109910 146684
rect 109950 146644 109992 146684
rect 109664 146635 110032 146644
rect 108424 145928 108792 145937
rect 108464 145888 108506 145928
rect 108546 145888 108588 145928
rect 108628 145888 108670 145928
rect 108710 145888 108752 145928
rect 108424 145879 108792 145888
rect 109664 145172 110032 145181
rect 109704 145132 109746 145172
rect 109786 145132 109828 145172
rect 109868 145132 109910 145172
rect 109950 145132 109992 145172
rect 109664 145123 110032 145132
rect 108424 144416 108792 144425
rect 108464 144376 108506 144416
rect 108546 144376 108588 144416
rect 108628 144376 108670 144416
rect 108710 144376 108752 144416
rect 108424 144367 108792 144376
rect 109664 143660 110032 143669
rect 109704 143620 109746 143660
rect 109786 143620 109828 143660
rect 109868 143620 109910 143660
rect 109950 143620 109992 143660
rect 109664 143611 110032 143620
rect 108424 142904 108792 142913
rect 108464 142864 108506 142904
rect 108546 142864 108588 142904
rect 108628 142864 108670 142904
rect 108710 142864 108752 142904
rect 108424 142855 108792 142864
rect 109664 142148 110032 142157
rect 109704 142108 109746 142148
rect 109786 142108 109828 142148
rect 109868 142108 109910 142148
rect 109950 142108 109992 142148
rect 109664 142099 110032 142108
rect 108424 141392 108792 141401
rect 108464 141352 108506 141392
rect 108546 141352 108588 141392
rect 108628 141352 108670 141392
rect 108710 141352 108752 141392
rect 108424 141343 108792 141352
rect 109664 140636 110032 140645
rect 109704 140596 109746 140636
rect 109786 140596 109828 140636
rect 109868 140596 109910 140636
rect 109950 140596 109992 140636
rect 109664 140587 110032 140596
rect 108424 139880 108792 139889
rect 108464 139840 108506 139880
rect 108546 139840 108588 139880
rect 108628 139840 108670 139880
rect 108710 139840 108752 139880
rect 108424 139831 108792 139840
rect 109664 139124 110032 139133
rect 109704 139084 109746 139124
rect 109786 139084 109828 139124
rect 109868 139084 109910 139124
rect 109950 139084 109992 139124
rect 109664 139075 110032 139084
rect 108424 138368 108792 138377
rect 108464 138328 108506 138368
rect 108546 138328 108588 138368
rect 108628 138328 108670 138368
rect 108710 138328 108752 138368
rect 108424 138319 108792 138328
rect 109664 137612 110032 137621
rect 109704 137572 109746 137612
rect 109786 137572 109828 137612
rect 109868 137572 109910 137612
rect 109950 137572 109992 137612
rect 109664 137563 110032 137572
rect 108424 136856 108792 136865
rect 108464 136816 108506 136856
rect 108546 136816 108588 136856
rect 108628 136816 108670 136856
rect 108710 136816 108752 136856
rect 108424 136807 108792 136816
rect 109664 136100 110032 136109
rect 109704 136060 109746 136100
rect 109786 136060 109828 136100
rect 109868 136060 109910 136100
rect 109950 136060 109992 136100
rect 109664 136051 110032 136060
rect 108424 135344 108792 135353
rect 108464 135304 108506 135344
rect 108546 135304 108588 135344
rect 108628 135304 108670 135344
rect 108710 135304 108752 135344
rect 108424 135295 108792 135304
rect 109664 134588 110032 134597
rect 109704 134548 109746 134588
rect 109786 134548 109828 134588
rect 109868 134548 109910 134588
rect 109950 134548 109992 134588
rect 109664 134539 110032 134548
rect 105099 134252 105141 134261
rect 105099 134212 105100 134252
rect 105140 134212 105141 134252
rect 105099 134203 105141 134212
rect 104236 132740 104276 132749
rect 104236 132068 104276 132700
rect 105100 132740 105140 134203
rect 108424 133832 108792 133841
rect 108464 133792 108506 133832
rect 108546 133792 108588 133832
rect 108628 133792 108670 133832
rect 108710 133792 108752 133832
rect 108424 133783 108792 133792
rect 109664 133076 110032 133085
rect 109704 133036 109746 133076
rect 109786 133036 109828 133076
rect 109868 133036 109910 133076
rect 109950 133036 109992 133076
rect 109664 133027 110032 133036
rect 104332 132068 104372 132077
rect 104236 132028 104332 132068
rect 104332 132019 104372 132028
rect 103947 131480 103989 131489
rect 103947 131440 103948 131480
rect 103988 131440 103989 131480
rect 103947 131431 103989 131440
rect 102220 131347 102260 131356
rect 103084 131356 103412 131396
rect 102123 131312 102165 131321
rect 102123 131272 102124 131312
rect 102164 131272 102165 131312
rect 102123 131263 102165 131272
rect 102027 131228 102069 131237
rect 102027 131188 102028 131228
rect 102068 131188 102069 131228
rect 102027 131179 102069 131188
rect 102124 131228 102164 131263
rect 102028 131094 102068 131179
rect 102124 131177 102164 131188
rect 102316 131228 102356 131237
rect 102219 131060 102261 131069
rect 102219 131020 102220 131060
rect 102260 131020 102261 131060
rect 102219 131011 102261 131020
rect 102220 130472 102260 131011
rect 102316 130640 102356 131188
rect 102508 130976 102548 130985
rect 102548 130936 103028 130976
rect 102508 130927 102548 130936
rect 102604 130640 102644 130649
rect 102316 130600 102604 130640
rect 102644 130600 102836 130640
rect 102604 130591 102644 130600
rect 102220 130432 102548 130472
rect 101643 130388 101685 130397
rect 101643 130348 101644 130388
rect 101684 130348 101685 130388
rect 101643 130339 101685 130348
rect 102508 130388 102548 130432
rect 102508 130339 102548 130348
rect 102796 130388 102836 130600
rect 102796 130339 102836 130348
rect 102988 130388 103028 130936
rect 103084 130556 103124 131356
rect 103084 130507 103124 130516
rect 103180 131228 103220 131237
rect 102988 130339 103028 130348
rect 103084 130388 103124 130399
rect 103084 130313 103124 130348
rect 103083 130304 103125 130313
rect 103083 130264 103084 130304
rect 103124 130264 103125 130304
rect 103083 130255 103125 130264
rect 100107 129884 100149 129893
rect 100107 129844 100108 129884
rect 100148 129844 100149 129884
rect 100107 129835 100149 129844
rect 103083 129884 103125 129893
rect 103083 129844 103084 129884
rect 103124 129844 103125 129884
rect 103083 129835 103125 129844
rect 103180 129884 103220 131188
rect 103372 131228 103412 131356
rect 103372 131179 103412 131188
rect 103467 131228 103509 131237
rect 103467 131188 103468 131228
rect 103508 131188 103509 131228
rect 103467 131179 103509 131188
rect 103468 130313 103508 131179
rect 104331 131144 104373 131153
rect 104331 131104 104332 131144
rect 104372 131104 104373 131144
rect 104331 131095 104373 131104
rect 103563 131060 103605 131069
rect 103563 131020 103564 131060
rect 103604 131020 103605 131060
rect 103563 131011 103605 131020
rect 104043 131060 104085 131069
rect 104043 131020 104044 131060
rect 104084 131020 104085 131060
rect 104043 131011 104085 131020
rect 103467 130304 103509 130313
rect 103467 130264 103468 130304
rect 103508 130264 103509 130304
rect 103467 130255 103509 130264
rect 103275 130220 103317 130229
rect 103275 130180 103276 130220
rect 103316 130180 103317 130220
rect 103275 130171 103317 130180
rect 103180 129835 103220 129844
rect 103084 129716 103124 129835
rect 103084 129667 103124 129676
rect 103276 129716 103316 130171
rect 103564 129800 103604 131011
rect 104044 130926 104084 131011
rect 103564 129751 103604 129760
rect 103276 129667 103316 129676
rect 103948 129716 103988 129725
rect 103948 129044 103988 129676
rect 104044 129044 104084 129053
rect 103948 129004 104044 129044
rect 104044 128995 104084 129004
rect 99188 128140 99189 128189
rect 99244 128155 99284 128164
rect 99147 128131 99189 128140
rect 99052 128071 99092 128080
rect 98956 127987 98996 127996
rect 95500 126811 95540 126820
rect 95559 126692 95599 126701
rect 95559 126533 95599 126652
rect 95672 126692 95712 126701
rect 95788 126692 95828 126703
rect 95712 126652 95732 126692
rect 95672 126643 95732 126652
rect 95559 126524 95637 126533
rect 95559 126484 95596 126524
rect 95636 126484 95637 126524
rect 95595 126475 95637 126484
rect 95692 126449 95732 126643
rect 95788 126617 95828 126652
rect 95883 126692 95925 126701
rect 95883 126652 95884 126692
rect 95924 126652 95925 126692
rect 95883 126643 95925 126652
rect 95787 126608 95829 126617
rect 95787 126568 95788 126608
rect 95828 126568 95829 126608
rect 95787 126559 95829 126568
rect 95884 126558 95924 126643
rect 104043 126608 104085 126617
rect 104043 126568 104044 126608
rect 104084 126568 104085 126608
rect 104043 126559 104085 126568
rect 94868 126400 95156 126440
rect 95691 126440 95733 126449
rect 95691 126400 95692 126440
rect 95732 126400 95733 126440
rect 94828 126391 94868 126400
rect 95691 126391 95733 126400
rect 94444 125644 94772 125684
rect 94444 105029 94484 125644
rect 94544 125516 94912 125525
rect 94584 125476 94626 125516
rect 94666 125476 94708 125516
rect 94748 125476 94790 125516
rect 94830 125476 94872 125516
rect 94544 125467 94912 125476
rect 94544 124004 94912 124013
rect 94584 123964 94626 124004
rect 94666 123964 94708 124004
rect 94748 123964 94790 124004
rect 94830 123964 94872 124004
rect 94544 123955 94912 123964
rect 94544 122492 94912 122501
rect 94584 122452 94626 122492
rect 94666 122452 94708 122492
rect 94748 122452 94790 122492
rect 94830 122452 94872 122492
rect 94544 122443 94912 122452
rect 94544 120980 94912 120989
rect 94584 120940 94626 120980
rect 94666 120940 94708 120980
rect 94748 120940 94790 120980
rect 94830 120940 94872 120980
rect 94544 120931 94912 120940
rect 94544 119468 94912 119477
rect 94584 119428 94626 119468
rect 94666 119428 94708 119468
rect 94748 119428 94790 119468
rect 94830 119428 94872 119468
rect 94544 119419 94912 119428
rect 94544 117956 94912 117965
rect 94584 117916 94626 117956
rect 94666 117916 94708 117956
rect 94748 117916 94790 117956
rect 94830 117916 94872 117956
rect 94544 117907 94912 117916
rect 94544 116444 94912 116453
rect 94584 116404 94626 116444
rect 94666 116404 94708 116444
rect 94748 116404 94790 116444
rect 94830 116404 94872 116444
rect 94544 116395 94912 116404
rect 94544 114932 94912 114941
rect 94584 114892 94626 114932
rect 94666 114892 94708 114932
rect 94748 114892 94790 114932
rect 94830 114892 94872 114932
rect 94544 114883 94912 114892
rect 94544 113420 94912 113429
rect 94584 113380 94626 113420
rect 94666 113380 94708 113420
rect 94748 113380 94790 113420
rect 94830 113380 94872 113420
rect 94544 113371 94912 113380
rect 94544 111908 94912 111917
rect 94584 111868 94626 111908
rect 94666 111868 94708 111908
rect 94748 111868 94790 111908
rect 94830 111868 94872 111908
rect 94544 111859 94912 111868
rect 94544 110396 94912 110405
rect 94584 110356 94626 110396
rect 94666 110356 94708 110396
rect 94748 110356 94790 110396
rect 94830 110356 94872 110396
rect 94544 110347 94912 110356
rect 94544 108884 94912 108893
rect 94584 108844 94626 108884
rect 94666 108844 94708 108884
rect 94748 108844 94790 108884
rect 94830 108844 94872 108884
rect 94544 108835 94912 108844
rect 94544 107372 94912 107381
rect 94584 107332 94626 107372
rect 94666 107332 94708 107372
rect 94748 107332 94790 107372
rect 94830 107332 94872 107372
rect 94544 107323 94912 107332
rect 94544 105860 94912 105869
rect 94584 105820 94626 105860
rect 94666 105820 94708 105860
rect 94748 105820 94790 105860
rect 94830 105820 94872 105860
rect 94544 105811 94912 105820
rect 94443 105020 94485 105029
rect 94443 104980 94444 105020
rect 94484 104980 94485 105020
rect 94443 104971 94485 104980
rect 94544 104348 94912 104357
rect 94584 104308 94626 104348
rect 94666 104308 94708 104348
rect 94748 104308 94790 104348
rect 94830 104308 94872 104348
rect 94544 104299 94912 104308
rect 94544 102836 94912 102845
rect 94584 102796 94626 102836
rect 94666 102796 94708 102836
rect 94748 102796 94790 102836
rect 94830 102796 94872 102836
rect 94544 102787 94912 102796
rect 94544 101324 94912 101333
rect 94584 101284 94626 101324
rect 94666 101284 94708 101324
rect 94748 101284 94790 101324
rect 94830 101284 94872 101324
rect 94544 101275 94912 101284
rect 94544 99812 94912 99821
rect 94584 99772 94626 99812
rect 94666 99772 94708 99812
rect 94748 99772 94790 99812
rect 94830 99772 94872 99812
rect 94544 99763 94912 99772
rect 94544 98300 94912 98309
rect 94584 98260 94626 98300
rect 94666 98260 94708 98300
rect 94748 98260 94790 98300
rect 94830 98260 94872 98300
rect 94544 98251 94912 98260
rect 94544 96788 94912 96797
rect 94584 96748 94626 96788
rect 94666 96748 94708 96788
rect 94748 96748 94790 96788
rect 94830 96748 94872 96788
rect 94544 96739 94912 96748
rect 103659 95612 103701 95621
rect 103659 95572 103660 95612
rect 103700 95572 103701 95612
rect 103659 95563 103701 95572
rect 103660 95478 103700 95563
rect 94544 95276 94912 95285
rect 94584 95236 94626 95276
rect 94666 95236 94708 95276
rect 94748 95236 94790 95276
rect 94830 95236 94872 95276
rect 94544 95227 94912 95236
rect 94544 93764 94912 93773
rect 94584 93724 94626 93764
rect 94666 93724 94708 93764
rect 94748 93724 94790 93764
rect 94830 93724 94872 93764
rect 94544 93715 94912 93724
rect 94544 92252 94912 92261
rect 94584 92212 94626 92252
rect 94666 92212 94708 92252
rect 94748 92212 94790 92252
rect 94830 92212 94872 92252
rect 94544 92203 94912 92212
rect 94544 90740 94912 90749
rect 94584 90700 94626 90740
rect 94666 90700 94708 90740
rect 94748 90700 94790 90740
rect 94830 90700 94872 90740
rect 94544 90691 94912 90700
rect 94544 89228 94912 89237
rect 94584 89188 94626 89228
rect 94666 89188 94708 89228
rect 94748 89188 94790 89228
rect 94830 89188 94872 89228
rect 94544 89179 94912 89188
rect 94251 89144 94293 89153
rect 94251 89104 94252 89144
rect 94292 89104 94293 89144
rect 94251 89095 94293 89104
rect 94544 87716 94912 87725
rect 94584 87676 94626 87716
rect 94666 87676 94708 87716
rect 94748 87676 94790 87716
rect 94830 87676 94872 87716
rect 94544 87667 94912 87676
rect 94544 86204 94912 86213
rect 94584 86164 94626 86204
rect 94666 86164 94708 86204
rect 94748 86164 94790 86204
rect 94830 86164 94872 86204
rect 94544 86155 94912 86164
rect 94544 84692 94912 84701
rect 94584 84652 94626 84692
rect 94666 84652 94708 84692
rect 94748 84652 94790 84692
rect 94830 84652 94872 84692
rect 94544 84643 94912 84652
rect 94544 83180 94912 83189
rect 94584 83140 94626 83180
rect 94666 83140 94708 83180
rect 94748 83140 94790 83180
rect 94830 83140 94872 83180
rect 94544 83131 94912 83140
rect 94544 81668 94912 81677
rect 94584 81628 94626 81668
rect 94666 81628 94708 81668
rect 94748 81628 94790 81668
rect 94830 81628 94872 81668
rect 94544 81619 94912 81628
rect 94544 80156 94912 80165
rect 94584 80116 94626 80156
rect 94666 80116 94708 80156
rect 94748 80116 94790 80156
rect 94830 80116 94872 80156
rect 94544 80107 94912 80116
rect 94544 78644 94912 78653
rect 94584 78604 94626 78644
rect 94666 78604 94708 78644
rect 94748 78604 94790 78644
rect 94830 78604 94872 78644
rect 94544 78595 94912 78604
rect 94544 77132 94912 77141
rect 94584 77092 94626 77132
rect 94666 77092 94708 77132
rect 94748 77092 94790 77132
rect 94830 77092 94872 77132
rect 94544 77083 94912 77092
rect 94544 75620 94912 75629
rect 94584 75580 94626 75620
rect 94666 75580 94708 75620
rect 94748 75580 94790 75620
rect 94830 75580 94872 75620
rect 94544 75571 94912 75580
rect 93771 71252 93813 71261
rect 93771 71212 93772 71252
rect 93812 71212 93813 71252
rect 93771 71203 93813 71212
rect 104044 64364 104084 126559
rect 104332 95864 104372 131095
rect 105100 130733 105140 132700
rect 106251 132656 106293 132665
rect 106251 132616 106252 132656
rect 106292 132616 106293 132656
rect 106251 132607 106293 132616
rect 106252 132522 106292 132607
rect 109900 132572 109940 132581
rect 109804 132532 109900 132572
rect 108424 132320 108792 132329
rect 108464 132280 108506 132320
rect 108546 132280 108588 132320
rect 108628 132280 108670 132320
rect 108710 132280 108752 132320
rect 108424 132271 108792 132280
rect 109804 131900 109844 132532
rect 109900 132523 109940 132532
rect 109804 131851 109844 131860
rect 110668 131900 110708 131909
rect 109420 131816 109460 131825
rect 108747 131648 108789 131657
rect 108747 131608 108748 131648
rect 108788 131608 108789 131648
rect 108747 131599 108789 131608
rect 108748 131153 108788 131599
rect 109420 131405 109460 131776
rect 109664 131564 110032 131573
rect 109704 131524 109746 131564
rect 109786 131524 109828 131564
rect 109868 131524 109910 131564
rect 109950 131524 109992 131564
rect 109664 131515 110032 131524
rect 108844 131396 108884 131405
rect 109419 131396 109461 131405
rect 108884 131356 109364 131396
rect 108844 131347 108884 131356
rect 108940 131228 108980 131239
rect 108940 131153 108980 131188
rect 109035 131228 109077 131237
rect 109035 131188 109036 131228
rect 109076 131188 109077 131228
rect 109035 131179 109077 131188
rect 109132 131228 109172 131239
rect 108747 131144 108789 131153
rect 108747 131104 108748 131144
rect 108788 131104 108789 131144
rect 108747 131095 108789 131104
rect 108939 131144 108981 131153
rect 108939 131104 108940 131144
rect 108980 131104 108981 131144
rect 108939 131095 108981 131104
rect 109036 131094 109076 131179
rect 109132 131153 109172 131188
rect 109324 131228 109364 131356
rect 109419 131356 109420 131396
rect 109460 131356 109461 131396
rect 109419 131347 109461 131356
rect 109803 131396 109845 131405
rect 109803 131356 109804 131396
rect 109844 131356 109845 131396
rect 109803 131347 109845 131356
rect 110379 131396 110421 131405
rect 110379 131356 110380 131396
rect 110420 131356 110421 131396
rect 110379 131347 110421 131356
rect 109804 131262 109844 131347
rect 109324 131179 109364 131188
rect 109419 131228 109461 131237
rect 109419 131188 109420 131228
rect 109460 131188 109461 131228
rect 109419 131179 109461 131188
rect 109612 131228 109652 131237
rect 109131 131144 109173 131153
rect 109131 131104 109132 131144
rect 109172 131104 109173 131144
rect 109131 131095 109173 131104
rect 109420 131094 109460 131179
rect 109612 131069 109652 131188
rect 110380 131153 110420 131347
rect 110475 131228 110517 131237
rect 110475 131188 110476 131228
rect 110516 131188 110517 131228
rect 110475 131179 110517 131188
rect 110379 131144 110421 131153
rect 110379 131104 110380 131144
rect 110420 131104 110421 131144
rect 110379 131095 110421 131104
rect 109611 131060 109653 131069
rect 109611 131020 109612 131060
rect 109652 131020 109653 131060
rect 109611 131011 109653 131020
rect 108424 130808 108792 130817
rect 108464 130768 108506 130808
rect 108546 130768 108588 130808
rect 108628 130768 108670 130808
rect 108710 130768 108752 130808
rect 108424 130759 108792 130768
rect 105099 130724 105141 130733
rect 105099 130684 105100 130724
rect 105140 130684 105141 130724
rect 105099 130675 105141 130684
rect 104715 130220 104757 130229
rect 104715 130180 104716 130220
rect 104756 130180 104757 130220
rect 104715 130171 104757 130180
rect 104716 130086 104756 130171
rect 104812 129716 104852 129725
rect 105100 129716 105140 130675
rect 108747 130640 108789 130649
rect 108747 130600 108748 130640
rect 108788 130600 108789 130640
rect 108747 130591 108789 130600
rect 108748 130472 108788 130591
rect 108748 130423 108788 130432
rect 105387 130388 105429 130397
rect 105387 130348 105388 130388
rect 105428 130348 105429 130388
rect 105387 130339 105429 130348
rect 105963 130388 106005 130397
rect 105963 130348 105964 130388
rect 106004 130348 106005 130388
rect 105963 130339 106005 130348
rect 110187 130388 110229 130397
rect 110187 130348 110188 130388
rect 110228 130348 110229 130388
rect 110380 130388 110420 131095
rect 110476 131094 110516 131179
rect 110571 131060 110613 131069
rect 110571 131020 110572 131060
rect 110612 131020 110613 131060
rect 110571 131011 110613 131020
rect 110476 130640 110516 130649
rect 110572 130640 110612 131011
rect 110668 130649 110708 131860
rect 112204 131900 112244 131909
rect 110763 131816 110805 131825
rect 110763 131776 110764 131816
rect 110804 131776 110805 131816
rect 110763 131767 110805 131776
rect 110764 131405 110804 131767
rect 111820 131732 111860 131741
rect 111820 131489 111860 131692
rect 111435 131480 111477 131489
rect 111435 131440 111436 131480
rect 111476 131440 111477 131480
rect 111435 131431 111477 131440
rect 111819 131480 111861 131489
rect 111819 131440 111820 131480
rect 111860 131440 111861 131480
rect 111819 131431 111861 131440
rect 110763 131396 110805 131405
rect 110763 131356 110764 131396
rect 110804 131356 110805 131396
rect 110763 131347 110805 131356
rect 110764 131262 110804 131347
rect 111436 131228 111476 131431
rect 111436 131179 111476 131188
rect 112204 130985 112244 131860
rect 112300 131900 112340 159655
rect 115947 151640 115989 151649
rect 115947 151600 115948 151640
rect 115988 151600 115989 151640
rect 115947 151591 115989 151600
rect 115948 134420 115988 151591
rect 124784 148196 125152 148205
rect 124824 148156 124866 148196
rect 124906 148156 124948 148196
rect 124988 148156 125030 148196
rect 125070 148156 125112 148196
rect 124784 148147 125152 148156
rect 123544 147440 123912 147449
rect 123584 147400 123626 147440
rect 123666 147400 123708 147440
rect 123748 147400 123790 147440
rect 123830 147400 123872 147440
rect 123544 147391 123912 147400
rect 124784 146684 125152 146693
rect 124824 146644 124866 146684
rect 124906 146644 124948 146684
rect 124988 146644 125030 146684
rect 125070 146644 125112 146684
rect 124784 146635 125152 146644
rect 123544 145928 123912 145937
rect 123584 145888 123626 145928
rect 123666 145888 123708 145928
rect 123748 145888 123790 145928
rect 123830 145888 123872 145928
rect 123544 145879 123912 145888
rect 124784 145172 125152 145181
rect 124824 145132 124866 145172
rect 124906 145132 124948 145172
rect 124988 145132 125030 145172
rect 125070 145132 125112 145172
rect 124784 145123 125152 145132
rect 123544 144416 123912 144425
rect 123584 144376 123626 144416
rect 123666 144376 123708 144416
rect 123748 144376 123790 144416
rect 123830 144376 123872 144416
rect 123544 144367 123912 144376
rect 124784 143660 125152 143669
rect 124824 143620 124866 143660
rect 124906 143620 124948 143660
rect 124988 143620 125030 143660
rect 125070 143620 125112 143660
rect 124784 143611 125152 143620
rect 123544 142904 123912 142913
rect 123584 142864 123626 142904
rect 123666 142864 123708 142904
rect 123748 142864 123790 142904
rect 123830 142864 123872 142904
rect 123544 142855 123912 142864
rect 124784 142148 125152 142157
rect 124824 142108 124866 142148
rect 124906 142108 124948 142148
rect 124988 142108 125030 142148
rect 125070 142108 125112 142148
rect 124784 142099 125152 142108
rect 123544 141392 123912 141401
rect 123584 141352 123626 141392
rect 123666 141352 123708 141392
rect 123748 141352 123790 141392
rect 123830 141352 123872 141392
rect 123544 141343 123912 141352
rect 124784 140636 125152 140645
rect 124824 140596 124866 140636
rect 124906 140596 124948 140636
rect 124988 140596 125030 140636
rect 125070 140596 125112 140636
rect 124784 140587 125152 140596
rect 123544 139880 123912 139889
rect 123584 139840 123626 139880
rect 123666 139840 123708 139880
rect 123748 139840 123790 139880
rect 123830 139840 123872 139880
rect 123544 139831 123912 139840
rect 124784 139124 125152 139133
rect 124824 139084 124866 139124
rect 124906 139084 124948 139124
rect 124988 139084 125030 139124
rect 125070 139084 125112 139124
rect 124784 139075 125152 139084
rect 123544 138368 123912 138377
rect 123584 138328 123626 138368
rect 123666 138328 123708 138368
rect 123748 138328 123790 138368
rect 123830 138328 123872 138368
rect 123544 138319 123912 138328
rect 124784 137612 125152 137621
rect 124824 137572 124866 137612
rect 124906 137572 124948 137612
rect 124988 137572 125030 137612
rect 125070 137572 125112 137612
rect 124784 137563 125152 137572
rect 123544 136856 123912 136865
rect 123584 136816 123626 136856
rect 123666 136816 123708 136856
rect 123748 136816 123790 136856
rect 123830 136816 123872 136856
rect 123544 136807 123912 136816
rect 124784 136100 125152 136109
rect 124824 136060 124866 136100
rect 124906 136060 124948 136100
rect 124988 136060 125030 136100
rect 125070 136060 125112 136100
rect 124784 136051 125152 136060
rect 121803 135596 121845 135605
rect 121803 135556 121804 135596
rect 121844 135556 121845 135596
rect 121803 135547 121845 135556
rect 115948 134371 115988 134380
rect 113548 134252 113588 134261
rect 113356 134212 113548 134252
rect 112875 133244 112917 133253
rect 112875 133204 112876 133244
rect 112916 133204 112917 133244
rect 112875 133195 112917 133204
rect 112300 131816 112340 131860
rect 112780 131900 112820 131909
rect 112297 131776 112340 131816
rect 112395 131816 112444 131825
rect 112395 131776 112396 131816
rect 112297 131732 112337 131776
rect 112395 131767 112444 131776
rect 112297 131692 112340 131732
rect 112300 131564 112340 131692
rect 112404 131689 112444 131767
rect 112588 131741 112628 131826
rect 112492 131732 112532 131741
rect 112492 131573 112532 131692
rect 112587 131732 112629 131741
rect 112587 131692 112588 131732
rect 112628 131692 112629 131732
rect 112587 131683 112629 131692
rect 112491 131564 112533 131573
rect 112300 131524 112436 131564
rect 112299 131396 112341 131405
rect 112299 131356 112300 131396
rect 112340 131356 112341 131396
rect 112299 131347 112341 131356
rect 112300 131262 112340 131347
rect 110763 130976 110805 130985
rect 110763 130936 110764 130976
rect 110804 130936 110805 130976
rect 110763 130927 110805 130936
rect 112203 130976 112245 130985
rect 112203 130936 112204 130976
rect 112244 130936 112245 130976
rect 112203 130927 112245 130936
rect 110516 130600 110612 130640
rect 110667 130640 110709 130649
rect 110667 130600 110668 130640
rect 110708 130600 110709 130640
rect 110476 130591 110516 130600
rect 110667 130591 110709 130600
rect 110476 130388 110516 130397
rect 110380 130348 110476 130388
rect 110187 130339 110229 130348
rect 110476 130339 110516 130348
rect 110668 130388 110708 130397
rect 105388 130254 105428 130339
rect 105964 130229 106004 130339
rect 110188 130254 110228 130339
rect 110668 130229 110708 130348
rect 110764 130388 110804 130927
rect 105963 130220 106005 130229
rect 105963 130180 105964 130220
rect 106004 130180 106005 130220
rect 105963 130171 106005 130180
rect 110667 130220 110709 130229
rect 110667 130180 110668 130220
rect 110708 130180 110709 130220
rect 110667 130171 110709 130180
rect 105964 129884 106004 130171
rect 109664 130052 110032 130061
rect 109704 130012 109746 130052
rect 109786 130012 109828 130052
rect 109868 130012 109910 130052
rect 109950 130012 109992 130052
rect 109664 130003 110032 130012
rect 110764 129893 110804 130348
rect 112011 130388 112053 130397
rect 112011 130348 112012 130388
rect 112052 130348 112053 130388
rect 112011 130339 112053 130348
rect 105964 129835 106004 129844
rect 110763 129884 110805 129893
rect 110763 129844 110764 129884
rect 110804 129844 110805 129884
rect 110763 129835 110805 129844
rect 112012 129725 112052 130339
rect 112396 130229 112436 131524
rect 112491 131524 112492 131564
rect 112532 131524 112533 131564
rect 112491 131515 112533 131524
rect 112780 131405 112820 131860
rect 112779 131396 112821 131405
rect 112779 131356 112780 131396
rect 112820 131356 112821 131396
rect 112779 131347 112821 131356
rect 112492 131228 112532 131237
rect 112492 131069 112532 131188
rect 112588 131228 112628 131237
rect 112876 131228 112916 133195
rect 113163 131732 113205 131741
rect 113163 131692 113164 131732
rect 113204 131692 113205 131732
rect 113163 131683 113205 131692
rect 113067 131648 113109 131657
rect 113067 131608 113068 131648
rect 113108 131608 113109 131648
rect 113067 131599 113109 131608
rect 113068 131396 113108 131599
rect 112628 131188 112916 131228
rect 112972 131356 113068 131396
rect 112588 131179 112628 131188
rect 112491 131060 112533 131069
rect 112491 131020 112492 131060
rect 112532 131020 112533 131060
rect 112491 131011 112533 131020
rect 112972 130481 113012 131356
rect 113068 131347 113108 131356
rect 113164 131237 113204 131683
rect 113356 131312 113396 134212
rect 113548 134203 113588 134212
rect 113932 134252 113972 134261
rect 113932 133580 113972 134212
rect 114796 134252 114836 134261
rect 114028 133580 114068 133589
rect 113932 133540 114028 133580
rect 114028 133531 114068 133540
rect 114796 133421 114836 134212
rect 119884 134084 119924 134093
rect 119788 134044 119884 134084
rect 115083 134000 115125 134009
rect 115083 133960 115084 134000
rect 115124 133960 115125 134000
rect 115083 133951 115125 133960
rect 115947 134000 115989 134009
rect 115947 133960 115948 134000
rect 115988 133960 115989 134000
rect 115947 133951 115989 133960
rect 114795 133412 114837 133421
rect 114795 133372 114796 133412
rect 114836 133372 114837 133412
rect 114795 133363 114837 133372
rect 115084 133412 115124 133951
rect 115948 133866 115988 133951
rect 114411 133244 114453 133253
rect 114411 133204 114412 133244
rect 114452 133204 114453 133244
rect 114411 133195 114453 133204
rect 114412 133110 114452 133195
rect 113356 131263 113396 131272
rect 113452 131732 113492 131741
rect 113068 131228 113108 131237
rect 113068 131060 113108 131188
rect 113163 131228 113205 131237
rect 113163 131188 113164 131228
rect 113204 131188 113205 131228
rect 113163 131179 113205 131188
rect 113452 131060 113492 131692
rect 113068 131020 113492 131060
rect 112971 130472 113013 130481
rect 112971 130432 112972 130472
rect 113012 130432 113013 130472
rect 112971 130423 113013 130432
rect 112395 130220 112437 130229
rect 112395 130180 112396 130220
rect 112436 130180 112437 130220
rect 112395 130171 112437 130180
rect 104852 129676 105140 129716
rect 110571 129716 110613 129725
rect 110571 129676 110572 129716
rect 110612 129676 110613 129716
rect 104812 129667 104852 129676
rect 110571 129667 110613 129676
rect 112011 129716 112053 129725
rect 112011 129676 112012 129716
rect 112052 129676 112053 129716
rect 112011 129667 112053 129676
rect 113931 129716 113973 129725
rect 113931 129676 113932 129716
rect 113972 129676 113973 129716
rect 114796 129716 114836 133363
rect 115084 131573 115124 133372
rect 119788 133412 119828 134044
rect 119884 134035 119924 134044
rect 121804 133664 121844 135547
rect 123544 135344 123912 135353
rect 123584 135304 123626 135344
rect 123666 135304 123708 135344
rect 123748 135304 123790 135344
rect 123830 135304 123872 135344
rect 123544 135295 123912 135304
rect 124784 134588 125152 134597
rect 124824 134548 124866 134588
rect 124906 134548 124948 134588
rect 124988 134548 125030 134588
rect 125070 134548 125112 134588
rect 124784 134539 125152 134548
rect 123544 133832 123912 133841
rect 123584 133792 123626 133832
rect 123666 133792 123708 133832
rect 123748 133792 123790 133832
rect 123830 133792 123872 133832
rect 123544 133783 123912 133792
rect 121804 133615 121844 133624
rect 119788 133363 119828 133372
rect 120459 133412 120501 133421
rect 120459 133372 120460 133412
rect 120500 133372 120501 133412
rect 120459 133363 120501 133372
rect 120651 133412 120693 133421
rect 120651 133372 120652 133412
rect 120692 133372 120693 133412
rect 120651 133363 120693 133372
rect 119404 133328 119444 133337
rect 119404 132908 119444 133288
rect 119404 132859 119444 132868
rect 115179 132824 115221 132833
rect 115179 132784 115180 132824
rect 115220 132784 115221 132824
rect 115179 132775 115221 132784
rect 115083 131564 115125 131573
rect 115083 131524 115084 131564
rect 115124 131524 115125 131564
rect 115083 131515 115125 131524
rect 114987 131480 115029 131489
rect 114987 131440 114988 131480
rect 115028 131440 115029 131480
rect 114987 131431 115029 131440
rect 114891 131228 114933 131237
rect 114891 131188 114892 131228
rect 114932 131188 114933 131228
rect 114891 131179 114933 131188
rect 114988 131228 115028 131431
rect 115084 131312 115124 131515
rect 115180 131396 115220 132775
rect 119307 132740 119349 132749
rect 119307 132700 119308 132740
rect 119348 132700 119349 132740
rect 119307 132691 119349 132700
rect 120075 132740 120117 132749
rect 120075 132700 120076 132740
rect 120116 132700 120117 132740
rect 120075 132691 120117 132700
rect 118539 132572 118581 132581
rect 118539 132532 118540 132572
rect 118580 132532 118581 132572
rect 118539 132523 118581 132532
rect 118540 131900 118580 132523
rect 118540 131851 118580 131860
rect 115180 131347 115220 131356
rect 118444 131732 118484 131741
rect 115084 131263 115124 131272
rect 118251 131312 118293 131321
rect 118251 131272 118252 131312
rect 118292 131272 118293 131312
rect 118251 131263 118293 131272
rect 114988 131179 115028 131188
rect 117579 131228 117621 131237
rect 117579 131188 117580 131228
rect 117620 131188 117621 131228
rect 117579 131179 117621 131188
rect 114892 131094 114932 131179
rect 115180 130976 115220 130985
rect 115180 130397 115220 130936
rect 117580 130640 117620 131179
rect 118252 131153 118292 131263
rect 118251 131144 118293 131153
rect 118251 131104 118252 131144
rect 118292 131104 118293 131144
rect 118251 131095 118293 131104
rect 117580 130591 117620 130600
rect 117675 130472 117717 130481
rect 117675 130432 117676 130472
rect 117716 130432 117717 130472
rect 117675 130423 117717 130432
rect 115179 130388 115221 130397
rect 115179 130348 115180 130388
rect 115220 130348 115221 130388
rect 115179 130339 115221 130348
rect 117483 130388 117525 130397
rect 117483 130348 117484 130388
rect 117524 130348 117525 130388
rect 117483 130339 117525 130348
rect 117676 130388 117716 130423
rect 117484 130254 117524 130339
rect 117676 130337 117716 130348
rect 115372 129716 115412 129725
rect 114796 129676 115372 129716
rect 113931 129667 113973 129676
rect 115372 129667 115412 129676
rect 110572 129582 110612 129667
rect 112012 129582 112052 129667
rect 113932 129582 113972 129667
rect 108424 129296 108792 129305
rect 108464 129256 108506 129296
rect 108546 129256 108588 129296
rect 108628 129256 108670 129296
rect 108710 129256 108752 129296
rect 108424 129247 108792 129256
rect 109664 128540 110032 128549
rect 109704 128500 109746 128540
rect 109786 128500 109828 128540
rect 109868 128500 109910 128540
rect 109950 128500 109992 128540
rect 109664 128491 110032 128500
rect 118252 128204 118292 131095
rect 118252 128155 118292 128164
rect 118444 131060 118484 131692
rect 119308 131396 119348 132691
rect 120076 132606 120116 132691
rect 120267 132572 120309 132581
rect 120267 132532 120268 132572
rect 120308 132532 120309 132572
rect 120267 132523 120309 132532
rect 120268 132438 120308 132523
rect 119308 131347 119348 131356
rect 119115 131312 119157 131321
rect 119115 131272 119116 131312
rect 119156 131272 119157 131312
rect 119115 131263 119157 131272
rect 119116 131228 119156 131263
rect 119404 131237 119444 131322
rect 119116 131177 119156 131188
rect 119212 131228 119252 131237
rect 119212 131060 119252 131188
rect 119403 131228 119445 131237
rect 119403 131188 119404 131228
rect 119444 131188 119445 131228
rect 119403 131179 119445 131188
rect 118444 131020 119252 131060
rect 118444 128202 118484 131020
rect 119211 130472 119253 130481
rect 119211 130432 119212 130472
rect 119252 130432 119253 130472
rect 119211 130423 119253 130432
rect 119115 130388 119157 130397
rect 119115 130348 119116 130388
rect 119156 130348 119157 130388
rect 119115 130339 119157 130348
rect 118540 128297 118580 128299
rect 119020 128297 119060 128299
rect 118539 128288 118581 128297
rect 118539 128248 118540 128288
rect 118580 128248 118581 128288
rect 118539 128239 118581 128248
rect 118731 128288 118773 128297
rect 118731 128248 118732 128288
rect 118772 128248 118773 128288
rect 118731 128239 118773 128248
rect 119019 128288 119061 128297
rect 119019 128248 119020 128288
rect 119060 128248 119061 128288
rect 119019 128239 119061 128248
rect 118444 128153 118484 128162
rect 118540 128204 118580 128239
rect 118540 128155 118580 128164
rect 118636 128204 118676 128213
rect 108424 127784 108792 127793
rect 108464 127744 108506 127784
rect 108546 127744 108588 127784
rect 108628 127744 108670 127784
rect 108710 127744 108752 127784
rect 108424 127735 108792 127744
rect 118636 127196 118676 128164
rect 118732 127364 118772 128239
rect 119020 128204 119060 128239
rect 119116 128213 119156 130339
rect 119020 128155 119060 128164
rect 119115 128204 119157 128213
rect 119115 128164 119116 128204
rect 119156 128164 119157 128204
rect 119115 128155 119157 128164
rect 119212 128204 119252 130423
rect 119500 128876 119540 128885
rect 120364 128876 120404 128885
rect 119308 128836 119500 128876
rect 119308 128372 119348 128836
rect 119500 128827 119540 128836
rect 119788 128836 120364 128876
rect 119691 128708 119733 128717
rect 119691 128668 119692 128708
rect 119732 128668 119733 128708
rect 119691 128659 119733 128668
rect 119308 128323 119348 128332
rect 119596 128213 119636 128298
rect 119692 128297 119732 128659
rect 119788 128372 119828 128836
rect 120364 128827 120404 128836
rect 120172 128708 120212 128717
rect 119788 128323 119828 128332
rect 119884 128668 120172 128708
rect 119691 128288 119733 128297
rect 119691 128248 119692 128288
rect 119732 128248 119733 128288
rect 119691 128239 119733 128248
rect 119595 128204 119637 128213
rect 119252 128164 119348 128180
rect 118827 127952 118869 127961
rect 118827 127912 118828 127952
rect 118868 127912 118869 127952
rect 118827 127903 118869 127912
rect 118828 127818 118868 127903
rect 119116 127784 119156 128155
rect 119212 128140 119348 128164
rect 119595 128164 119596 128204
rect 119636 128164 119637 128204
rect 119595 128155 119637 128164
rect 119692 128204 119732 128239
rect 119692 128155 119732 128164
rect 119884 128204 119924 128668
rect 120172 128659 120212 128668
rect 120460 128213 120500 133363
rect 120652 133278 120692 133363
rect 121804 133244 121844 133253
rect 121804 132749 121844 133204
rect 124784 133076 125152 133085
rect 124824 133036 124866 133076
rect 124906 133036 124948 133076
rect 124988 133036 125030 133076
rect 125070 133036 125112 133076
rect 124784 133027 125152 133036
rect 120939 132740 120981 132749
rect 120939 132700 120940 132740
rect 120980 132700 120981 132740
rect 120939 132691 120981 132700
rect 121803 132740 121845 132749
rect 121803 132700 121804 132740
rect 121844 132700 121845 132740
rect 121803 132691 121845 132700
rect 120940 132606 120980 132691
rect 135724 132665 135764 160020
rect 139904 148196 140272 148205
rect 139944 148156 139986 148196
rect 140026 148156 140068 148196
rect 140108 148156 140150 148196
rect 140190 148156 140232 148196
rect 139904 148147 140272 148156
rect 138664 147440 139032 147449
rect 138704 147400 138746 147440
rect 138786 147400 138828 147440
rect 138868 147400 138910 147440
rect 138950 147400 138992 147440
rect 138664 147391 139032 147400
rect 139904 146684 140272 146693
rect 139944 146644 139986 146684
rect 140026 146644 140068 146684
rect 140108 146644 140150 146684
rect 140190 146644 140232 146684
rect 139904 146635 140272 146644
rect 138664 145928 139032 145937
rect 138704 145888 138746 145928
rect 138786 145888 138828 145928
rect 138868 145888 138910 145928
rect 138950 145888 138992 145928
rect 138664 145879 139032 145888
rect 139904 145172 140272 145181
rect 139944 145132 139986 145172
rect 140026 145132 140068 145172
rect 140108 145132 140150 145172
rect 140190 145132 140232 145172
rect 139904 145123 140272 145132
rect 138664 144416 139032 144425
rect 138704 144376 138746 144416
rect 138786 144376 138828 144416
rect 138868 144376 138910 144416
rect 138950 144376 138992 144416
rect 138664 144367 139032 144376
rect 139904 143660 140272 143669
rect 139944 143620 139986 143660
rect 140026 143620 140068 143660
rect 140108 143620 140150 143660
rect 140190 143620 140232 143660
rect 139904 143611 140272 143620
rect 138664 142904 139032 142913
rect 138704 142864 138746 142904
rect 138786 142864 138828 142904
rect 138868 142864 138910 142904
rect 138950 142864 138992 142904
rect 138664 142855 139032 142864
rect 139904 142148 140272 142157
rect 139944 142108 139986 142148
rect 140026 142108 140068 142148
rect 140108 142108 140150 142148
rect 140190 142108 140232 142148
rect 139904 142099 140272 142108
rect 138664 141392 139032 141401
rect 138704 141352 138746 141392
rect 138786 141352 138828 141392
rect 138868 141352 138910 141392
rect 138950 141352 138992 141392
rect 138664 141343 139032 141352
rect 139904 140636 140272 140645
rect 139944 140596 139986 140636
rect 140026 140596 140068 140636
rect 140108 140596 140150 140636
rect 140190 140596 140232 140636
rect 139904 140587 140272 140596
rect 138664 139880 139032 139889
rect 138704 139840 138746 139880
rect 138786 139840 138828 139880
rect 138868 139840 138910 139880
rect 138950 139840 138992 139880
rect 138664 139831 139032 139840
rect 139904 139124 140272 139133
rect 139944 139084 139986 139124
rect 140026 139084 140068 139124
rect 140108 139084 140150 139124
rect 140190 139084 140232 139124
rect 139904 139075 140272 139084
rect 138664 138368 139032 138377
rect 138704 138328 138746 138368
rect 138786 138328 138828 138368
rect 138868 138328 138910 138368
rect 138950 138328 138992 138368
rect 138664 138319 139032 138328
rect 139904 137612 140272 137621
rect 139944 137572 139986 137612
rect 140026 137572 140068 137612
rect 140108 137572 140150 137612
rect 140190 137572 140232 137612
rect 139904 137563 140272 137572
rect 138664 136856 139032 136865
rect 138704 136816 138746 136856
rect 138786 136816 138828 136856
rect 138868 136816 138910 136856
rect 138950 136816 138992 136856
rect 138664 136807 139032 136816
rect 139904 136100 140272 136109
rect 139944 136060 139986 136100
rect 140026 136060 140068 136100
rect 140108 136060 140150 136100
rect 140190 136060 140232 136100
rect 139904 136051 140272 136060
rect 138664 135344 139032 135353
rect 138704 135304 138746 135344
rect 138786 135304 138828 135344
rect 138868 135304 138910 135344
rect 138950 135304 138992 135344
rect 138664 135295 139032 135304
rect 139904 134588 140272 134597
rect 139944 134548 139986 134588
rect 140026 134548 140068 134588
rect 140108 134548 140150 134588
rect 140190 134548 140232 134588
rect 139904 134539 140272 134548
rect 151660 134093 151700 160020
rect 151659 134084 151701 134093
rect 151659 134044 151660 134084
rect 151700 134044 151701 134084
rect 151659 134035 151701 134044
rect 138664 133832 139032 133841
rect 138704 133792 138746 133832
rect 138786 133792 138828 133832
rect 138868 133792 138910 133832
rect 138950 133792 138992 133832
rect 138664 133783 139032 133792
rect 139904 133076 140272 133085
rect 139944 133036 139986 133076
rect 140026 133036 140068 133076
rect 140108 133036 140150 133076
rect 140190 133036 140232 133076
rect 139904 133027 140272 133036
rect 135723 132656 135765 132665
rect 135723 132616 135724 132656
rect 135764 132616 135765 132656
rect 135723 132607 135765 132616
rect 123544 132320 123912 132329
rect 123584 132280 123626 132320
rect 123666 132280 123708 132320
rect 123748 132280 123790 132320
rect 123830 132280 123872 132320
rect 123544 132271 123912 132280
rect 138664 132320 139032 132329
rect 138704 132280 138746 132320
rect 138786 132280 138828 132320
rect 138868 132280 138910 132320
rect 138950 132280 138992 132320
rect 138664 132271 139032 132280
rect 124784 131564 125152 131573
rect 124824 131524 124866 131564
rect 124906 131524 124948 131564
rect 124988 131524 125030 131564
rect 125070 131524 125112 131564
rect 124784 131515 125152 131524
rect 139904 131564 140272 131573
rect 139944 131524 139986 131564
rect 140026 131524 140068 131564
rect 140108 131524 140150 131564
rect 140190 131524 140232 131564
rect 139904 131515 140272 131524
rect 123544 130808 123912 130817
rect 123584 130768 123626 130808
rect 123666 130768 123708 130808
rect 123748 130768 123790 130808
rect 123830 130768 123872 130808
rect 123544 130759 123912 130768
rect 138664 130808 139032 130817
rect 138704 130768 138746 130808
rect 138786 130768 138828 130808
rect 138868 130768 138910 130808
rect 138950 130768 138992 130808
rect 138664 130759 139032 130768
rect 124784 130052 125152 130061
rect 124824 130012 124866 130052
rect 124906 130012 124948 130052
rect 124988 130012 125030 130052
rect 125070 130012 125112 130052
rect 124784 130003 125152 130012
rect 139904 130052 140272 130061
rect 139944 130012 139986 130052
rect 140026 130012 140068 130052
rect 140108 130012 140150 130052
rect 140190 130012 140232 130052
rect 139904 130003 140272 130012
rect 123544 129296 123912 129305
rect 123584 129256 123626 129296
rect 123666 129256 123708 129296
rect 123748 129256 123790 129296
rect 123830 129256 123872 129296
rect 123544 129247 123912 129256
rect 138664 129296 139032 129305
rect 138704 129256 138746 129296
rect 138786 129256 138828 129296
rect 138868 129256 138910 129296
rect 138950 129256 138992 129296
rect 138664 129247 139032 129256
rect 121228 129044 121268 129053
rect 121132 129004 121228 129044
rect 121036 128708 121076 128717
rect 120748 128668 121036 128708
rect 120748 128288 120788 128668
rect 121036 128659 121076 128668
rect 120748 128239 120788 128248
rect 119884 128155 119924 128164
rect 120459 128204 120501 128213
rect 120459 128164 120460 128204
rect 120500 128164 120501 128204
rect 120459 128155 120501 128164
rect 121132 128204 121172 129004
rect 121228 128995 121268 129004
rect 121995 128876 122037 128885
rect 121995 128836 121996 128876
rect 122036 128836 122037 128876
rect 121995 128827 122037 128836
rect 123147 128876 123189 128885
rect 123147 128836 123148 128876
rect 123188 128836 123189 128876
rect 123147 128827 123189 128836
rect 121996 128742 122036 128827
rect 121899 128708 121941 128717
rect 121899 128668 121900 128708
rect 121940 128668 121941 128708
rect 121899 128659 121941 128668
rect 121900 128574 121940 128659
rect 123148 128372 123188 128827
rect 124784 128540 125152 128549
rect 124824 128500 124866 128540
rect 124906 128500 124948 128540
rect 124988 128500 125030 128540
rect 125070 128500 125112 128540
rect 124784 128491 125152 128500
rect 139904 128540 140272 128549
rect 139944 128500 139986 128540
rect 140026 128500 140068 128540
rect 140108 128500 140150 128540
rect 140190 128500 140232 128540
rect 139904 128491 140272 128500
rect 123148 128323 123188 128332
rect 121996 128213 122036 128298
rect 121132 128155 121172 128164
rect 121995 128204 122037 128213
rect 121995 128164 121996 128204
rect 122036 128164 122037 128204
rect 121995 128155 122037 128164
rect 119211 127952 119253 127961
rect 119211 127912 119212 127952
rect 119252 127912 119253 127952
rect 119211 127903 119253 127912
rect 118924 127744 119156 127784
rect 118828 127364 118868 127373
rect 118732 127324 118828 127364
rect 118828 127315 118868 127324
rect 118924 127364 118964 127744
rect 118924 127315 118964 127324
rect 119020 127364 119060 127373
rect 119020 127196 119060 127324
rect 118636 127156 119060 127196
rect 109664 127028 110032 127037
rect 109704 126988 109746 127028
rect 109786 126988 109828 127028
rect 109868 126988 109910 127028
rect 109950 126988 109992 127028
rect 109664 126979 110032 126988
rect 108424 126272 108792 126281
rect 108464 126232 108506 126272
rect 108546 126232 108588 126272
rect 108628 126232 108670 126272
rect 108710 126232 108752 126272
rect 108424 126223 108792 126232
rect 109664 125516 110032 125525
rect 109704 125476 109746 125516
rect 109786 125476 109828 125516
rect 109868 125476 109910 125516
rect 109950 125476 109992 125516
rect 109664 125467 110032 125476
rect 119020 125357 119060 127156
rect 119116 127196 119156 127205
rect 119116 125852 119156 127156
rect 119212 125877 119252 127903
rect 119212 125828 119252 125837
rect 119116 125803 119156 125812
rect 119116 125684 119156 125693
rect 119308 125684 119348 128140
rect 119979 126692 120021 126701
rect 119979 126652 119980 126692
rect 120020 126652 120021 126692
rect 119979 126643 120021 126652
rect 119156 125644 119348 125684
rect 119404 125768 119444 125777
rect 119116 125635 119156 125644
rect 119019 125348 119061 125357
rect 119019 125308 119020 125348
rect 119060 125308 119061 125348
rect 119019 125299 119061 125308
rect 108424 124760 108792 124769
rect 108464 124720 108506 124760
rect 108546 124720 108588 124760
rect 108628 124720 108670 124760
rect 108710 124720 108752 124760
rect 108424 124711 108792 124720
rect 109664 124004 110032 124013
rect 109704 123964 109746 124004
rect 109786 123964 109828 124004
rect 109868 123964 109910 124004
rect 109950 123964 109992 124004
rect 109664 123955 110032 123964
rect 119212 123752 119252 123761
rect 119404 123752 119444 125728
rect 119252 123712 119444 123752
rect 119212 123703 119252 123712
rect 119596 123668 119636 123677
rect 108424 123248 108792 123257
rect 108464 123208 108506 123248
rect 108546 123208 108588 123248
rect 108628 123208 108670 123248
rect 108710 123208 108752 123248
rect 108424 123199 108792 123208
rect 119596 122996 119636 123628
rect 119692 122996 119732 123005
rect 119596 122956 119692 122996
rect 119692 122947 119732 122956
rect 109664 122492 110032 122501
rect 109704 122452 109746 122492
rect 109786 122452 109828 122492
rect 109868 122452 109910 122492
rect 109950 122452 109992 122492
rect 109664 122443 110032 122452
rect 108424 121736 108792 121745
rect 108464 121696 108506 121736
rect 108546 121696 108588 121736
rect 108628 121696 108670 121736
rect 108710 121696 108752 121736
rect 108424 121687 108792 121696
rect 109664 120980 110032 120989
rect 109704 120940 109746 120980
rect 109786 120940 109828 120980
rect 109868 120940 109910 120980
rect 109950 120940 109992 120980
rect 109664 120931 110032 120940
rect 108424 120224 108792 120233
rect 108464 120184 108506 120224
rect 108546 120184 108588 120224
rect 108628 120184 108670 120224
rect 108710 120184 108752 120224
rect 108424 120175 108792 120184
rect 109664 119468 110032 119477
rect 109704 119428 109746 119468
rect 109786 119428 109828 119468
rect 109868 119428 109910 119468
rect 109950 119428 109992 119468
rect 109664 119419 110032 119428
rect 108424 118712 108792 118721
rect 108464 118672 108506 118712
rect 108546 118672 108588 118712
rect 108628 118672 108670 118712
rect 108710 118672 108752 118712
rect 108424 118663 108792 118672
rect 109664 117956 110032 117965
rect 109704 117916 109746 117956
rect 109786 117916 109828 117956
rect 109868 117916 109910 117956
rect 109950 117916 109992 117956
rect 109664 117907 110032 117916
rect 108424 117200 108792 117209
rect 108464 117160 108506 117200
rect 108546 117160 108588 117200
rect 108628 117160 108670 117200
rect 108710 117160 108752 117200
rect 108424 117151 108792 117160
rect 109664 116444 110032 116453
rect 109704 116404 109746 116444
rect 109786 116404 109828 116444
rect 109868 116404 109910 116444
rect 109950 116404 109992 116444
rect 109664 116395 110032 116404
rect 108424 115688 108792 115697
rect 108464 115648 108506 115688
rect 108546 115648 108588 115688
rect 108628 115648 108670 115688
rect 108710 115648 108752 115688
rect 108424 115639 108792 115648
rect 109664 114932 110032 114941
rect 109704 114892 109746 114932
rect 109786 114892 109828 114932
rect 109868 114892 109910 114932
rect 109950 114892 109992 114932
rect 109664 114883 110032 114892
rect 108424 114176 108792 114185
rect 108464 114136 108506 114176
rect 108546 114136 108588 114176
rect 108628 114136 108670 114176
rect 108710 114136 108752 114176
rect 108424 114127 108792 114136
rect 109664 113420 110032 113429
rect 109704 113380 109746 113420
rect 109786 113380 109828 113420
rect 109868 113380 109910 113420
rect 109950 113380 109992 113420
rect 109664 113371 110032 113380
rect 108424 112664 108792 112673
rect 108464 112624 108506 112664
rect 108546 112624 108588 112664
rect 108628 112624 108670 112664
rect 108710 112624 108752 112664
rect 108424 112615 108792 112624
rect 109664 111908 110032 111917
rect 109704 111868 109746 111908
rect 109786 111868 109828 111908
rect 109868 111868 109910 111908
rect 109950 111868 109992 111908
rect 109664 111859 110032 111868
rect 108424 111152 108792 111161
rect 108464 111112 108506 111152
rect 108546 111112 108588 111152
rect 108628 111112 108670 111152
rect 108710 111112 108752 111152
rect 108424 111103 108792 111112
rect 109664 110396 110032 110405
rect 109704 110356 109746 110396
rect 109786 110356 109828 110396
rect 109868 110356 109910 110396
rect 109950 110356 109992 110396
rect 109664 110347 110032 110356
rect 108424 109640 108792 109649
rect 108464 109600 108506 109640
rect 108546 109600 108588 109640
rect 108628 109600 108670 109640
rect 108710 109600 108752 109640
rect 108424 109591 108792 109600
rect 109664 108884 110032 108893
rect 109704 108844 109746 108884
rect 109786 108844 109828 108884
rect 109868 108844 109910 108884
rect 109950 108844 109992 108884
rect 109664 108835 110032 108844
rect 108424 108128 108792 108137
rect 108464 108088 108506 108128
rect 108546 108088 108588 108128
rect 108628 108088 108670 108128
rect 108710 108088 108752 108128
rect 108424 108079 108792 108088
rect 109664 107372 110032 107381
rect 109704 107332 109746 107372
rect 109786 107332 109828 107372
rect 109868 107332 109910 107372
rect 109950 107332 109992 107372
rect 109664 107323 110032 107332
rect 108424 106616 108792 106625
rect 108464 106576 108506 106616
rect 108546 106576 108588 106616
rect 108628 106576 108670 106616
rect 108710 106576 108752 106616
rect 108424 106567 108792 106576
rect 109664 105860 110032 105869
rect 109704 105820 109746 105860
rect 109786 105820 109828 105860
rect 109868 105820 109910 105860
rect 109950 105820 109992 105860
rect 109664 105811 110032 105820
rect 108424 105104 108792 105113
rect 108464 105064 108506 105104
rect 108546 105064 108588 105104
rect 108628 105064 108670 105104
rect 108710 105064 108752 105104
rect 108424 105055 108792 105064
rect 109664 104348 110032 104357
rect 109704 104308 109746 104348
rect 109786 104308 109828 104348
rect 109868 104308 109910 104348
rect 109950 104308 109992 104348
rect 109664 104299 110032 104308
rect 108424 103592 108792 103601
rect 108464 103552 108506 103592
rect 108546 103552 108588 103592
rect 108628 103552 108670 103592
rect 108710 103552 108752 103592
rect 108424 103543 108792 103552
rect 109664 102836 110032 102845
rect 109704 102796 109746 102836
rect 109786 102796 109828 102836
rect 109868 102796 109910 102836
rect 109950 102796 109992 102836
rect 109664 102787 110032 102796
rect 108424 102080 108792 102089
rect 108464 102040 108506 102080
rect 108546 102040 108588 102080
rect 108628 102040 108670 102080
rect 108710 102040 108752 102080
rect 108424 102031 108792 102040
rect 109664 101324 110032 101333
rect 109704 101284 109746 101324
rect 109786 101284 109828 101324
rect 109868 101284 109910 101324
rect 109950 101284 109992 101324
rect 109664 101275 110032 101284
rect 108424 100568 108792 100577
rect 108464 100528 108506 100568
rect 108546 100528 108588 100568
rect 108628 100528 108670 100568
rect 108710 100528 108752 100568
rect 108424 100519 108792 100528
rect 109664 99812 110032 99821
rect 109704 99772 109746 99812
rect 109786 99772 109828 99812
rect 109868 99772 109910 99812
rect 109950 99772 109992 99812
rect 109664 99763 110032 99772
rect 108424 99056 108792 99065
rect 108464 99016 108506 99056
rect 108546 99016 108588 99056
rect 108628 99016 108670 99056
rect 108710 99016 108752 99056
rect 108424 99007 108792 99016
rect 109664 98300 110032 98309
rect 109704 98260 109746 98300
rect 109786 98260 109828 98300
rect 109868 98260 109910 98300
rect 109950 98260 109992 98300
rect 109664 98251 110032 98260
rect 108424 97544 108792 97553
rect 108464 97504 108506 97544
rect 108546 97504 108588 97544
rect 108628 97504 108670 97544
rect 108710 97504 108752 97544
rect 108424 97495 108792 97504
rect 109664 96788 110032 96797
rect 109704 96748 109746 96788
rect 109786 96748 109828 96788
rect 109868 96748 109910 96788
rect 109950 96748 109992 96788
rect 109664 96739 110032 96748
rect 108424 96032 108792 96041
rect 108464 95992 108506 96032
rect 108546 95992 108588 96032
rect 108628 95992 108670 96032
rect 108710 95992 108752 96032
rect 108424 95983 108792 95992
rect 104332 95815 104372 95824
rect 109664 95276 110032 95285
rect 109704 95236 109746 95276
rect 109786 95236 109828 95276
rect 109868 95236 109910 95276
rect 109950 95236 109992 95276
rect 109664 95227 110032 95236
rect 108424 94520 108792 94529
rect 108464 94480 108506 94520
rect 108546 94480 108588 94520
rect 108628 94480 108670 94520
rect 108710 94480 108752 94520
rect 108424 94471 108792 94480
rect 109664 93764 110032 93773
rect 109704 93724 109746 93764
rect 109786 93724 109828 93764
rect 109868 93724 109910 93764
rect 109950 93724 109992 93764
rect 109664 93715 110032 93724
rect 108424 93008 108792 93017
rect 108464 92968 108506 93008
rect 108546 92968 108588 93008
rect 108628 92968 108670 93008
rect 108710 92968 108752 93008
rect 108424 92959 108792 92968
rect 109664 92252 110032 92261
rect 109704 92212 109746 92252
rect 109786 92212 109828 92252
rect 109868 92212 109910 92252
rect 109950 92212 109992 92252
rect 109664 92203 110032 92212
rect 108424 91496 108792 91505
rect 108464 91456 108506 91496
rect 108546 91456 108588 91496
rect 108628 91456 108670 91496
rect 108710 91456 108752 91496
rect 108424 91447 108792 91456
rect 109664 90740 110032 90749
rect 109704 90700 109746 90740
rect 109786 90700 109828 90740
rect 109868 90700 109910 90740
rect 109950 90700 109992 90740
rect 109664 90691 110032 90700
rect 108424 89984 108792 89993
rect 108464 89944 108506 89984
rect 108546 89944 108588 89984
rect 108628 89944 108670 89984
rect 108710 89944 108752 89984
rect 108424 89935 108792 89944
rect 109664 89228 110032 89237
rect 109704 89188 109746 89228
rect 109786 89188 109828 89228
rect 109868 89188 109910 89228
rect 109950 89188 109992 89228
rect 109664 89179 110032 89188
rect 108424 88472 108792 88481
rect 108464 88432 108506 88472
rect 108546 88432 108588 88472
rect 108628 88432 108670 88472
rect 108710 88432 108752 88472
rect 108424 88423 108792 88432
rect 109664 87716 110032 87725
rect 109704 87676 109746 87716
rect 109786 87676 109828 87716
rect 109868 87676 109910 87716
rect 109950 87676 109992 87716
rect 109664 87667 110032 87676
rect 108424 86960 108792 86969
rect 108464 86920 108506 86960
rect 108546 86920 108588 86960
rect 108628 86920 108670 86960
rect 108710 86920 108752 86960
rect 108424 86911 108792 86920
rect 109664 86204 110032 86213
rect 109704 86164 109746 86204
rect 109786 86164 109828 86204
rect 109868 86164 109910 86204
rect 109950 86164 109992 86204
rect 109664 86155 110032 86164
rect 108424 85448 108792 85457
rect 108464 85408 108506 85448
rect 108546 85408 108588 85448
rect 108628 85408 108670 85448
rect 108710 85408 108752 85448
rect 108424 85399 108792 85408
rect 109664 84692 110032 84701
rect 109704 84652 109746 84692
rect 109786 84652 109828 84692
rect 109868 84652 109910 84692
rect 109950 84652 109992 84692
rect 109664 84643 110032 84652
rect 108424 83936 108792 83945
rect 108464 83896 108506 83936
rect 108546 83896 108588 83936
rect 108628 83896 108670 83936
rect 108710 83896 108752 83936
rect 108424 83887 108792 83896
rect 109664 83180 110032 83189
rect 109704 83140 109746 83180
rect 109786 83140 109828 83180
rect 109868 83140 109910 83180
rect 109950 83140 109992 83180
rect 109664 83131 110032 83140
rect 108424 82424 108792 82433
rect 108464 82384 108506 82424
rect 108546 82384 108588 82424
rect 108628 82384 108670 82424
rect 108710 82384 108752 82424
rect 108424 82375 108792 82384
rect 109664 81668 110032 81677
rect 109704 81628 109746 81668
rect 109786 81628 109828 81668
rect 109868 81628 109910 81668
rect 109950 81628 109992 81668
rect 109664 81619 110032 81628
rect 108424 80912 108792 80921
rect 108464 80872 108506 80912
rect 108546 80872 108588 80912
rect 108628 80872 108670 80912
rect 108710 80872 108752 80912
rect 108424 80863 108792 80872
rect 109664 80156 110032 80165
rect 109704 80116 109746 80156
rect 109786 80116 109828 80156
rect 109868 80116 109910 80156
rect 109950 80116 109992 80156
rect 109664 80107 110032 80116
rect 108424 79400 108792 79409
rect 108464 79360 108506 79400
rect 108546 79360 108588 79400
rect 108628 79360 108670 79400
rect 108710 79360 108752 79400
rect 108424 79351 108792 79360
rect 109664 78644 110032 78653
rect 109704 78604 109746 78644
rect 109786 78604 109828 78644
rect 109868 78604 109910 78644
rect 109950 78604 109992 78644
rect 109664 78595 110032 78604
rect 108424 77888 108792 77897
rect 108464 77848 108506 77888
rect 108546 77848 108588 77888
rect 108628 77848 108670 77888
rect 108710 77848 108752 77888
rect 108424 77839 108792 77848
rect 109664 77132 110032 77141
rect 109704 77092 109746 77132
rect 109786 77092 109828 77132
rect 109868 77092 109910 77132
rect 109950 77092 109992 77132
rect 109664 77083 110032 77092
rect 108424 76376 108792 76385
rect 108464 76336 108506 76376
rect 108546 76336 108588 76376
rect 108628 76336 108670 76376
rect 108710 76336 108752 76376
rect 108424 76327 108792 76336
rect 109664 75620 110032 75629
rect 109704 75580 109746 75620
rect 109786 75580 109828 75620
rect 109868 75580 109910 75620
rect 109950 75580 109992 75620
rect 109664 75571 110032 75580
rect 119980 64364 120020 126643
rect 120460 123668 120500 128155
rect 123148 127952 123188 127961
rect 121035 125348 121077 125357
rect 121035 125308 121036 125348
rect 121076 125308 121077 125348
rect 121035 125299 121077 125308
rect 121036 125214 121076 125299
rect 121132 125180 121172 125189
rect 121516 125180 121556 125189
rect 121172 125140 121516 125180
rect 121132 125131 121172 125140
rect 121516 125131 121556 125140
rect 122188 125180 122228 125189
rect 121612 123836 121652 123845
rect 122188 123836 122228 125140
rect 121652 123796 122228 123836
rect 121612 123787 121652 123796
rect 120460 123619 120500 123628
rect 121612 123416 121652 123425
rect 121612 103769 121652 123376
rect 123148 119645 123188 127912
rect 123544 127784 123912 127793
rect 123584 127744 123626 127784
rect 123666 127744 123708 127784
rect 123748 127744 123790 127784
rect 123830 127744 123872 127784
rect 123544 127735 123912 127744
rect 138664 127784 139032 127793
rect 138704 127744 138746 127784
rect 138786 127744 138828 127784
rect 138868 127744 138910 127784
rect 138950 127744 138992 127784
rect 138664 127735 139032 127744
rect 124784 127028 125152 127037
rect 124824 126988 124866 127028
rect 124906 126988 124948 127028
rect 124988 126988 125030 127028
rect 125070 126988 125112 127028
rect 124784 126979 125152 126988
rect 139904 127028 140272 127037
rect 139944 126988 139986 127028
rect 140026 126988 140068 127028
rect 140108 126988 140150 127028
rect 140190 126988 140232 127028
rect 139904 126979 140272 126988
rect 123544 126272 123912 126281
rect 123584 126232 123626 126272
rect 123666 126232 123708 126272
rect 123748 126232 123790 126272
rect 123830 126232 123872 126272
rect 123544 126223 123912 126232
rect 138664 126272 139032 126281
rect 138704 126232 138746 126272
rect 138786 126232 138828 126272
rect 138868 126232 138910 126272
rect 138950 126232 138992 126272
rect 138664 126223 139032 126232
rect 124784 125516 125152 125525
rect 124824 125476 124866 125516
rect 124906 125476 124948 125516
rect 124988 125476 125030 125516
rect 125070 125476 125112 125516
rect 124784 125467 125152 125476
rect 139904 125516 140272 125525
rect 139944 125476 139986 125516
rect 140026 125476 140068 125516
rect 140108 125476 140150 125516
rect 140190 125476 140232 125516
rect 139904 125467 140272 125476
rect 123544 124760 123912 124769
rect 123584 124720 123626 124760
rect 123666 124720 123708 124760
rect 123748 124720 123790 124760
rect 123830 124720 123872 124760
rect 123544 124711 123912 124720
rect 138664 124760 139032 124769
rect 138704 124720 138746 124760
rect 138786 124720 138828 124760
rect 138868 124720 138910 124760
rect 138950 124720 138992 124760
rect 138664 124711 139032 124720
rect 124784 124004 125152 124013
rect 124824 123964 124866 124004
rect 124906 123964 124948 124004
rect 124988 123964 125030 124004
rect 125070 123964 125112 124004
rect 124784 123955 125152 123964
rect 139904 124004 140272 124013
rect 139944 123964 139986 124004
rect 140026 123964 140068 124004
rect 140108 123964 140150 124004
rect 140190 123964 140232 124004
rect 139904 123955 140272 123964
rect 123544 123248 123912 123257
rect 123584 123208 123626 123248
rect 123666 123208 123708 123248
rect 123748 123208 123790 123248
rect 123830 123208 123872 123248
rect 123544 123199 123912 123208
rect 138664 123248 139032 123257
rect 138704 123208 138746 123248
rect 138786 123208 138828 123248
rect 138868 123208 138910 123248
rect 138950 123208 138992 123248
rect 138664 123199 139032 123208
rect 124784 122492 125152 122501
rect 124824 122452 124866 122492
rect 124906 122452 124948 122492
rect 124988 122452 125030 122492
rect 125070 122452 125112 122492
rect 124784 122443 125152 122452
rect 139904 122492 140272 122501
rect 139944 122452 139986 122492
rect 140026 122452 140068 122492
rect 140108 122452 140150 122492
rect 140190 122452 140232 122492
rect 139904 122443 140272 122452
rect 123544 121736 123912 121745
rect 123584 121696 123626 121736
rect 123666 121696 123708 121736
rect 123748 121696 123790 121736
rect 123830 121696 123872 121736
rect 123544 121687 123912 121696
rect 138664 121736 139032 121745
rect 138704 121696 138746 121736
rect 138786 121696 138828 121736
rect 138868 121696 138910 121736
rect 138950 121696 138992 121736
rect 138664 121687 139032 121696
rect 124784 120980 125152 120989
rect 124824 120940 124866 120980
rect 124906 120940 124948 120980
rect 124988 120940 125030 120980
rect 125070 120940 125112 120980
rect 124784 120931 125152 120940
rect 139904 120980 140272 120989
rect 139944 120940 139986 120980
rect 140026 120940 140068 120980
rect 140108 120940 140150 120980
rect 140190 120940 140232 120980
rect 139904 120931 140272 120940
rect 123544 120224 123912 120233
rect 123584 120184 123626 120224
rect 123666 120184 123708 120224
rect 123748 120184 123790 120224
rect 123830 120184 123872 120224
rect 123544 120175 123912 120184
rect 138664 120224 139032 120233
rect 138704 120184 138746 120224
rect 138786 120184 138828 120224
rect 138868 120184 138910 120224
rect 138950 120184 138992 120224
rect 138664 120175 139032 120184
rect 123147 119636 123189 119645
rect 123147 119596 123148 119636
rect 123188 119596 123189 119636
rect 123147 119587 123189 119596
rect 124784 119468 125152 119477
rect 124824 119428 124866 119468
rect 124906 119428 124948 119468
rect 124988 119428 125030 119468
rect 125070 119428 125112 119468
rect 124784 119419 125152 119428
rect 139904 119468 140272 119477
rect 139944 119428 139986 119468
rect 140026 119428 140068 119468
rect 140108 119428 140150 119468
rect 140190 119428 140232 119468
rect 139904 119419 140272 119428
rect 123544 118712 123912 118721
rect 123584 118672 123626 118712
rect 123666 118672 123708 118712
rect 123748 118672 123790 118712
rect 123830 118672 123872 118712
rect 123544 118663 123912 118672
rect 138664 118712 139032 118721
rect 138704 118672 138746 118712
rect 138786 118672 138828 118712
rect 138868 118672 138910 118712
rect 138950 118672 138992 118712
rect 138664 118663 139032 118672
rect 124784 117956 125152 117965
rect 124824 117916 124866 117956
rect 124906 117916 124948 117956
rect 124988 117916 125030 117956
rect 125070 117916 125112 117956
rect 124784 117907 125152 117916
rect 139904 117956 140272 117965
rect 139944 117916 139986 117956
rect 140026 117916 140068 117956
rect 140108 117916 140150 117956
rect 140190 117916 140232 117956
rect 139904 117907 140272 117916
rect 123544 117200 123912 117209
rect 123584 117160 123626 117200
rect 123666 117160 123708 117200
rect 123748 117160 123790 117200
rect 123830 117160 123872 117200
rect 123544 117151 123912 117160
rect 138664 117200 139032 117209
rect 138704 117160 138746 117200
rect 138786 117160 138828 117200
rect 138868 117160 138910 117200
rect 138950 117160 138992 117200
rect 138664 117151 139032 117160
rect 124784 116444 125152 116453
rect 124824 116404 124866 116444
rect 124906 116404 124948 116444
rect 124988 116404 125030 116444
rect 125070 116404 125112 116444
rect 124784 116395 125152 116404
rect 139904 116444 140272 116453
rect 139944 116404 139986 116444
rect 140026 116404 140068 116444
rect 140108 116404 140150 116444
rect 140190 116404 140232 116444
rect 139904 116395 140272 116404
rect 123544 115688 123912 115697
rect 123584 115648 123626 115688
rect 123666 115648 123708 115688
rect 123748 115648 123790 115688
rect 123830 115648 123872 115688
rect 123544 115639 123912 115648
rect 138664 115688 139032 115697
rect 138704 115648 138746 115688
rect 138786 115648 138828 115688
rect 138868 115648 138910 115688
rect 138950 115648 138992 115688
rect 138664 115639 139032 115648
rect 124784 114932 125152 114941
rect 124824 114892 124866 114932
rect 124906 114892 124948 114932
rect 124988 114892 125030 114932
rect 125070 114892 125112 114932
rect 124784 114883 125152 114892
rect 139904 114932 140272 114941
rect 139944 114892 139986 114932
rect 140026 114892 140068 114932
rect 140108 114892 140150 114932
rect 140190 114892 140232 114932
rect 139904 114883 140272 114892
rect 123544 114176 123912 114185
rect 123584 114136 123626 114176
rect 123666 114136 123708 114176
rect 123748 114136 123790 114176
rect 123830 114136 123872 114176
rect 123544 114127 123912 114136
rect 138664 114176 139032 114185
rect 138704 114136 138746 114176
rect 138786 114136 138828 114176
rect 138868 114136 138910 114176
rect 138950 114136 138992 114176
rect 138664 114127 139032 114136
rect 124784 113420 125152 113429
rect 124824 113380 124866 113420
rect 124906 113380 124948 113420
rect 124988 113380 125030 113420
rect 125070 113380 125112 113420
rect 124784 113371 125152 113380
rect 139904 113420 140272 113429
rect 139944 113380 139986 113420
rect 140026 113380 140068 113420
rect 140108 113380 140150 113420
rect 140190 113380 140232 113420
rect 139904 113371 140272 113380
rect 123544 112664 123912 112673
rect 123584 112624 123626 112664
rect 123666 112624 123708 112664
rect 123748 112624 123790 112664
rect 123830 112624 123872 112664
rect 123544 112615 123912 112624
rect 138664 112664 139032 112673
rect 138704 112624 138746 112664
rect 138786 112624 138828 112664
rect 138868 112624 138910 112664
rect 138950 112624 138992 112664
rect 138664 112615 139032 112624
rect 124784 111908 125152 111917
rect 124824 111868 124866 111908
rect 124906 111868 124948 111908
rect 124988 111868 125030 111908
rect 125070 111868 125112 111908
rect 124784 111859 125152 111868
rect 139904 111908 140272 111917
rect 139944 111868 139986 111908
rect 140026 111868 140068 111908
rect 140108 111868 140150 111908
rect 140190 111868 140232 111908
rect 139904 111859 140272 111868
rect 123544 111152 123912 111161
rect 123584 111112 123626 111152
rect 123666 111112 123708 111152
rect 123748 111112 123790 111152
rect 123830 111112 123872 111152
rect 123544 111103 123912 111112
rect 138664 111152 139032 111161
rect 138704 111112 138746 111152
rect 138786 111112 138828 111152
rect 138868 111112 138910 111152
rect 138950 111112 138992 111152
rect 138664 111103 139032 111112
rect 124784 110396 125152 110405
rect 124824 110356 124866 110396
rect 124906 110356 124948 110396
rect 124988 110356 125030 110396
rect 125070 110356 125112 110396
rect 124784 110347 125152 110356
rect 139904 110396 140272 110405
rect 139944 110356 139986 110396
rect 140026 110356 140068 110396
rect 140108 110356 140150 110396
rect 140190 110356 140232 110396
rect 139904 110347 140272 110356
rect 123544 109640 123912 109649
rect 123584 109600 123626 109640
rect 123666 109600 123708 109640
rect 123748 109600 123790 109640
rect 123830 109600 123872 109640
rect 123544 109591 123912 109600
rect 138664 109640 139032 109649
rect 138704 109600 138746 109640
rect 138786 109600 138828 109640
rect 138868 109600 138910 109640
rect 138950 109600 138992 109640
rect 138664 109591 139032 109600
rect 124784 108884 125152 108893
rect 124824 108844 124866 108884
rect 124906 108844 124948 108884
rect 124988 108844 125030 108884
rect 125070 108844 125112 108884
rect 124784 108835 125152 108844
rect 139904 108884 140272 108893
rect 139944 108844 139986 108884
rect 140026 108844 140068 108884
rect 140108 108844 140150 108884
rect 140190 108844 140232 108884
rect 139904 108835 140272 108844
rect 123544 108128 123912 108137
rect 123584 108088 123626 108128
rect 123666 108088 123708 108128
rect 123748 108088 123790 108128
rect 123830 108088 123872 108128
rect 123544 108079 123912 108088
rect 138664 108128 139032 108137
rect 138704 108088 138746 108128
rect 138786 108088 138828 108128
rect 138868 108088 138910 108128
rect 138950 108088 138992 108128
rect 138664 108079 139032 108088
rect 124784 107372 125152 107381
rect 124824 107332 124866 107372
rect 124906 107332 124948 107372
rect 124988 107332 125030 107372
rect 125070 107332 125112 107372
rect 124784 107323 125152 107332
rect 139904 107372 140272 107381
rect 139944 107332 139986 107372
rect 140026 107332 140068 107372
rect 140108 107332 140150 107372
rect 140190 107332 140232 107372
rect 139904 107323 140272 107332
rect 123544 106616 123912 106625
rect 123584 106576 123626 106616
rect 123666 106576 123708 106616
rect 123748 106576 123790 106616
rect 123830 106576 123872 106616
rect 123544 106567 123912 106576
rect 138664 106616 139032 106625
rect 138704 106576 138746 106616
rect 138786 106576 138828 106616
rect 138868 106576 138910 106616
rect 138950 106576 138992 106616
rect 138664 106567 139032 106576
rect 124784 105860 125152 105869
rect 124824 105820 124866 105860
rect 124906 105820 124948 105860
rect 124988 105820 125030 105860
rect 125070 105820 125112 105860
rect 124784 105811 125152 105820
rect 139904 105860 140272 105869
rect 139944 105820 139986 105860
rect 140026 105820 140068 105860
rect 140108 105820 140150 105860
rect 140190 105820 140232 105860
rect 139904 105811 140272 105820
rect 123544 105104 123912 105113
rect 123584 105064 123626 105104
rect 123666 105064 123708 105104
rect 123748 105064 123790 105104
rect 123830 105064 123872 105104
rect 123544 105055 123912 105064
rect 138664 105104 139032 105113
rect 138704 105064 138746 105104
rect 138786 105064 138828 105104
rect 138868 105064 138910 105104
rect 138950 105064 138992 105104
rect 138664 105055 139032 105064
rect 124784 104348 125152 104357
rect 124824 104308 124866 104348
rect 124906 104308 124948 104348
rect 124988 104308 125030 104348
rect 125070 104308 125112 104348
rect 124784 104299 125152 104308
rect 139904 104348 140272 104357
rect 139944 104308 139986 104348
rect 140026 104308 140068 104348
rect 140108 104308 140150 104348
rect 140190 104308 140232 104348
rect 139904 104299 140272 104308
rect 121611 103760 121653 103769
rect 121611 103720 121612 103760
rect 121652 103720 121653 103760
rect 121611 103711 121653 103720
rect 123544 103592 123912 103601
rect 123584 103552 123626 103592
rect 123666 103552 123708 103592
rect 123748 103552 123790 103592
rect 123830 103552 123872 103592
rect 123544 103543 123912 103552
rect 138664 103592 139032 103601
rect 138704 103552 138746 103592
rect 138786 103552 138828 103592
rect 138868 103552 138910 103592
rect 138950 103552 138992 103592
rect 138664 103543 139032 103552
rect 124784 102836 125152 102845
rect 124824 102796 124866 102836
rect 124906 102796 124948 102836
rect 124988 102796 125030 102836
rect 125070 102796 125112 102836
rect 124784 102787 125152 102796
rect 139904 102836 140272 102845
rect 139944 102796 139986 102836
rect 140026 102796 140068 102836
rect 140108 102796 140150 102836
rect 140190 102796 140232 102836
rect 139904 102787 140272 102796
rect 123544 102080 123912 102089
rect 123584 102040 123626 102080
rect 123666 102040 123708 102080
rect 123748 102040 123790 102080
rect 123830 102040 123872 102080
rect 123544 102031 123912 102040
rect 138664 102080 139032 102089
rect 138704 102040 138746 102080
rect 138786 102040 138828 102080
rect 138868 102040 138910 102080
rect 138950 102040 138992 102080
rect 138664 102031 139032 102040
rect 124784 101324 125152 101333
rect 124824 101284 124866 101324
rect 124906 101284 124948 101324
rect 124988 101284 125030 101324
rect 125070 101284 125112 101324
rect 124784 101275 125152 101284
rect 139904 101324 140272 101333
rect 139944 101284 139986 101324
rect 140026 101284 140068 101324
rect 140108 101284 140150 101324
rect 140190 101284 140232 101324
rect 139904 101275 140272 101284
rect 123544 100568 123912 100577
rect 123584 100528 123626 100568
rect 123666 100528 123708 100568
rect 123748 100528 123790 100568
rect 123830 100528 123872 100568
rect 123544 100519 123912 100528
rect 138664 100568 139032 100577
rect 138704 100528 138746 100568
rect 138786 100528 138828 100568
rect 138868 100528 138910 100568
rect 138950 100528 138992 100568
rect 138664 100519 139032 100528
rect 124784 99812 125152 99821
rect 124824 99772 124866 99812
rect 124906 99772 124948 99812
rect 124988 99772 125030 99812
rect 125070 99772 125112 99812
rect 124784 99763 125152 99772
rect 139904 99812 140272 99821
rect 139944 99772 139986 99812
rect 140026 99772 140068 99812
rect 140108 99772 140150 99812
rect 140190 99772 140232 99812
rect 139904 99763 140272 99772
rect 123544 99056 123912 99065
rect 123584 99016 123626 99056
rect 123666 99016 123708 99056
rect 123748 99016 123790 99056
rect 123830 99016 123872 99056
rect 123544 99007 123912 99016
rect 138664 99056 139032 99065
rect 138704 99016 138746 99056
rect 138786 99016 138828 99056
rect 138868 99016 138910 99056
rect 138950 99016 138992 99056
rect 138664 99007 139032 99016
rect 124784 98300 125152 98309
rect 124824 98260 124866 98300
rect 124906 98260 124948 98300
rect 124988 98260 125030 98300
rect 125070 98260 125112 98300
rect 124784 98251 125152 98260
rect 139904 98300 140272 98309
rect 139944 98260 139986 98300
rect 140026 98260 140068 98300
rect 140108 98260 140150 98300
rect 140190 98260 140232 98300
rect 139904 98251 140272 98260
rect 123544 97544 123912 97553
rect 123584 97504 123626 97544
rect 123666 97504 123708 97544
rect 123748 97504 123790 97544
rect 123830 97504 123872 97544
rect 123544 97495 123912 97504
rect 138664 97544 139032 97553
rect 138704 97504 138746 97544
rect 138786 97504 138828 97544
rect 138868 97504 138910 97544
rect 138950 97504 138992 97544
rect 138664 97495 139032 97504
rect 124784 96788 125152 96797
rect 124824 96748 124866 96788
rect 124906 96748 124948 96788
rect 124988 96748 125030 96788
rect 125070 96748 125112 96788
rect 124784 96739 125152 96748
rect 139904 96788 140272 96797
rect 139944 96748 139986 96788
rect 140026 96748 140068 96788
rect 140108 96748 140150 96788
rect 140190 96748 140232 96788
rect 139904 96739 140272 96748
rect 123544 96032 123912 96041
rect 123584 95992 123626 96032
rect 123666 95992 123708 96032
rect 123748 95992 123790 96032
rect 123830 95992 123872 96032
rect 123544 95983 123912 95992
rect 138664 96032 139032 96041
rect 138704 95992 138746 96032
rect 138786 95992 138828 96032
rect 138868 95992 138910 96032
rect 138950 95992 138992 96032
rect 138664 95983 139032 95992
rect 124784 95276 125152 95285
rect 124824 95236 124866 95276
rect 124906 95236 124948 95276
rect 124988 95236 125030 95276
rect 125070 95236 125112 95276
rect 124784 95227 125152 95236
rect 139904 95276 140272 95285
rect 139944 95236 139986 95276
rect 140026 95236 140068 95276
rect 140108 95236 140150 95276
rect 140190 95236 140232 95276
rect 139904 95227 140272 95236
rect 123544 94520 123912 94529
rect 123584 94480 123626 94520
rect 123666 94480 123708 94520
rect 123748 94480 123790 94520
rect 123830 94480 123872 94520
rect 123544 94471 123912 94480
rect 138664 94520 139032 94529
rect 138704 94480 138746 94520
rect 138786 94480 138828 94520
rect 138868 94480 138910 94520
rect 138950 94480 138992 94520
rect 138664 94471 139032 94480
rect 124784 93764 125152 93773
rect 124824 93724 124866 93764
rect 124906 93724 124948 93764
rect 124988 93724 125030 93764
rect 125070 93724 125112 93764
rect 124784 93715 125152 93724
rect 139904 93764 140272 93773
rect 139944 93724 139986 93764
rect 140026 93724 140068 93764
rect 140108 93724 140150 93764
rect 140190 93724 140232 93764
rect 139904 93715 140272 93724
rect 123544 93008 123912 93017
rect 123584 92968 123626 93008
rect 123666 92968 123708 93008
rect 123748 92968 123790 93008
rect 123830 92968 123872 93008
rect 123544 92959 123912 92968
rect 138664 93008 139032 93017
rect 138704 92968 138746 93008
rect 138786 92968 138828 93008
rect 138868 92968 138910 93008
rect 138950 92968 138992 93008
rect 138664 92959 139032 92968
rect 124784 92252 125152 92261
rect 124824 92212 124866 92252
rect 124906 92212 124948 92252
rect 124988 92212 125030 92252
rect 125070 92212 125112 92252
rect 124784 92203 125152 92212
rect 139904 92252 140272 92261
rect 139944 92212 139986 92252
rect 140026 92212 140068 92252
rect 140108 92212 140150 92252
rect 140190 92212 140232 92252
rect 139904 92203 140272 92212
rect 123544 91496 123912 91505
rect 123584 91456 123626 91496
rect 123666 91456 123708 91496
rect 123748 91456 123790 91496
rect 123830 91456 123872 91496
rect 123544 91447 123912 91456
rect 138664 91496 139032 91505
rect 138704 91456 138746 91496
rect 138786 91456 138828 91496
rect 138868 91456 138910 91496
rect 138950 91456 138992 91496
rect 138664 91447 139032 91456
rect 124784 90740 125152 90749
rect 124824 90700 124866 90740
rect 124906 90700 124948 90740
rect 124988 90700 125030 90740
rect 125070 90700 125112 90740
rect 124784 90691 125152 90700
rect 139904 90740 140272 90749
rect 139944 90700 139986 90740
rect 140026 90700 140068 90740
rect 140108 90700 140150 90740
rect 140190 90700 140232 90740
rect 139904 90691 140272 90700
rect 123544 89984 123912 89993
rect 123584 89944 123626 89984
rect 123666 89944 123708 89984
rect 123748 89944 123790 89984
rect 123830 89944 123872 89984
rect 123544 89935 123912 89944
rect 138664 89984 139032 89993
rect 138704 89944 138746 89984
rect 138786 89944 138828 89984
rect 138868 89944 138910 89984
rect 138950 89944 138992 89984
rect 138664 89935 139032 89944
rect 124784 89228 125152 89237
rect 124824 89188 124866 89228
rect 124906 89188 124948 89228
rect 124988 89188 125030 89228
rect 125070 89188 125112 89228
rect 124784 89179 125152 89188
rect 139904 89228 140272 89237
rect 139944 89188 139986 89228
rect 140026 89188 140068 89228
rect 140108 89188 140150 89228
rect 140190 89188 140232 89228
rect 139904 89179 140272 89188
rect 123544 88472 123912 88481
rect 123584 88432 123626 88472
rect 123666 88432 123708 88472
rect 123748 88432 123790 88472
rect 123830 88432 123872 88472
rect 123544 88423 123912 88432
rect 138664 88472 139032 88481
rect 138704 88432 138746 88472
rect 138786 88432 138828 88472
rect 138868 88432 138910 88472
rect 138950 88432 138992 88472
rect 138664 88423 139032 88432
rect 148204 87893 148244 87978
rect 148203 87884 148245 87893
rect 148203 87844 148204 87884
rect 148244 87844 148245 87884
rect 148203 87835 148245 87844
rect 124784 87716 125152 87725
rect 124824 87676 124866 87716
rect 124906 87676 124948 87716
rect 124988 87676 125030 87716
rect 125070 87676 125112 87716
rect 124784 87667 125152 87676
rect 139904 87716 140272 87725
rect 139944 87676 139986 87716
rect 140026 87676 140068 87716
rect 140108 87676 140150 87716
rect 140190 87676 140232 87716
rect 139904 87667 140272 87676
rect 123544 86960 123912 86969
rect 123584 86920 123626 86960
rect 123666 86920 123708 86960
rect 123748 86920 123790 86960
rect 123830 86920 123872 86960
rect 123544 86911 123912 86920
rect 138664 86960 139032 86969
rect 138704 86920 138746 86960
rect 138786 86920 138828 86960
rect 138868 86920 138910 86960
rect 138950 86920 138992 86960
rect 138664 86911 139032 86920
rect 124784 86204 125152 86213
rect 124824 86164 124866 86204
rect 124906 86164 124948 86204
rect 124988 86164 125030 86204
rect 125070 86164 125112 86204
rect 124784 86155 125152 86164
rect 139904 86204 140272 86213
rect 139944 86164 139986 86204
rect 140026 86164 140068 86204
rect 140108 86164 140150 86204
rect 140190 86164 140232 86204
rect 139904 86155 140272 86164
rect 123544 85448 123912 85457
rect 123584 85408 123626 85448
rect 123666 85408 123708 85448
rect 123748 85408 123790 85448
rect 123830 85408 123872 85448
rect 123544 85399 123912 85408
rect 138664 85448 139032 85457
rect 138704 85408 138746 85448
rect 138786 85408 138828 85448
rect 138868 85408 138910 85448
rect 138950 85408 138992 85448
rect 138664 85399 139032 85408
rect 124784 84692 125152 84701
rect 124824 84652 124866 84692
rect 124906 84652 124948 84692
rect 124988 84652 125030 84692
rect 125070 84652 125112 84692
rect 124784 84643 125152 84652
rect 139904 84692 140272 84701
rect 139944 84652 139986 84692
rect 140026 84652 140068 84692
rect 140108 84652 140150 84692
rect 140190 84652 140232 84692
rect 139904 84643 140272 84652
rect 123544 83936 123912 83945
rect 123584 83896 123626 83936
rect 123666 83896 123708 83936
rect 123748 83896 123790 83936
rect 123830 83896 123872 83936
rect 123544 83887 123912 83896
rect 138664 83936 139032 83945
rect 138704 83896 138746 83936
rect 138786 83896 138828 83936
rect 138868 83896 138910 83936
rect 138950 83896 138992 83936
rect 138664 83887 139032 83896
rect 124784 83180 125152 83189
rect 124824 83140 124866 83180
rect 124906 83140 124948 83180
rect 124988 83140 125030 83180
rect 125070 83140 125112 83180
rect 124784 83131 125152 83140
rect 139904 83180 140272 83189
rect 139944 83140 139986 83180
rect 140026 83140 140068 83180
rect 140108 83140 140150 83180
rect 140190 83140 140232 83180
rect 139904 83131 140272 83140
rect 123544 82424 123912 82433
rect 123584 82384 123626 82424
rect 123666 82384 123708 82424
rect 123748 82384 123790 82424
rect 123830 82384 123872 82424
rect 123544 82375 123912 82384
rect 138664 82424 139032 82433
rect 138704 82384 138746 82424
rect 138786 82384 138828 82424
rect 138868 82384 138910 82424
rect 138950 82384 138992 82424
rect 138664 82375 139032 82384
rect 124784 81668 125152 81677
rect 124824 81628 124866 81668
rect 124906 81628 124948 81668
rect 124988 81628 125030 81668
rect 125070 81628 125112 81668
rect 124784 81619 125152 81628
rect 139904 81668 140272 81677
rect 139944 81628 139986 81668
rect 140026 81628 140068 81668
rect 140108 81628 140150 81668
rect 140190 81628 140232 81668
rect 139904 81619 140272 81628
rect 123544 80912 123912 80921
rect 123584 80872 123626 80912
rect 123666 80872 123708 80912
rect 123748 80872 123790 80912
rect 123830 80872 123872 80912
rect 123544 80863 123912 80872
rect 138664 80912 139032 80921
rect 138704 80872 138746 80912
rect 138786 80872 138828 80912
rect 138868 80872 138910 80912
rect 138950 80872 138992 80912
rect 138664 80863 139032 80872
rect 124784 80156 125152 80165
rect 124824 80116 124866 80156
rect 124906 80116 124948 80156
rect 124988 80116 125030 80156
rect 125070 80116 125112 80156
rect 124784 80107 125152 80116
rect 139904 80156 140272 80165
rect 139944 80116 139986 80156
rect 140026 80116 140068 80156
rect 140108 80116 140150 80156
rect 140190 80116 140232 80156
rect 139904 80107 140272 80116
rect 123544 79400 123912 79409
rect 123584 79360 123626 79400
rect 123666 79360 123708 79400
rect 123748 79360 123790 79400
rect 123830 79360 123872 79400
rect 123544 79351 123912 79360
rect 138664 79400 139032 79409
rect 138704 79360 138746 79400
rect 138786 79360 138828 79400
rect 138868 79360 138910 79400
rect 138950 79360 138992 79400
rect 138664 79351 139032 79360
rect 124784 78644 125152 78653
rect 124824 78604 124866 78644
rect 124906 78604 124948 78644
rect 124988 78604 125030 78644
rect 125070 78604 125112 78644
rect 124784 78595 125152 78604
rect 139904 78644 140272 78653
rect 139944 78604 139986 78644
rect 140026 78604 140068 78644
rect 140108 78604 140150 78644
rect 140190 78604 140232 78644
rect 139904 78595 140272 78604
rect 123544 77888 123912 77897
rect 123584 77848 123626 77888
rect 123666 77848 123708 77888
rect 123748 77848 123790 77888
rect 123830 77848 123872 77888
rect 123544 77839 123912 77848
rect 138664 77888 139032 77897
rect 138704 77848 138746 77888
rect 138786 77848 138828 77888
rect 138868 77848 138910 77888
rect 138950 77848 138992 77888
rect 138664 77839 139032 77848
rect 124784 77132 125152 77141
rect 124824 77092 124866 77132
rect 124906 77092 124948 77132
rect 124988 77092 125030 77132
rect 125070 77092 125112 77132
rect 124784 77083 125152 77092
rect 139904 77132 140272 77141
rect 139944 77092 139986 77132
rect 140026 77092 140068 77132
rect 140108 77092 140150 77132
rect 140190 77092 140232 77132
rect 139904 77083 140272 77092
rect 123544 76376 123912 76385
rect 123584 76336 123626 76376
rect 123666 76336 123708 76376
rect 123748 76336 123790 76376
rect 123830 76336 123872 76376
rect 123544 76327 123912 76336
rect 138664 76376 139032 76385
rect 138704 76336 138746 76376
rect 138786 76336 138828 76376
rect 138868 76336 138910 76376
rect 138950 76336 138992 76376
rect 138664 76327 139032 76336
rect 148204 75788 148244 75797
rect 124784 75620 125152 75629
rect 124824 75580 124866 75620
rect 124906 75580 124948 75620
rect 124988 75580 125030 75620
rect 125070 75580 125112 75620
rect 124784 75571 125152 75580
rect 139904 75620 140272 75629
rect 139944 75580 139986 75620
rect 140026 75580 140068 75620
rect 140108 75580 140150 75620
rect 140190 75580 140232 75620
rect 139904 75571 140272 75580
rect 148204 72437 148244 75748
rect 148203 72428 148245 72437
rect 148203 72388 148204 72428
rect 148244 72388 148245 72428
rect 148203 72379 148245 72388
rect 87975 64324 88052 64364
rect 103975 64324 104084 64364
rect 119975 64324 120020 64364
rect 73323 64196 73365 64205
rect 73323 64156 73324 64196
rect 73364 64156 73365 64196
rect 73323 64147 73365 64156
rect 87975 63966 88015 64324
rect 103975 63966 104015 64324
rect 119975 63966 120015 64324
<< via2 >>
rect 112300 159664 112340 159704
rect 64108 152020 64148 152060
rect 94060 152020 94100 152060
rect 79424 148156 79464 148196
rect 79506 148156 79546 148196
rect 79588 148156 79628 148196
rect 79670 148156 79710 148196
rect 79752 148156 79792 148196
rect 78184 147400 78224 147440
rect 78266 147400 78306 147440
rect 78348 147400 78388 147440
rect 78430 147400 78470 147440
rect 78512 147400 78552 147440
rect 93304 147400 93344 147440
rect 93386 147400 93426 147440
rect 93468 147400 93508 147440
rect 93550 147400 93590 147440
rect 93632 147400 93672 147440
rect 79424 146644 79464 146684
rect 79506 146644 79546 146684
rect 79588 146644 79628 146684
rect 79670 146644 79710 146684
rect 79752 146644 79792 146684
rect 78184 145888 78224 145928
rect 78266 145888 78306 145928
rect 78348 145888 78388 145928
rect 78430 145888 78470 145928
rect 78512 145888 78552 145928
rect 93304 145888 93344 145928
rect 93386 145888 93426 145928
rect 93468 145888 93508 145928
rect 93550 145888 93590 145928
rect 93632 145888 93672 145928
rect 79424 145132 79464 145172
rect 79506 145132 79546 145172
rect 79588 145132 79628 145172
rect 79670 145132 79710 145172
rect 79752 145132 79792 145172
rect 78184 144376 78224 144416
rect 78266 144376 78306 144416
rect 78348 144376 78388 144416
rect 78430 144376 78470 144416
rect 78512 144376 78552 144416
rect 93304 144376 93344 144416
rect 93386 144376 93426 144416
rect 93468 144376 93508 144416
rect 93550 144376 93590 144416
rect 93632 144376 93672 144416
rect 79424 143620 79464 143660
rect 79506 143620 79546 143660
rect 79588 143620 79628 143660
rect 79670 143620 79710 143660
rect 79752 143620 79792 143660
rect 78184 142864 78224 142904
rect 78266 142864 78306 142904
rect 78348 142864 78388 142904
rect 78430 142864 78470 142904
rect 78512 142864 78552 142904
rect 93304 142864 93344 142904
rect 93386 142864 93426 142904
rect 93468 142864 93508 142904
rect 93550 142864 93590 142904
rect 93632 142864 93672 142904
rect 79424 142108 79464 142148
rect 79506 142108 79546 142148
rect 79588 142108 79628 142148
rect 79670 142108 79710 142148
rect 79752 142108 79792 142148
rect 78184 141352 78224 141392
rect 78266 141352 78306 141392
rect 78348 141352 78388 141392
rect 78430 141352 78470 141392
rect 78512 141352 78552 141392
rect 93304 141352 93344 141392
rect 93386 141352 93426 141392
rect 93468 141352 93508 141392
rect 93550 141352 93590 141392
rect 93632 141352 93672 141392
rect 79424 140596 79464 140636
rect 79506 140596 79546 140636
rect 79588 140596 79628 140636
rect 79670 140596 79710 140636
rect 79752 140596 79792 140636
rect 78184 139840 78224 139880
rect 78266 139840 78306 139880
rect 78348 139840 78388 139880
rect 78430 139840 78470 139880
rect 78512 139840 78552 139880
rect 93304 139840 93344 139880
rect 93386 139840 93426 139880
rect 93468 139840 93508 139880
rect 93550 139840 93590 139880
rect 93632 139840 93672 139880
rect 79424 139084 79464 139124
rect 79506 139084 79546 139124
rect 79588 139084 79628 139124
rect 79670 139084 79710 139124
rect 79752 139084 79792 139124
rect 78184 138328 78224 138368
rect 78266 138328 78306 138368
rect 78348 138328 78388 138368
rect 78430 138328 78470 138368
rect 78512 138328 78552 138368
rect 93304 138328 93344 138368
rect 93386 138328 93426 138368
rect 93468 138328 93508 138368
rect 93550 138328 93590 138368
rect 93632 138328 93672 138368
rect 79424 137572 79464 137612
rect 79506 137572 79546 137612
rect 79588 137572 79628 137612
rect 79670 137572 79710 137612
rect 79752 137572 79792 137612
rect 78184 136816 78224 136856
rect 78266 136816 78306 136856
rect 78348 136816 78388 136856
rect 78430 136816 78470 136856
rect 78512 136816 78552 136856
rect 93304 136816 93344 136856
rect 93386 136816 93426 136856
rect 93468 136816 93508 136856
rect 93550 136816 93590 136856
rect 93632 136816 93672 136856
rect 79424 136060 79464 136100
rect 79506 136060 79546 136100
rect 79588 136060 79628 136100
rect 79670 136060 79710 136100
rect 79752 136060 79792 136100
rect 78604 135472 78644 135512
rect 64108 135388 64148 135428
rect 78184 135304 78224 135344
rect 78266 135304 78306 135344
rect 78348 135304 78388 135344
rect 78430 135304 78470 135344
rect 78512 135304 78552 135344
rect 78184 133792 78224 133832
rect 78266 133792 78306 133832
rect 78348 133792 78388 133832
rect 78430 133792 78470 133832
rect 78512 133792 78552 133832
rect 93304 135304 93344 135344
rect 93386 135304 93426 135344
rect 93468 135304 93508 135344
rect 93550 135304 93590 135344
rect 93632 135304 93672 135344
rect 79424 134548 79464 134588
rect 79506 134548 79546 134588
rect 79588 134548 79628 134588
rect 79670 134548 79710 134588
rect 79752 134548 79792 134588
rect 93304 133792 93344 133832
rect 93386 133792 93426 133832
rect 93468 133792 93508 133832
rect 93550 133792 93590 133832
rect 93632 133792 93672 133832
rect 79424 133036 79464 133076
rect 79506 133036 79546 133076
rect 79588 133036 79628 133076
rect 79670 133036 79710 133076
rect 79752 133036 79792 133076
rect 79276 132532 79316 132572
rect 78184 132280 78224 132320
rect 78266 132280 78306 132320
rect 78348 132280 78388 132320
rect 78430 132280 78470 132320
rect 78512 132280 78552 132320
rect 93304 132280 93344 132320
rect 93386 132280 93426 132320
rect 93468 132280 93508 132320
rect 93550 132280 93590 132320
rect 93632 132280 93672 132320
rect 79424 131524 79464 131564
rect 79506 131524 79546 131564
rect 79588 131524 79628 131564
rect 79670 131524 79710 131564
rect 79752 131524 79792 131564
rect 78184 130768 78224 130808
rect 78266 130768 78306 130808
rect 78348 130768 78388 130808
rect 78430 130768 78470 130808
rect 78512 130768 78552 130808
rect 93304 130768 93344 130808
rect 93386 130768 93426 130808
rect 93468 130768 93508 130808
rect 93550 130768 93590 130808
rect 93632 130768 93672 130808
rect 79424 130012 79464 130052
rect 79506 130012 79546 130052
rect 79588 130012 79628 130052
rect 79670 130012 79710 130052
rect 79752 130012 79792 130052
rect 73324 129676 73364 129716
rect 64108 120856 64148 120896
rect 64108 104980 64148 105020
rect 64108 87970 64148 88010
rect 64108 71968 64148 72008
rect 78184 129256 78224 129296
rect 78266 129256 78306 129296
rect 78348 129256 78388 129296
rect 78430 129256 78470 129296
rect 78512 129256 78552 129296
rect 93304 129256 93344 129296
rect 93386 129256 93426 129296
rect 93468 129256 93508 129296
rect 93550 129256 93590 129296
rect 93632 129256 93672 129296
rect 79424 128500 79464 128540
rect 79506 128500 79546 128540
rect 79588 128500 79628 128540
rect 79670 128500 79710 128540
rect 79752 128500 79792 128540
rect 78184 127744 78224 127784
rect 78266 127744 78306 127784
rect 78348 127744 78388 127784
rect 78430 127744 78470 127784
rect 78512 127744 78552 127784
rect 93304 127744 93344 127784
rect 93386 127744 93426 127784
rect 93468 127744 93508 127784
rect 93550 127744 93590 127784
rect 93632 127744 93672 127784
rect 79852 127240 79892 127280
rect 79424 126988 79464 127028
rect 79506 126988 79546 127028
rect 79588 126988 79628 127028
rect 79670 126988 79710 127028
rect 79752 126988 79792 127028
rect 78184 126232 78224 126272
rect 78266 126232 78306 126272
rect 78348 126232 78388 126272
rect 78430 126232 78470 126272
rect 78512 126232 78552 126272
rect 79424 125476 79464 125516
rect 79506 125476 79546 125516
rect 79588 125476 79628 125516
rect 79670 125476 79710 125516
rect 79752 125476 79792 125516
rect 78184 124720 78224 124760
rect 78266 124720 78306 124760
rect 78348 124720 78388 124760
rect 78430 124720 78470 124760
rect 78512 124720 78552 124760
rect 93772 126568 93812 126608
rect 93304 126232 93344 126272
rect 93386 126232 93426 126272
rect 93468 126232 93508 126272
rect 93550 126232 93590 126272
rect 93632 126232 93672 126272
rect 93772 125224 93812 125264
rect 93304 124720 93344 124760
rect 93386 124720 93426 124760
rect 93468 124720 93508 124760
rect 93550 124720 93590 124760
rect 93632 124720 93672 124760
rect 94544 148156 94584 148196
rect 94626 148156 94666 148196
rect 94708 148156 94748 148196
rect 94790 148156 94830 148196
rect 94872 148156 94912 148196
rect 94544 146644 94584 146684
rect 94626 146644 94666 146684
rect 94708 146644 94748 146684
rect 94790 146644 94830 146684
rect 94872 146644 94912 146684
rect 94544 145132 94584 145172
rect 94626 145132 94666 145172
rect 94708 145132 94748 145172
rect 94790 145132 94830 145172
rect 94872 145132 94912 145172
rect 94544 143620 94584 143660
rect 94626 143620 94666 143660
rect 94708 143620 94748 143660
rect 94790 143620 94830 143660
rect 94872 143620 94912 143660
rect 94544 142108 94584 142148
rect 94626 142108 94666 142148
rect 94708 142108 94748 142148
rect 94790 142108 94830 142148
rect 94872 142108 94912 142148
rect 94544 140596 94584 140636
rect 94626 140596 94666 140636
rect 94708 140596 94748 140636
rect 94790 140596 94830 140636
rect 94872 140596 94912 140636
rect 94544 139084 94584 139124
rect 94626 139084 94666 139124
rect 94708 139084 94748 139124
rect 94790 139084 94830 139124
rect 94872 139084 94912 139124
rect 94544 137572 94584 137612
rect 94626 137572 94666 137612
rect 94708 137572 94748 137612
rect 94790 137572 94830 137612
rect 94872 137572 94912 137612
rect 94544 136060 94584 136100
rect 94626 136060 94666 136100
rect 94708 136060 94748 136100
rect 94790 136060 94830 136100
rect 94872 136060 94912 136100
rect 94544 134548 94584 134588
rect 94626 134548 94666 134588
rect 94708 134548 94748 134588
rect 94790 134548 94830 134588
rect 94872 134548 94912 134588
rect 97420 134212 97460 134252
rect 98188 134212 98228 134252
rect 98668 134212 98708 134252
rect 99820 134044 99860 134084
rect 100012 134044 100052 134084
rect 94544 133036 94584 133076
rect 94626 133036 94666 133076
rect 94708 133036 94748 133076
rect 94790 133036 94830 133076
rect 94872 133036 94912 133076
rect 94252 132532 94292 132572
rect 94156 129844 94196 129884
rect 94544 131524 94584 131564
rect 94626 131524 94666 131564
rect 94708 131524 94748 131564
rect 94790 131524 94830 131564
rect 94872 131524 94912 131564
rect 98764 132700 98804 132740
rect 100012 132700 100052 132740
rect 102220 132700 102260 132740
rect 102988 132700 103028 132740
rect 98860 132028 98900 132068
rect 99052 132028 99092 132068
rect 99436 132028 99476 132068
rect 99244 131692 99284 131732
rect 96844 130348 96884 130388
rect 94544 130012 94584 130052
rect 94626 130012 94666 130052
rect 94708 130012 94748 130052
rect 94790 130012 94830 130052
rect 94872 130012 94912 130052
rect 95020 129928 95060 129968
rect 94544 128500 94584 128540
rect 94626 128500 94666 128540
rect 94708 128500 94748 128540
rect 94790 128500 94830 128540
rect 94872 128500 94912 128540
rect 94828 128332 94868 128372
rect 96172 129844 96212 129884
rect 98092 130348 98132 130388
rect 99052 130348 99092 130388
rect 97228 130096 97268 130136
rect 97132 129928 97172 129968
rect 97420 129844 97460 129884
rect 96076 128332 96116 128372
rect 98956 129844 98996 129884
rect 95500 128248 95540 128288
rect 97996 128248 98036 128288
rect 94732 127324 94752 127364
rect 94752 127324 94772 127364
rect 94060 126820 94100 126860
rect 93964 126736 94004 126776
rect 94544 126988 94584 127028
rect 94626 126988 94666 127028
rect 94708 126988 94748 127028
rect 94790 126988 94830 127028
rect 94872 126988 94912 127028
rect 94636 126820 94676 126860
rect 94732 126736 94772 126776
rect 94252 126400 94292 126440
rect 78892 124300 78932 124340
rect 93868 124300 93908 124340
rect 78184 123208 78224 123248
rect 78266 123208 78306 123248
rect 78348 123208 78388 123248
rect 78430 123208 78470 123248
rect 78512 123208 78552 123248
rect 78184 121696 78224 121736
rect 78266 121696 78306 121736
rect 78348 121696 78388 121736
rect 78430 121696 78470 121736
rect 78512 121696 78552 121736
rect 79424 123964 79464 124004
rect 79506 123964 79546 124004
rect 79588 123964 79628 124004
rect 79670 123964 79710 124004
rect 79752 123964 79792 124004
rect 93304 123208 93344 123248
rect 93386 123208 93426 123248
rect 93468 123208 93508 123248
rect 93550 123208 93590 123248
rect 93632 123208 93672 123248
rect 79424 122452 79464 122492
rect 79506 122452 79546 122492
rect 79588 122452 79628 122492
rect 79670 122452 79710 122492
rect 79752 122452 79792 122492
rect 93772 122368 93812 122408
rect 93304 121696 93344 121736
rect 93386 121696 93426 121736
rect 93468 121696 93508 121736
rect 93550 121696 93590 121736
rect 93632 121696 93672 121736
rect 79424 120940 79464 120980
rect 79506 120940 79546 120980
rect 79588 120940 79628 120980
rect 79670 120940 79710 120980
rect 79752 120940 79792 120980
rect 78892 120856 78932 120896
rect 78184 120184 78224 120224
rect 78266 120184 78306 120224
rect 78348 120184 78388 120224
rect 78430 120184 78470 120224
rect 78512 120184 78552 120224
rect 93304 120184 93344 120224
rect 93386 120184 93426 120224
rect 93468 120184 93508 120224
rect 93550 120184 93590 120224
rect 93632 120184 93672 120224
rect 79424 119428 79464 119468
rect 79506 119428 79546 119468
rect 79588 119428 79628 119468
rect 79670 119428 79710 119468
rect 79752 119428 79792 119468
rect 78184 118672 78224 118712
rect 78266 118672 78306 118712
rect 78348 118672 78388 118712
rect 78430 118672 78470 118712
rect 78512 118672 78552 118712
rect 93304 118672 93344 118712
rect 93386 118672 93426 118712
rect 93468 118672 93508 118712
rect 93550 118672 93590 118712
rect 93632 118672 93672 118712
rect 79424 117916 79464 117956
rect 79506 117916 79546 117956
rect 79588 117916 79628 117956
rect 79670 117916 79710 117956
rect 79752 117916 79792 117956
rect 78184 117160 78224 117200
rect 78266 117160 78306 117200
rect 78348 117160 78388 117200
rect 78430 117160 78470 117200
rect 78512 117160 78552 117200
rect 93304 117160 93344 117200
rect 93386 117160 93426 117200
rect 93468 117160 93508 117200
rect 93550 117160 93590 117200
rect 93632 117160 93672 117200
rect 79424 116404 79464 116444
rect 79506 116404 79546 116444
rect 79588 116404 79628 116444
rect 79670 116404 79710 116444
rect 79752 116404 79792 116444
rect 78184 115648 78224 115688
rect 78266 115648 78306 115688
rect 78348 115648 78388 115688
rect 78430 115648 78470 115688
rect 78512 115648 78552 115688
rect 93304 115648 93344 115688
rect 93386 115648 93426 115688
rect 93468 115648 93508 115688
rect 93550 115648 93590 115688
rect 93632 115648 93672 115688
rect 79424 114892 79464 114932
rect 79506 114892 79546 114932
rect 79588 114892 79628 114932
rect 79670 114892 79710 114932
rect 79752 114892 79792 114932
rect 78184 114136 78224 114176
rect 78266 114136 78306 114176
rect 78348 114136 78388 114176
rect 78430 114136 78470 114176
rect 78512 114136 78552 114176
rect 93304 114136 93344 114176
rect 93386 114136 93426 114176
rect 93468 114136 93508 114176
rect 93550 114136 93590 114176
rect 93632 114136 93672 114176
rect 79424 113380 79464 113420
rect 79506 113380 79546 113420
rect 79588 113380 79628 113420
rect 79670 113380 79710 113420
rect 79752 113380 79792 113420
rect 78184 112624 78224 112664
rect 78266 112624 78306 112664
rect 78348 112624 78388 112664
rect 78430 112624 78470 112664
rect 78512 112624 78552 112664
rect 93304 112624 93344 112664
rect 93386 112624 93426 112664
rect 93468 112624 93508 112664
rect 93550 112624 93590 112664
rect 93632 112624 93672 112664
rect 79424 111868 79464 111908
rect 79506 111868 79546 111908
rect 79588 111868 79628 111908
rect 79670 111868 79710 111908
rect 79752 111868 79792 111908
rect 78184 111112 78224 111152
rect 78266 111112 78306 111152
rect 78348 111112 78388 111152
rect 78430 111112 78470 111152
rect 78512 111112 78552 111152
rect 93304 111112 93344 111152
rect 93386 111112 93426 111152
rect 93468 111112 93508 111152
rect 93550 111112 93590 111152
rect 93632 111112 93672 111152
rect 79424 110356 79464 110396
rect 79506 110356 79546 110396
rect 79588 110356 79628 110396
rect 79670 110356 79710 110396
rect 79752 110356 79792 110396
rect 78184 109600 78224 109640
rect 78266 109600 78306 109640
rect 78348 109600 78388 109640
rect 78430 109600 78470 109640
rect 78512 109600 78552 109640
rect 93304 109600 93344 109640
rect 93386 109600 93426 109640
rect 93468 109600 93508 109640
rect 93550 109600 93590 109640
rect 93632 109600 93672 109640
rect 79424 108844 79464 108884
rect 79506 108844 79546 108884
rect 79588 108844 79628 108884
rect 79670 108844 79710 108884
rect 79752 108844 79792 108884
rect 78184 108088 78224 108128
rect 78266 108088 78306 108128
rect 78348 108088 78388 108128
rect 78430 108088 78470 108128
rect 78512 108088 78552 108128
rect 93304 108088 93344 108128
rect 93386 108088 93426 108128
rect 93468 108088 93508 108128
rect 93550 108088 93590 108128
rect 93632 108088 93672 108128
rect 79424 107332 79464 107372
rect 79506 107332 79546 107372
rect 79588 107332 79628 107372
rect 79670 107332 79710 107372
rect 79752 107332 79792 107372
rect 78184 106576 78224 106616
rect 78266 106576 78306 106616
rect 78348 106576 78388 106616
rect 78430 106576 78470 106616
rect 78512 106576 78552 106616
rect 93304 106576 93344 106616
rect 93386 106576 93426 106616
rect 93468 106576 93508 106616
rect 93550 106576 93590 106616
rect 93632 106576 93672 106616
rect 79424 105820 79464 105860
rect 79506 105820 79546 105860
rect 79588 105820 79628 105860
rect 79670 105820 79710 105860
rect 79752 105820 79792 105860
rect 78184 105064 78224 105104
rect 78266 105064 78306 105104
rect 78348 105064 78388 105104
rect 78430 105064 78470 105104
rect 78512 105064 78552 105104
rect 93304 105064 93344 105104
rect 93386 105064 93426 105104
rect 93468 105064 93508 105104
rect 93550 105064 93590 105104
rect 93632 105064 93672 105104
rect 79424 104308 79464 104348
rect 79506 104308 79546 104348
rect 79588 104308 79628 104348
rect 79670 104308 79710 104348
rect 79752 104308 79792 104348
rect 78184 103552 78224 103592
rect 78266 103552 78306 103592
rect 78348 103552 78388 103592
rect 78430 103552 78470 103592
rect 78512 103552 78552 103592
rect 93304 103552 93344 103592
rect 93386 103552 93426 103592
rect 93468 103552 93508 103592
rect 93550 103552 93590 103592
rect 93632 103552 93672 103592
rect 79424 102796 79464 102836
rect 79506 102796 79546 102836
rect 79588 102796 79628 102836
rect 79670 102796 79710 102836
rect 79752 102796 79792 102836
rect 78184 102040 78224 102080
rect 78266 102040 78306 102080
rect 78348 102040 78388 102080
rect 78430 102040 78470 102080
rect 78512 102040 78552 102080
rect 93304 102040 93344 102080
rect 93386 102040 93426 102080
rect 93468 102040 93508 102080
rect 93550 102040 93590 102080
rect 93632 102040 93672 102080
rect 79424 101284 79464 101324
rect 79506 101284 79546 101324
rect 79588 101284 79628 101324
rect 79670 101284 79710 101324
rect 79752 101284 79792 101324
rect 78184 100528 78224 100568
rect 78266 100528 78306 100568
rect 78348 100528 78388 100568
rect 78430 100528 78470 100568
rect 78512 100528 78552 100568
rect 93304 100528 93344 100568
rect 93386 100528 93426 100568
rect 93468 100528 93508 100568
rect 93550 100528 93590 100568
rect 93632 100528 93672 100568
rect 79424 99772 79464 99812
rect 79506 99772 79546 99812
rect 79588 99772 79628 99812
rect 79670 99772 79710 99812
rect 79752 99772 79792 99812
rect 78184 99016 78224 99056
rect 78266 99016 78306 99056
rect 78348 99016 78388 99056
rect 78430 99016 78470 99056
rect 78512 99016 78552 99056
rect 93304 99016 93344 99056
rect 93386 99016 93426 99056
rect 93468 99016 93508 99056
rect 93550 99016 93590 99056
rect 93632 99016 93672 99056
rect 79424 98260 79464 98300
rect 79506 98260 79546 98300
rect 79588 98260 79628 98300
rect 79670 98260 79710 98300
rect 79752 98260 79792 98300
rect 78184 97504 78224 97544
rect 78266 97504 78306 97544
rect 78348 97504 78388 97544
rect 78430 97504 78470 97544
rect 78512 97504 78552 97544
rect 93304 97504 93344 97544
rect 93386 97504 93426 97544
rect 93468 97504 93508 97544
rect 93550 97504 93590 97544
rect 93632 97504 93672 97544
rect 79424 96748 79464 96788
rect 79506 96748 79546 96788
rect 79588 96748 79628 96788
rect 79670 96748 79710 96788
rect 79752 96748 79792 96788
rect 78184 95992 78224 96032
rect 78266 95992 78306 96032
rect 78348 95992 78388 96032
rect 78430 95992 78470 96032
rect 78512 95992 78552 96032
rect 93304 95992 93344 96032
rect 93386 95992 93426 96032
rect 93468 95992 93508 96032
rect 93550 95992 93590 96032
rect 93632 95992 93672 96032
rect 88012 95572 88052 95612
rect 79424 95236 79464 95276
rect 79506 95236 79546 95276
rect 79588 95236 79628 95276
rect 79670 95236 79710 95276
rect 79752 95236 79792 95276
rect 78184 94480 78224 94520
rect 78266 94480 78306 94520
rect 78348 94480 78388 94520
rect 78430 94480 78470 94520
rect 78512 94480 78552 94520
rect 79424 93724 79464 93764
rect 79506 93724 79546 93764
rect 79588 93724 79628 93764
rect 79670 93724 79710 93764
rect 79752 93724 79792 93764
rect 78184 92968 78224 93008
rect 78266 92968 78306 93008
rect 78348 92968 78388 93008
rect 78430 92968 78470 93008
rect 78512 92968 78552 93008
rect 79424 92212 79464 92252
rect 79506 92212 79546 92252
rect 79588 92212 79628 92252
rect 79670 92212 79710 92252
rect 79752 92212 79792 92252
rect 78184 91456 78224 91496
rect 78266 91456 78306 91496
rect 78348 91456 78388 91496
rect 78430 91456 78470 91496
rect 78512 91456 78552 91496
rect 79424 90700 79464 90740
rect 79506 90700 79546 90740
rect 79588 90700 79628 90740
rect 79670 90700 79710 90740
rect 79752 90700 79792 90740
rect 78184 89944 78224 89984
rect 78266 89944 78306 89984
rect 78348 89944 78388 89984
rect 78430 89944 78470 89984
rect 78512 89944 78552 89984
rect 79424 89188 79464 89228
rect 79506 89188 79546 89228
rect 79588 89188 79628 89228
rect 79670 89188 79710 89228
rect 79752 89188 79792 89228
rect 78184 88432 78224 88472
rect 78266 88432 78306 88472
rect 78348 88432 78388 88472
rect 78430 88432 78470 88472
rect 78512 88432 78552 88472
rect 79424 87676 79464 87716
rect 79506 87676 79546 87716
rect 79588 87676 79628 87716
rect 79670 87676 79710 87716
rect 79752 87676 79792 87716
rect 78184 86920 78224 86960
rect 78266 86920 78306 86960
rect 78348 86920 78388 86960
rect 78430 86920 78470 86960
rect 78512 86920 78552 86960
rect 79424 86164 79464 86204
rect 79506 86164 79546 86204
rect 79588 86164 79628 86204
rect 79670 86164 79710 86204
rect 79752 86164 79792 86204
rect 78184 85408 78224 85448
rect 78266 85408 78306 85448
rect 78348 85408 78388 85448
rect 78430 85408 78470 85448
rect 78512 85408 78552 85448
rect 79424 84652 79464 84692
rect 79506 84652 79546 84692
rect 79588 84652 79628 84692
rect 79670 84652 79710 84692
rect 79752 84652 79792 84692
rect 78184 83896 78224 83936
rect 78266 83896 78306 83936
rect 78348 83896 78388 83936
rect 78430 83896 78470 83936
rect 78512 83896 78552 83936
rect 79424 83140 79464 83180
rect 79506 83140 79546 83180
rect 79588 83140 79628 83180
rect 79670 83140 79710 83180
rect 79752 83140 79792 83180
rect 78184 82384 78224 82424
rect 78266 82384 78306 82424
rect 78348 82384 78388 82424
rect 78430 82384 78470 82424
rect 78512 82384 78552 82424
rect 79424 81628 79464 81668
rect 79506 81628 79546 81668
rect 79588 81628 79628 81668
rect 79670 81628 79710 81668
rect 79752 81628 79792 81668
rect 78184 80872 78224 80912
rect 78266 80872 78306 80912
rect 78348 80872 78388 80912
rect 78430 80872 78470 80912
rect 78512 80872 78552 80912
rect 79424 80116 79464 80156
rect 79506 80116 79546 80156
rect 79588 80116 79628 80156
rect 79670 80116 79710 80156
rect 79752 80116 79792 80156
rect 78184 79360 78224 79400
rect 78266 79360 78306 79400
rect 78348 79360 78388 79400
rect 78430 79360 78470 79400
rect 78512 79360 78552 79400
rect 79424 78604 79464 78644
rect 79506 78604 79546 78644
rect 79588 78604 79628 78644
rect 79670 78604 79710 78644
rect 79752 78604 79792 78644
rect 78184 77848 78224 77888
rect 78266 77848 78306 77888
rect 78348 77848 78388 77888
rect 78430 77848 78470 77888
rect 78512 77848 78552 77888
rect 79424 77092 79464 77132
rect 79506 77092 79546 77132
rect 79588 77092 79628 77132
rect 79670 77092 79710 77132
rect 79752 77092 79792 77132
rect 78184 76336 78224 76376
rect 78266 76336 78306 76376
rect 78348 76336 78388 76376
rect 78430 76336 78470 76376
rect 78512 76336 78552 76376
rect 79424 75580 79464 75620
rect 79506 75580 79546 75620
rect 79588 75580 79628 75620
rect 79670 75580 79710 75620
rect 79752 75580 79792 75620
rect 93304 94480 93344 94520
rect 93386 94480 93426 94520
rect 93468 94480 93508 94520
rect 93550 94480 93590 94520
rect 93632 94480 93672 94520
rect 93304 92968 93344 93008
rect 93386 92968 93426 93008
rect 93468 92968 93508 93008
rect 93550 92968 93590 93008
rect 93632 92968 93672 93008
rect 93304 91456 93344 91496
rect 93386 91456 93426 91496
rect 93468 91456 93508 91496
rect 93550 91456 93590 91496
rect 93632 91456 93672 91496
rect 93304 89944 93344 89984
rect 93386 89944 93426 89984
rect 93468 89944 93508 89984
rect 93550 89944 93590 89984
rect 93632 89944 93672 89984
rect 93304 88432 93344 88472
rect 93386 88432 93426 88472
rect 93468 88432 93508 88472
rect 93550 88432 93590 88472
rect 93632 88432 93672 88472
rect 93304 86920 93344 86960
rect 93386 86920 93426 86960
rect 93468 86920 93508 86960
rect 93550 86920 93590 86960
rect 93632 86920 93672 86960
rect 93304 85408 93344 85448
rect 93386 85408 93426 85448
rect 93468 85408 93508 85448
rect 93550 85408 93590 85448
rect 93632 85408 93672 85448
rect 93304 83896 93344 83936
rect 93386 83896 93426 83936
rect 93468 83896 93508 83936
rect 93550 83896 93590 83936
rect 93632 83896 93672 83936
rect 93304 82384 93344 82424
rect 93386 82384 93426 82424
rect 93468 82384 93508 82424
rect 93550 82384 93590 82424
rect 93632 82384 93672 82424
rect 93304 80872 93344 80912
rect 93386 80872 93426 80912
rect 93468 80872 93508 80912
rect 93550 80872 93590 80912
rect 93632 80872 93672 80912
rect 93304 79360 93344 79400
rect 93386 79360 93426 79400
rect 93468 79360 93508 79400
rect 93550 79360 93590 79400
rect 93632 79360 93672 79400
rect 93304 77848 93344 77888
rect 93386 77848 93426 77888
rect 93468 77848 93508 77888
rect 93550 77848 93590 77888
rect 93632 77848 93672 77888
rect 93304 76336 93344 76376
rect 93386 76336 93426 76376
rect 93468 76336 93508 76376
rect 93550 76336 93590 76376
rect 93632 76336 93672 76376
rect 94924 126652 94964 126692
rect 94828 126568 94868 126608
rect 95020 126568 95060 126608
rect 99148 130264 99188 130304
rect 101356 132616 101396 132656
rect 101068 132028 101108 132068
rect 99532 131944 99572 131984
rect 100012 131944 100052 131984
rect 100204 131860 100244 131900
rect 101164 131944 101204 131984
rect 99340 131020 99380 131060
rect 99916 130096 99956 130136
rect 99916 129928 99956 129968
rect 101356 131860 101396 131900
rect 101548 131692 101588 131732
rect 101260 131272 101300 131312
rect 100588 131188 100628 131228
rect 109664 148156 109704 148196
rect 109746 148156 109786 148196
rect 109828 148156 109868 148196
rect 109910 148156 109950 148196
rect 109992 148156 110032 148196
rect 108424 147400 108464 147440
rect 108506 147400 108546 147440
rect 108588 147400 108628 147440
rect 108670 147400 108710 147440
rect 108752 147400 108792 147440
rect 109664 146644 109704 146684
rect 109746 146644 109786 146684
rect 109828 146644 109868 146684
rect 109910 146644 109950 146684
rect 109992 146644 110032 146684
rect 108424 145888 108464 145928
rect 108506 145888 108546 145928
rect 108588 145888 108628 145928
rect 108670 145888 108710 145928
rect 108752 145888 108792 145928
rect 109664 145132 109704 145172
rect 109746 145132 109786 145172
rect 109828 145132 109868 145172
rect 109910 145132 109950 145172
rect 109992 145132 110032 145172
rect 108424 144376 108464 144416
rect 108506 144376 108546 144416
rect 108588 144376 108628 144416
rect 108670 144376 108710 144416
rect 108752 144376 108792 144416
rect 109664 143620 109704 143660
rect 109746 143620 109786 143660
rect 109828 143620 109868 143660
rect 109910 143620 109950 143660
rect 109992 143620 110032 143660
rect 108424 142864 108464 142904
rect 108506 142864 108546 142904
rect 108588 142864 108628 142904
rect 108670 142864 108710 142904
rect 108752 142864 108792 142904
rect 109664 142108 109704 142148
rect 109746 142108 109786 142148
rect 109828 142108 109868 142148
rect 109910 142108 109950 142148
rect 109992 142108 110032 142148
rect 108424 141352 108464 141392
rect 108506 141352 108546 141392
rect 108588 141352 108628 141392
rect 108670 141352 108710 141392
rect 108752 141352 108792 141392
rect 109664 140596 109704 140636
rect 109746 140596 109786 140636
rect 109828 140596 109868 140636
rect 109910 140596 109950 140636
rect 109992 140596 110032 140636
rect 108424 139840 108464 139880
rect 108506 139840 108546 139880
rect 108588 139840 108628 139880
rect 108670 139840 108710 139880
rect 108752 139840 108792 139880
rect 109664 139084 109704 139124
rect 109746 139084 109786 139124
rect 109828 139084 109868 139124
rect 109910 139084 109950 139124
rect 109992 139084 110032 139124
rect 108424 138328 108464 138368
rect 108506 138328 108546 138368
rect 108588 138328 108628 138368
rect 108670 138328 108710 138368
rect 108752 138328 108792 138368
rect 109664 137572 109704 137612
rect 109746 137572 109786 137612
rect 109828 137572 109868 137612
rect 109910 137572 109950 137612
rect 109992 137572 110032 137612
rect 108424 136816 108464 136856
rect 108506 136816 108546 136856
rect 108588 136816 108628 136856
rect 108670 136816 108710 136856
rect 108752 136816 108792 136856
rect 109664 136060 109704 136100
rect 109746 136060 109786 136100
rect 109828 136060 109868 136100
rect 109910 136060 109950 136100
rect 109992 136060 110032 136100
rect 108424 135304 108464 135344
rect 108506 135304 108546 135344
rect 108588 135304 108628 135344
rect 108670 135304 108710 135344
rect 108752 135304 108792 135344
rect 109664 134548 109704 134588
rect 109746 134548 109786 134588
rect 109828 134548 109868 134588
rect 109910 134548 109950 134588
rect 109992 134548 110032 134588
rect 105100 134212 105140 134252
rect 108424 133792 108464 133832
rect 108506 133792 108546 133832
rect 108588 133792 108628 133832
rect 108670 133792 108710 133832
rect 108752 133792 108792 133832
rect 109664 133036 109704 133076
rect 109746 133036 109786 133076
rect 109828 133036 109868 133076
rect 109910 133036 109950 133076
rect 109992 133036 110032 133076
rect 103948 131440 103988 131480
rect 102124 131272 102164 131312
rect 102028 131188 102068 131228
rect 102220 131020 102260 131060
rect 101644 130348 101684 130388
rect 103084 130264 103124 130304
rect 100108 129844 100148 129884
rect 103084 129844 103124 129884
rect 103468 131188 103508 131228
rect 104332 131104 104372 131144
rect 103564 131020 103604 131060
rect 104044 131020 104084 131060
rect 103468 130264 103508 130304
rect 103276 130180 103316 130220
rect 99148 128164 99188 128180
rect 99148 128140 99188 128164
rect 95596 126484 95636 126524
rect 95884 126652 95924 126692
rect 95788 126568 95828 126608
rect 104044 126568 104084 126608
rect 95692 126400 95732 126440
rect 94544 125476 94584 125516
rect 94626 125476 94666 125516
rect 94708 125476 94748 125516
rect 94790 125476 94830 125516
rect 94872 125476 94912 125516
rect 94544 123964 94584 124004
rect 94626 123964 94666 124004
rect 94708 123964 94748 124004
rect 94790 123964 94830 124004
rect 94872 123964 94912 124004
rect 94544 122452 94584 122492
rect 94626 122452 94666 122492
rect 94708 122452 94748 122492
rect 94790 122452 94830 122492
rect 94872 122452 94912 122492
rect 94544 120940 94584 120980
rect 94626 120940 94666 120980
rect 94708 120940 94748 120980
rect 94790 120940 94830 120980
rect 94872 120940 94912 120980
rect 94544 119428 94584 119468
rect 94626 119428 94666 119468
rect 94708 119428 94748 119468
rect 94790 119428 94830 119468
rect 94872 119428 94912 119468
rect 94544 117916 94584 117956
rect 94626 117916 94666 117956
rect 94708 117916 94748 117956
rect 94790 117916 94830 117956
rect 94872 117916 94912 117956
rect 94544 116404 94584 116444
rect 94626 116404 94666 116444
rect 94708 116404 94748 116444
rect 94790 116404 94830 116444
rect 94872 116404 94912 116444
rect 94544 114892 94584 114932
rect 94626 114892 94666 114932
rect 94708 114892 94748 114932
rect 94790 114892 94830 114932
rect 94872 114892 94912 114932
rect 94544 113380 94584 113420
rect 94626 113380 94666 113420
rect 94708 113380 94748 113420
rect 94790 113380 94830 113420
rect 94872 113380 94912 113420
rect 94544 111868 94584 111908
rect 94626 111868 94666 111908
rect 94708 111868 94748 111908
rect 94790 111868 94830 111908
rect 94872 111868 94912 111908
rect 94544 110356 94584 110396
rect 94626 110356 94666 110396
rect 94708 110356 94748 110396
rect 94790 110356 94830 110396
rect 94872 110356 94912 110396
rect 94544 108844 94584 108884
rect 94626 108844 94666 108884
rect 94708 108844 94748 108884
rect 94790 108844 94830 108884
rect 94872 108844 94912 108884
rect 94544 107332 94584 107372
rect 94626 107332 94666 107372
rect 94708 107332 94748 107372
rect 94790 107332 94830 107372
rect 94872 107332 94912 107372
rect 94544 105820 94584 105860
rect 94626 105820 94666 105860
rect 94708 105820 94748 105860
rect 94790 105820 94830 105860
rect 94872 105820 94912 105860
rect 94444 104980 94484 105020
rect 94544 104308 94584 104348
rect 94626 104308 94666 104348
rect 94708 104308 94748 104348
rect 94790 104308 94830 104348
rect 94872 104308 94912 104348
rect 94544 102796 94584 102836
rect 94626 102796 94666 102836
rect 94708 102796 94748 102836
rect 94790 102796 94830 102836
rect 94872 102796 94912 102836
rect 94544 101284 94584 101324
rect 94626 101284 94666 101324
rect 94708 101284 94748 101324
rect 94790 101284 94830 101324
rect 94872 101284 94912 101324
rect 94544 99772 94584 99812
rect 94626 99772 94666 99812
rect 94708 99772 94748 99812
rect 94790 99772 94830 99812
rect 94872 99772 94912 99812
rect 94544 98260 94584 98300
rect 94626 98260 94666 98300
rect 94708 98260 94748 98300
rect 94790 98260 94830 98300
rect 94872 98260 94912 98300
rect 94544 96748 94584 96788
rect 94626 96748 94666 96788
rect 94708 96748 94748 96788
rect 94790 96748 94830 96788
rect 94872 96748 94912 96788
rect 103660 95572 103700 95612
rect 94544 95236 94584 95276
rect 94626 95236 94666 95276
rect 94708 95236 94748 95276
rect 94790 95236 94830 95276
rect 94872 95236 94912 95276
rect 94544 93724 94584 93764
rect 94626 93724 94666 93764
rect 94708 93724 94748 93764
rect 94790 93724 94830 93764
rect 94872 93724 94912 93764
rect 94544 92212 94584 92252
rect 94626 92212 94666 92252
rect 94708 92212 94748 92252
rect 94790 92212 94830 92252
rect 94872 92212 94912 92252
rect 94544 90700 94584 90740
rect 94626 90700 94666 90740
rect 94708 90700 94748 90740
rect 94790 90700 94830 90740
rect 94872 90700 94912 90740
rect 94544 89188 94584 89228
rect 94626 89188 94666 89228
rect 94708 89188 94748 89228
rect 94790 89188 94830 89228
rect 94872 89188 94912 89228
rect 94252 89104 94292 89144
rect 94544 87676 94584 87716
rect 94626 87676 94666 87716
rect 94708 87676 94748 87716
rect 94790 87676 94830 87716
rect 94872 87676 94912 87716
rect 94544 86164 94584 86204
rect 94626 86164 94666 86204
rect 94708 86164 94748 86204
rect 94790 86164 94830 86204
rect 94872 86164 94912 86204
rect 94544 84652 94584 84692
rect 94626 84652 94666 84692
rect 94708 84652 94748 84692
rect 94790 84652 94830 84692
rect 94872 84652 94912 84692
rect 94544 83140 94584 83180
rect 94626 83140 94666 83180
rect 94708 83140 94748 83180
rect 94790 83140 94830 83180
rect 94872 83140 94912 83180
rect 94544 81628 94584 81668
rect 94626 81628 94666 81668
rect 94708 81628 94748 81668
rect 94790 81628 94830 81668
rect 94872 81628 94912 81668
rect 94544 80116 94584 80156
rect 94626 80116 94666 80156
rect 94708 80116 94748 80156
rect 94790 80116 94830 80156
rect 94872 80116 94912 80156
rect 94544 78604 94584 78644
rect 94626 78604 94666 78644
rect 94708 78604 94748 78644
rect 94790 78604 94830 78644
rect 94872 78604 94912 78644
rect 94544 77092 94584 77132
rect 94626 77092 94666 77132
rect 94708 77092 94748 77132
rect 94790 77092 94830 77132
rect 94872 77092 94912 77132
rect 94544 75580 94584 75620
rect 94626 75580 94666 75620
rect 94708 75580 94748 75620
rect 94790 75580 94830 75620
rect 94872 75580 94912 75620
rect 93772 71212 93812 71252
rect 106252 132616 106292 132656
rect 108424 132280 108464 132320
rect 108506 132280 108546 132320
rect 108588 132280 108628 132320
rect 108670 132280 108710 132320
rect 108752 132280 108792 132320
rect 108748 131608 108788 131648
rect 109664 131524 109704 131564
rect 109746 131524 109786 131564
rect 109828 131524 109868 131564
rect 109910 131524 109950 131564
rect 109992 131524 110032 131564
rect 109036 131188 109076 131228
rect 108748 131104 108788 131144
rect 108940 131104 108980 131144
rect 109420 131356 109460 131396
rect 109804 131356 109844 131396
rect 110380 131356 110420 131396
rect 109420 131188 109460 131228
rect 109132 131104 109172 131144
rect 110476 131188 110516 131228
rect 110380 131104 110420 131144
rect 109612 131020 109652 131060
rect 108424 130768 108464 130808
rect 108506 130768 108546 130808
rect 108588 130768 108628 130808
rect 108670 130768 108710 130808
rect 108752 130768 108792 130808
rect 105100 130684 105140 130724
rect 104716 130180 104756 130220
rect 108748 130600 108788 130640
rect 105388 130348 105428 130388
rect 105964 130348 106004 130388
rect 110188 130348 110228 130388
rect 110572 131020 110612 131060
rect 110764 131776 110804 131816
rect 111436 131440 111476 131480
rect 111820 131440 111860 131480
rect 110764 131356 110804 131396
rect 115948 151600 115988 151640
rect 124784 148156 124824 148196
rect 124866 148156 124906 148196
rect 124948 148156 124988 148196
rect 125030 148156 125070 148196
rect 125112 148156 125152 148196
rect 123544 147400 123584 147440
rect 123626 147400 123666 147440
rect 123708 147400 123748 147440
rect 123790 147400 123830 147440
rect 123872 147400 123912 147440
rect 124784 146644 124824 146684
rect 124866 146644 124906 146684
rect 124948 146644 124988 146684
rect 125030 146644 125070 146684
rect 125112 146644 125152 146684
rect 123544 145888 123584 145928
rect 123626 145888 123666 145928
rect 123708 145888 123748 145928
rect 123790 145888 123830 145928
rect 123872 145888 123912 145928
rect 124784 145132 124824 145172
rect 124866 145132 124906 145172
rect 124948 145132 124988 145172
rect 125030 145132 125070 145172
rect 125112 145132 125152 145172
rect 123544 144376 123584 144416
rect 123626 144376 123666 144416
rect 123708 144376 123748 144416
rect 123790 144376 123830 144416
rect 123872 144376 123912 144416
rect 124784 143620 124824 143660
rect 124866 143620 124906 143660
rect 124948 143620 124988 143660
rect 125030 143620 125070 143660
rect 125112 143620 125152 143660
rect 123544 142864 123584 142904
rect 123626 142864 123666 142904
rect 123708 142864 123748 142904
rect 123790 142864 123830 142904
rect 123872 142864 123912 142904
rect 124784 142108 124824 142148
rect 124866 142108 124906 142148
rect 124948 142108 124988 142148
rect 125030 142108 125070 142148
rect 125112 142108 125152 142148
rect 123544 141352 123584 141392
rect 123626 141352 123666 141392
rect 123708 141352 123748 141392
rect 123790 141352 123830 141392
rect 123872 141352 123912 141392
rect 124784 140596 124824 140636
rect 124866 140596 124906 140636
rect 124948 140596 124988 140636
rect 125030 140596 125070 140636
rect 125112 140596 125152 140636
rect 123544 139840 123584 139880
rect 123626 139840 123666 139880
rect 123708 139840 123748 139880
rect 123790 139840 123830 139880
rect 123872 139840 123912 139880
rect 124784 139084 124824 139124
rect 124866 139084 124906 139124
rect 124948 139084 124988 139124
rect 125030 139084 125070 139124
rect 125112 139084 125152 139124
rect 123544 138328 123584 138368
rect 123626 138328 123666 138368
rect 123708 138328 123748 138368
rect 123790 138328 123830 138368
rect 123872 138328 123912 138368
rect 124784 137572 124824 137612
rect 124866 137572 124906 137612
rect 124948 137572 124988 137612
rect 125030 137572 125070 137612
rect 125112 137572 125152 137612
rect 123544 136816 123584 136856
rect 123626 136816 123666 136856
rect 123708 136816 123748 136856
rect 123790 136816 123830 136856
rect 123872 136816 123912 136856
rect 124784 136060 124824 136100
rect 124866 136060 124906 136100
rect 124948 136060 124988 136100
rect 125030 136060 125070 136100
rect 125112 136060 125152 136100
rect 121804 135556 121844 135596
rect 112876 133204 112916 133244
rect 112396 131776 112404 131816
rect 112404 131776 112436 131816
rect 112588 131692 112628 131732
rect 112300 131356 112340 131396
rect 110764 130936 110804 130976
rect 112204 130936 112244 130976
rect 110668 130600 110708 130640
rect 105964 130180 106004 130220
rect 110668 130180 110708 130220
rect 109664 130012 109704 130052
rect 109746 130012 109786 130052
rect 109828 130012 109868 130052
rect 109910 130012 109950 130052
rect 109992 130012 110032 130052
rect 112012 130348 112052 130388
rect 110764 129844 110804 129884
rect 112492 131524 112532 131564
rect 112780 131356 112820 131396
rect 113164 131692 113204 131732
rect 113068 131608 113108 131648
rect 112492 131020 112532 131060
rect 115084 133960 115124 134000
rect 115948 133960 115988 134000
rect 114796 133372 114836 133412
rect 114412 133204 114452 133244
rect 113164 131188 113204 131228
rect 112972 130432 113012 130472
rect 112396 130180 112436 130220
rect 110572 129676 110612 129716
rect 112012 129676 112052 129716
rect 113932 129676 113972 129716
rect 123544 135304 123584 135344
rect 123626 135304 123666 135344
rect 123708 135304 123748 135344
rect 123790 135304 123830 135344
rect 123872 135304 123912 135344
rect 124784 134548 124824 134588
rect 124866 134548 124906 134588
rect 124948 134548 124988 134588
rect 125030 134548 125070 134588
rect 125112 134548 125152 134588
rect 123544 133792 123584 133832
rect 123626 133792 123666 133832
rect 123708 133792 123748 133832
rect 123790 133792 123830 133832
rect 123872 133792 123912 133832
rect 120460 133372 120500 133412
rect 120652 133372 120692 133412
rect 115180 132784 115220 132824
rect 115084 131524 115124 131564
rect 114988 131440 115028 131480
rect 114892 131188 114932 131228
rect 119308 132700 119348 132740
rect 120076 132700 120116 132740
rect 118540 132532 118580 132572
rect 118252 131272 118292 131312
rect 117580 131188 117620 131228
rect 118252 131104 118292 131144
rect 117676 130432 117716 130472
rect 115180 130348 115220 130388
rect 117484 130348 117524 130388
rect 108424 129256 108464 129296
rect 108506 129256 108546 129296
rect 108588 129256 108628 129296
rect 108670 129256 108710 129296
rect 108752 129256 108792 129296
rect 109664 128500 109704 128540
rect 109746 128500 109786 128540
rect 109828 128500 109868 128540
rect 109910 128500 109950 128540
rect 109992 128500 110032 128540
rect 120268 132532 120308 132572
rect 119116 131272 119156 131312
rect 119404 131188 119444 131228
rect 119212 130432 119252 130472
rect 119116 130348 119156 130388
rect 118540 128248 118580 128288
rect 118732 128248 118772 128288
rect 119020 128248 119060 128288
rect 108424 127744 108464 127784
rect 108506 127744 108546 127784
rect 108588 127744 108628 127784
rect 108670 127744 108710 127784
rect 108752 127744 108792 127784
rect 119116 128164 119156 128204
rect 119692 128668 119732 128708
rect 119692 128248 119732 128288
rect 118828 127912 118868 127952
rect 119596 128164 119636 128204
rect 124784 133036 124824 133076
rect 124866 133036 124906 133076
rect 124948 133036 124988 133076
rect 125030 133036 125070 133076
rect 125112 133036 125152 133076
rect 120940 132700 120980 132740
rect 121804 132700 121844 132740
rect 139904 148156 139944 148196
rect 139986 148156 140026 148196
rect 140068 148156 140108 148196
rect 140150 148156 140190 148196
rect 140232 148156 140272 148196
rect 138664 147400 138704 147440
rect 138746 147400 138786 147440
rect 138828 147400 138868 147440
rect 138910 147400 138950 147440
rect 138992 147400 139032 147440
rect 139904 146644 139944 146684
rect 139986 146644 140026 146684
rect 140068 146644 140108 146684
rect 140150 146644 140190 146684
rect 140232 146644 140272 146684
rect 138664 145888 138704 145928
rect 138746 145888 138786 145928
rect 138828 145888 138868 145928
rect 138910 145888 138950 145928
rect 138992 145888 139032 145928
rect 139904 145132 139944 145172
rect 139986 145132 140026 145172
rect 140068 145132 140108 145172
rect 140150 145132 140190 145172
rect 140232 145132 140272 145172
rect 138664 144376 138704 144416
rect 138746 144376 138786 144416
rect 138828 144376 138868 144416
rect 138910 144376 138950 144416
rect 138992 144376 139032 144416
rect 139904 143620 139944 143660
rect 139986 143620 140026 143660
rect 140068 143620 140108 143660
rect 140150 143620 140190 143660
rect 140232 143620 140272 143660
rect 138664 142864 138704 142904
rect 138746 142864 138786 142904
rect 138828 142864 138868 142904
rect 138910 142864 138950 142904
rect 138992 142864 139032 142904
rect 139904 142108 139944 142148
rect 139986 142108 140026 142148
rect 140068 142108 140108 142148
rect 140150 142108 140190 142148
rect 140232 142108 140272 142148
rect 138664 141352 138704 141392
rect 138746 141352 138786 141392
rect 138828 141352 138868 141392
rect 138910 141352 138950 141392
rect 138992 141352 139032 141392
rect 139904 140596 139944 140636
rect 139986 140596 140026 140636
rect 140068 140596 140108 140636
rect 140150 140596 140190 140636
rect 140232 140596 140272 140636
rect 138664 139840 138704 139880
rect 138746 139840 138786 139880
rect 138828 139840 138868 139880
rect 138910 139840 138950 139880
rect 138992 139840 139032 139880
rect 139904 139084 139944 139124
rect 139986 139084 140026 139124
rect 140068 139084 140108 139124
rect 140150 139084 140190 139124
rect 140232 139084 140272 139124
rect 138664 138328 138704 138368
rect 138746 138328 138786 138368
rect 138828 138328 138868 138368
rect 138910 138328 138950 138368
rect 138992 138328 139032 138368
rect 139904 137572 139944 137612
rect 139986 137572 140026 137612
rect 140068 137572 140108 137612
rect 140150 137572 140190 137612
rect 140232 137572 140272 137612
rect 138664 136816 138704 136856
rect 138746 136816 138786 136856
rect 138828 136816 138868 136856
rect 138910 136816 138950 136856
rect 138992 136816 139032 136856
rect 139904 136060 139944 136100
rect 139986 136060 140026 136100
rect 140068 136060 140108 136100
rect 140150 136060 140190 136100
rect 140232 136060 140272 136100
rect 138664 135304 138704 135344
rect 138746 135304 138786 135344
rect 138828 135304 138868 135344
rect 138910 135304 138950 135344
rect 138992 135304 139032 135344
rect 139904 134548 139944 134588
rect 139986 134548 140026 134588
rect 140068 134548 140108 134588
rect 140150 134548 140190 134588
rect 140232 134548 140272 134588
rect 151660 134044 151700 134084
rect 138664 133792 138704 133832
rect 138746 133792 138786 133832
rect 138828 133792 138868 133832
rect 138910 133792 138950 133832
rect 138992 133792 139032 133832
rect 139904 133036 139944 133076
rect 139986 133036 140026 133076
rect 140068 133036 140108 133076
rect 140150 133036 140190 133076
rect 140232 133036 140272 133076
rect 135724 132616 135764 132656
rect 123544 132280 123584 132320
rect 123626 132280 123666 132320
rect 123708 132280 123748 132320
rect 123790 132280 123830 132320
rect 123872 132280 123912 132320
rect 138664 132280 138704 132320
rect 138746 132280 138786 132320
rect 138828 132280 138868 132320
rect 138910 132280 138950 132320
rect 138992 132280 139032 132320
rect 124784 131524 124824 131564
rect 124866 131524 124906 131564
rect 124948 131524 124988 131564
rect 125030 131524 125070 131564
rect 125112 131524 125152 131564
rect 139904 131524 139944 131564
rect 139986 131524 140026 131564
rect 140068 131524 140108 131564
rect 140150 131524 140190 131564
rect 140232 131524 140272 131564
rect 123544 130768 123584 130808
rect 123626 130768 123666 130808
rect 123708 130768 123748 130808
rect 123790 130768 123830 130808
rect 123872 130768 123912 130808
rect 138664 130768 138704 130808
rect 138746 130768 138786 130808
rect 138828 130768 138868 130808
rect 138910 130768 138950 130808
rect 138992 130768 139032 130808
rect 124784 130012 124824 130052
rect 124866 130012 124906 130052
rect 124948 130012 124988 130052
rect 125030 130012 125070 130052
rect 125112 130012 125152 130052
rect 139904 130012 139944 130052
rect 139986 130012 140026 130052
rect 140068 130012 140108 130052
rect 140150 130012 140190 130052
rect 140232 130012 140272 130052
rect 123544 129256 123584 129296
rect 123626 129256 123666 129296
rect 123708 129256 123748 129296
rect 123790 129256 123830 129296
rect 123872 129256 123912 129296
rect 138664 129256 138704 129296
rect 138746 129256 138786 129296
rect 138828 129256 138868 129296
rect 138910 129256 138950 129296
rect 138992 129256 139032 129296
rect 120460 128164 120500 128204
rect 121996 128836 122036 128876
rect 123148 128836 123188 128876
rect 121900 128668 121940 128708
rect 124784 128500 124824 128540
rect 124866 128500 124906 128540
rect 124948 128500 124988 128540
rect 125030 128500 125070 128540
rect 125112 128500 125152 128540
rect 139904 128500 139944 128540
rect 139986 128500 140026 128540
rect 140068 128500 140108 128540
rect 140150 128500 140190 128540
rect 140232 128500 140272 128540
rect 121996 128164 122036 128204
rect 119212 127912 119252 127952
rect 109664 126988 109704 127028
rect 109746 126988 109786 127028
rect 109828 126988 109868 127028
rect 109910 126988 109950 127028
rect 109992 126988 110032 127028
rect 108424 126232 108464 126272
rect 108506 126232 108546 126272
rect 108588 126232 108628 126272
rect 108670 126232 108710 126272
rect 108752 126232 108792 126272
rect 109664 125476 109704 125516
rect 109746 125476 109786 125516
rect 109828 125476 109868 125516
rect 109910 125476 109950 125516
rect 109992 125476 110032 125516
rect 119980 126652 120020 126692
rect 119020 125308 119060 125348
rect 108424 124720 108464 124760
rect 108506 124720 108546 124760
rect 108588 124720 108628 124760
rect 108670 124720 108710 124760
rect 108752 124720 108792 124760
rect 109664 123964 109704 124004
rect 109746 123964 109786 124004
rect 109828 123964 109868 124004
rect 109910 123964 109950 124004
rect 109992 123964 110032 124004
rect 108424 123208 108464 123248
rect 108506 123208 108546 123248
rect 108588 123208 108628 123248
rect 108670 123208 108710 123248
rect 108752 123208 108792 123248
rect 109664 122452 109704 122492
rect 109746 122452 109786 122492
rect 109828 122452 109868 122492
rect 109910 122452 109950 122492
rect 109992 122452 110032 122492
rect 108424 121696 108464 121736
rect 108506 121696 108546 121736
rect 108588 121696 108628 121736
rect 108670 121696 108710 121736
rect 108752 121696 108792 121736
rect 109664 120940 109704 120980
rect 109746 120940 109786 120980
rect 109828 120940 109868 120980
rect 109910 120940 109950 120980
rect 109992 120940 110032 120980
rect 108424 120184 108464 120224
rect 108506 120184 108546 120224
rect 108588 120184 108628 120224
rect 108670 120184 108710 120224
rect 108752 120184 108792 120224
rect 109664 119428 109704 119468
rect 109746 119428 109786 119468
rect 109828 119428 109868 119468
rect 109910 119428 109950 119468
rect 109992 119428 110032 119468
rect 108424 118672 108464 118712
rect 108506 118672 108546 118712
rect 108588 118672 108628 118712
rect 108670 118672 108710 118712
rect 108752 118672 108792 118712
rect 109664 117916 109704 117956
rect 109746 117916 109786 117956
rect 109828 117916 109868 117956
rect 109910 117916 109950 117956
rect 109992 117916 110032 117956
rect 108424 117160 108464 117200
rect 108506 117160 108546 117200
rect 108588 117160 108628 117200
rect 108670 117160 108710 117200
rect 108752 117160 108792 117200
rect 109664 116404 109704 116444
rect 109746 116404 109786 116444
rect 109828 116404 109868 116444
rect 109910 116404 109950 116444
rect 109992 116404 110032 116444
rect 108424 115648 108464 115688
rect 108506 115648 108546 115688
rect 108588 115648 108628 115688
rect 108670 115648 108710 115688
rect 108752 115648 108792 115688
rect 109664 114892 109704 114932
rect 109746 114892 109786 114932
rect 109828 114892 109868 114932
rect 109910 114892 109950 114932
rect 109992 114892 110032 114932
rect 108424 114136 108464 114176
rect 108506 114136 108546 114176
rect 108588 114136 108628 114176
rect 108670 114136 108710 114176
rect 108752 114136 108792 114176
rect 109664 113380 109704 113420
rect 109746 113380 109786 113420
rect 109828 113380 109868 113420
rect 109910 113380 109950 113420
rect 109992 113380 110032 113420
rect 108424 112624 108464 112664
rect 108506 112624 108546 112664
rect 108588 112624 108628 112664
rect 108670 112624 108710 112664
rect 108752 112624 108792 112664
rect 109664 111868 109704 111908
rect 109746 111868 109786 111908
rect 109828 111868 109868 111908
rect 109910 111868 109950 111908
rect 109992 111868 110032 111908
rect 108424 111112 108464 111152
rect 108506 111112 108546 111152
rect 108588 111112 108628 111152
rect 108670 111112 108710 111152
rect 108752 111112 108792 111152
rect 109664 110356 109704 110396
rect 109746 110356 109786 110396
rect 109828 110356 109868 110396
rect 109910 110356 109950 110396
rect 109992 110356 110032 110396
rect 108424 109600 108464 109640
rect 108506 109600 108546 109640
rect 108588 109600 108628 109640
rect 108670 109600 108710 109640
rect 108752 109600 108792 109640
rect 109664 108844 109704 108884
rect 109746 108844 109786 108884
rect 109828 108844 109868 108884
rect 109910 108844 109950 108884
rect 109992 108844 110032 108884
rect 108424 108088 108464 108128
rect 108506 108088 108546 108128
rect 108588 108088 108628 108128
rect 108670 108088 108710 108128
rect 108752 108088 108792 108128
rect 109664 107332 109704 107372
rect 109746 107332 109786 107372
rect 109828 107332 109868 107372
rect 109910 107332 109950 107372
rect 109992 107332 110032 107372
rect 108424 106576 108464 106616
rect 108506 106576 108546 106616
rect 108588 106576 108628 106616
rect 108670 106576 108710 106616
rect 108752 106576 108792 106616
rect 109664 105820 109704 105860
rect 109746 105820 109786 105860
rect 109828 105820 109868 105860
rect 109910 105820 109950 105860
rect 109992 105820 110032 105860
rect 108424 105064 108464 105104
rect 108506 105064 108546 105104
rect 108588 105064 108628 105104
rect 108670 105064 108710 105104
rect 108752 105064 108792 105104
rect 109664 104308 109704 104348
rect 109746 104308 109786 104348
rect 109828 104308 109868 104348
rect 109910 104308 109950 104348
rect 109992 104308 110032 104348
rect 108424 103552 108464 103592
rect 108506 103552 108546 103592
rect 108588 103552 108628 103592
rect 108670 103552 108710 103592
rect 108752 103552 108792 103592
rect 109664 102796 109704 102836
rect 109746 102796 109786 102836
rect 109828 102796 109868 102836
rect 109910 102796 109950 102836
rect 109992 102796 110032 102836
rect 108424 102040 108464 102080
rect 108506 102040 108546 102080
rect 108588 102040 108628 102080
rect 108670 102040 108710 102080
rect 108752 102040 108792 102080
rect 109664 101284 109704 101324
rect 109746 101284 109786 101324
rect 109828 101284 109868 101324
rect 109910 101284 109950 101324
rect 109992 101284 110032 101324
rect 108424 100528 108464 100568
rect 108506 100528 108546 100568
rect 108588 100528 108628 100568
rect 108670 100528 108710 100568
rect 108752 100528 108792 100568
rect 109664 99772 109704 99812
rect 109746 99772 109786 99812
rect 109828 99772 109868 99812
rect 109910 99772 109950 99812
rect 109992 99772 110032 99812
rect 108424 99016 108464 99056
rect 108506 99016 108546 99056
rect 108588 99016 108628 99056
rect 108670 99016 108710 99056
rect 108752 99016 108792 99056
rect 109664 98260 109704 98300
rect 109746 98260 109786 98300
rect 109828 98260 109868 98300
rect 109910 98260 109950 98300
rect 109992 98260 110032 98300
rect 108424 97504 108464 97544
rect 108506 97504 108546 97544
rect 108588 97504 108628 97544
rect 108670 97504 108710 97544
rect 108752 97504 108792 97544
rect 109664 96748 109704 96788
rect 109746 96748 109786 96788
rect 109828 96748 109868 96788
rect 109910 96748 109950 96788
rect 109992 96748 110032 96788
rect 108424 95992 108464 96032
rect 108506 95992 108546 96032
rect 108588 95992 108628 96032
rect 108670 95992 108710 96032
rect 108752 95992 108792 96032
rect 109664 95236 109704 95276
rect 109746 95236 109786 95276
rect 109828 95236 109868 95276
rect 109910 95236 109950 95276
rect 109992 95236 110032 95276
rect 108424 94480 108464 94520
rect 108506 94480 108546 94520
rect 108588 94480 108628 94520
rect 108670 94480 108710 94520
rect 108752 94480 108792 94520
rect 109664 93724 109704 93764
rect 109746 93724 109786 93764
rect 109828 93724 109868 93764
rect 109910 93724 109950 93764
rect 109992 93724 110032 93764
rect 108424 92968 108464 93008
rect 108506 92968 108546 93008
rect 108588 92968 108628 93008
rect 108670 92968 108710 93008
rect 108752 92968 108792 93008
rect 109664 92212 109704 92252
rect 109746 92212 109786 92252
rect 109828 92212 109868 92252
rect 109910 92212 109950 92252
rect 109992 92212 110032 92252
rect 108424 91456 108464 91496
rect 108506 91456 108546 91496
rect 108588 91456 108628 91496
rect 108670 91456 108710 91496
rect 108752 91456 108792 91496
rect 109664 90700 109704 90740
rect 109746 90700 109786 90740
rect 109828 90700 109868 90740
rect 109910 90700 109950 90740
rect 109992 90700 110032 90740
rect 108424 89944 108464 89984
rect 108506 89944 108546 89984
rect 108588 89944 108628 89984
rect 108670 89944 108710 89984
rect 108752 89944 108792 89984
rect 109664 89188 109704 89228
rect 109746 89188 109786 89228
rect 109828 89188 109868 89228
rect 109910 89188 109950 89228
rect 109992 89188 110032 89228
rect 108424 88432 108464 88472
rect 108506 88432 108546 88472
rect 108588 88432 108628 88472
rect 108670 88432 108710 88472
rect 108752 88432 108792 88472
rect 109664 87676 109704 87716
rect 109746 87676 109786 87716
rect 109828 87676 109868 87716
rect 109910 87676 109950 87716
rect 109992 87676 110032 87716
rect 108424 86920 108464 86960
rect 108506 86920 108546 86960
rect 108588 86920 108628 86960
rect 108670 86920 108710 86960
rect 108752 86920 108792 86960
rect 109664 86164 109704 86204
rect 109746 86164 109786 86204
rect 109828 86164 109868 86204
rect 109910 86164 109950 86204
rect 109992 86164 110032 86204
rect 108424 85408 108464 85448
rect 108506 85408 108546 85448
rect 108588 85408 108628 85448
rect 108670 85408 108710 85448
rect 108752 85408 108792 85448
rect 109664 84652 109704 84692
rect 109746 84652 109786 84692
rect 109828 84652 109868 84692
rect 109910 84652 109950 84692
rect 109992 84652 110032 84692
rect 108424 83896 108464 83936
rect 108506 83896 108546 83936
rect 108588 83896 108628 83936
rect 108670 83896 108710 83936
rect 108752 83896 108792 83936
rect 109664 83140 109704 83180
rect 109746 83140 109786 83180
rect 109828 83140 109868 83180
rect 109910 83140 109950 83180
rect 109992 83140 110032 83180
rect 108424 82384 108464 82424
rect 108506 82384 108546 82424
rect 108588 82384 108628 82424
rect 108670 82384 108710 82424
rect 108752 82384 108792 82424
rect 109664 81628 109704 81668
rect 109746 81628 109786 81668
rect 109828 81628 109868 81668
rect 109910 81628 109950 81668
rect 109992 81628 110032 81668
rect 108424 80872 108464 80912
rect 108506 80872 108546 80912
rect 108588 80872 108628 80912
rect 108670 80872 108710 80912
rect 108752 80872 108792 80912
rect 109664 80116 109704 80156
rect 109746 80116 109786 80156
rect 109828 80116 109868 80156
rect 109910 80116 109950 80156
rect 109992 80116 110032 80156
rect 108424 79360 108464 79400
rect 108506 79360 108546 79400
rect 108588 79360 108628 79400
rect 108670 79360 108710 79400
rect 108752 79360 108792 79400
rect 109664 78604 109704 78644
rect 109746 78604 109786 78644
rect 109828 78604 109868 78644
rect 109910 78604 109950 78644
rect 109992 78604 110032 78644
rect 108424 77848 108464 77888
rect 108506 77848 108546 77888
rect 108588 77848 108628 77888
rect 108670 77848 108710 77888
rect 108752 77848 108792 77888
rect 109664 77092 109704 77132
rect 109746 77092 109786 77132
rect 109828 77092 109868 77132
rect 109910 77092 109950 77132
rect 109992 77092 110032 77132
rect 108424 76336 108464 76376
rect 108506 76336 108546 76376
rect 108588 76336 108628 76376
rect 108670 76336 108710 76376
rect 108752 76336 108792 76376
rect 109664 75580 109704 75620
rect 109746 75580 109786 75620
rect 109828 75580 109868 75620
rect 109910 75580 109950 75620
rect 109992 75580 110032 75620
rect 121036 125308 121076 125348
rect 123544 127744 123584 127784
rect 123626 127744 123666 127784
rect 123708 127744 123748 127784
rect 123790 127744 123830 127784
rect 123872 127744 123912 127784
rect 138664 127744 138704 127784
rect 138746 127744 138786 127784
rect 138828 127744 138868 127784
rect 138910 127744 138950 127784
rect 138992 127744 139032 127784
rect 124784 126988 124824 127028
rect 124866 126988 124906 127028
rect 124948 126988 124988 127028
rect 125030 126988 125070 127028
rect 125112 126988 125152 127028
rect 139904 126988 139944 127028
rect 139986 126988 140026 127028
rect 140068 126988 140108 127028
rect 140150 126988 140190 127028
rect 140232 126988 140272 127028
rect 123544 126232 123584 126272
rect 123626 126232 123666 126272
rect 123708 126232 123748 126272
rect 123790 126232 123830 126272
rect 123872 126232 123912 126272
rect 138664 126232 138704 126272
rect 138746 126232 138786 126272
rect 138828 126232 138868 126272
rect 138910 126232 138950 126272
rect 138992 126232 139032 126272
rect 124784 125476 124824 125516
rect 124866 125476 124906 125516
rect 124948 125476 124988 125516
rect 125030 125476 125070 125516
rect 125112 125476 125152 125516
rect 139904 125476 139944 125516
rect 139986 125476 140026 125516
rect 140068 125476 140108 125516
rect 140150 125476 140190 125516
rect 140232 125476 140272 125516
rect 123544 124720 123584 124760
rect 123626 124720 123666 124760
rect 123708 124720 123748 124760
rect 123790 124720 123830 124760
rect 123872 124720 123912 124760
rect 138664 124720 138704 124760
rect 138746 124720 138786 124760
rect 138828 124720 138868 124760
rect 138910 124720 138950 124760
rect 138992 124720 139032 124760
rect 124784 123964 124824 124004
rect 124866 123964 124906 124004
rect 124948 123964 124988 124004
rect 125030 123964 125070 124004
rect 125112 123964 125152 124004
rect 139904 123964 139944 124004
rect 139986 123964 140026 124004
rect 140068 123964 140108 124004
rect 140150 123964 140190 124004
rect 140232 123964 140272 124004
rect 123544 123208 123584 123248
rect 123626 123208 123666 123248
rect 123708 123208 123748 123248
rect 123790 123208 123830 123248
rect 123872 123208 123912 123248
rect 138664 123208 138704 123248
rect 138746 123208 138786 123248
rect 138828 123208 138868 123248
rect 138910 123208 138950 123248
rect 138992 123208 139032 123248
rect 124784 122452 124824 122492
rect 124866 122452 124906 122492
rect 124948 122452 124988 122492
rect 125030 122452 125070 122492
rect 125112 122452 125152 122492
rect 139904 122452 139944 122492
rect 139986 122452 140026 122492
rect 140068 122452 140108 122492
rect 140150 122452 140190 122492
rect 140232 122452 140272 122492
rect 123544 121696 123584 121736
rect 123626 121696 123666 121736
rect 123708 121696 123748 121736
rect 123790 121696 123830 121736
rect 123872 121696 123912 121736
rect 138664 121696 138704 121736
rect 138746 121696 138786 121736
rect 138828 121696 138868 121736
rect 138910 121696 138950 121736
rect 138992 121696 139032 121736
rect 124784 120940 124824 120980
rect 124866 120940 124906 120980
rect 124948 120940 124988 120980
rect 125030 120940 125070 120980
rect 125112 120940 125152 120980
rect 139904 120940 139944 120980
rect 139986 120940 140026 120980
rect 140068 120940 140108 120980
rect 140150 120940 140190 120980
rect 140232 120940 140272 120980
rect 123544 120184 123584 120224
rect 123626 120184 123666 120224
rect 123708 120184 123748 120224
rect 123790 120184 123830 120224
rect 123872 120184 123912 120224
rect 138664 120184 138704 120224
rect 138746 120184 138786 120224
rect 138828 120184 138868 120224
rect 138910 120184 138950 120224
rect 138992 120184 139032 120224
rect 123148 119596 123188 119636
rect 124784 119428 124824 119468
rect 124866 119428 124906 119468
rect 124948 119428 124988 119468
rect 125030 119428 125070 119468
rect 125112 119428 125152 119468
rect 139904 119428 139944 119468
rect 139986 119428 140026 119468
rect 140068 119428 140108 119468
rect 140150 119428 140190 119468
rect 140232 119428 140272 119468
rect 123544 118672 123584 118712
rect 123626 118672 123666 118712
rect 123708 118672 123748 118712
rect 123790 118672 123830 118712
rect 123872 118672 123912 118712
rect 138664 118672 138704 118712
rect 138746 118672 138786 118712
rect 138828 118672 138868 118712
rect 138910 118672 138950 118712
rect 138992 118672 139032 118712
rect 124784 117916 124824 117956
rect 124866 117916 124906 117956
rect 124948 117916 124988 117956
rect 125030 117916 125070 117956
rect 125112 117916 125152 117956
rect 139904 117916 139944 117956
rect 139986 117916 140026 117956
rect 140068 117916 140108 117956
rect 140150 117916 140190 117956
rect 140232 117916 140272 117956
rect 123544 117160 123584 117200
rect 123626 117160 123666 117200
rect 123708 117160 123748 117200
rect 123790 117160 123830 117200
rect 123872 117160 123912 117200
rect 138664 117160 138704 117200
rect 138746 117160 138786 117200
rect 138828 117160 138868 117200
rect 138910 117160 138950 117200
rect 138992 117160 139032 117200
rect 124784 116404 124824 116444
rect 124866 116404 124906 116444
rect 124948 116404 124988 116444
rect 125030 116404 125070 116444
rect 125112 116404 125152 116444
rect 139904 116404 139944 116444
rect 139986 116404 140026 116444
rect 140068 116404 140108 116444
rect 140150 116404 140190 116444
rect 140232 116404 140272 116444
rect 123544 115648 123584 115688
rect 123626 115648 123666 115688
rect 123708 115648 123748 115688
rect 123790 115648 123830 115688
rect 123872 115648 123912 115688
rect 138664 115648 138704 115688
rect 138746 115648 138786 115688
rect 138828 115648 138868 115688
rect 138910 115648 138950 115688
rect 138992 115648 139032 115688
rect 124784 114892 124824 114932
rect 124866 114892 124906 114932
rect 124948 114892 124988 114932
rect 125030 114892 125070 114932
rect 125112 114892 125152 114932
rect 139904 114892 139944 114932
rect 139986 114892 140026 114932
rect 140068 114892 140108 114932
rect 140150 114892 140190 114932
rect 140232 114892 140272 114932
rect 123544 114136 123584 114176
rect 123626 114136 123666 114176
rect 123708 114136 123748 114176
rect 123790 114136 123830 114176
rect 123872 114136 123912 114176
rect 138664 114136 138704 114176
rect 138746 114136 138786 114176
rect 138828 114136 138868 114176
rect 138910 114136 138950 114176
rect 138992 114136 139032 114176
rect 124784 113380 124824 113420
rect 124866 113380 124906 113420
rect 124948 113380 124988 113420
rect 125030 113380 125070 113420
rect 125112 113380 125152 113420
rect 139904 113380 139944 113420
rect 139986 113380 140026 113420
rect 140068 113380 140108 113420
rect 140150 113380 140190 113420
rect 140232 113380 140272 113420
rect 123544 112624 123584 112664
rect 123626 112624 123666 112664
rect 123708 112624 123748 112664
rect 123790 112624 123830 112664
rect 123872 112624 123912 112664
rect 138664 112624 138704 112664
rect 138746 112624 138786 112664
rect 138828 112624 138868 112664
rect 138910 112624 138950 112664
rect 138992 112624 139032 112664
rect 124784 111868 124824 111908
rect 124866 111868 124906 111908
rect 124948 111868 124988 111908
rect 125030 111868 125070 111908
rect 125112 111868 125152 111908
rect 139904 111868 139944 111908
rect 139986 111868 140026 111908
rect 140068 111868 140108 111908
rect 140150 111868 140190 111908
rect 140232 111868 140272 111908
rect 123544 111112 123584 111152
rect 123626 111112 123666 111152
rect 123708 111112 123748 111152
rect 123790 111112 123830 111152
rect 123872 111112 123912 111152
rect 138664 111112 138704 111152
rect 138746 111112 138786 111152
rect 138828 111112 138868 111152
rect 138910 111112 138950 111152
rect 138992 111112 139032 111152
rect 124784 110356 124824 110396
rect 124866 110356 124906 110396
rect 124948 110356 124988 110396
rect 125030 110356 125070 110396
rect 125112 110356 125152 110396
rect 139904 110356 139944 110396
rect 139986 110356 140026 110396
rect 140068 110356 140108 110396
rect 140150 110356 140190 110396
rect 140232 110356 140272 110396
rect 123544 109600 123584 109640
rect 123626 109600 123666 109640
rect 123708 109600 123748 109640
rect 123790 109600 123830 109640
rect 123872 109600 123912 109640
rect 138664 109600 138704 109640
rect 138746 109600 138786 109640
rect 138828 109600 138868 109640
rect 138910 109600 138950 109640
rect 138992 109600 139032 109640
rect 124784 108844 124824 108884
rect 124866 108844 124906 108884
rect 124948 108844 124988 108884
rect 125030 108844 125070 108884
rect 125112 108844 125152 108884
rect 139904 108844 139944 108884
rect 139986 108844 140026 108884
rect 140068 108844 140108 108884
rect 140150 108844 140190 108884
rect 140232 108844 140272 108884
rect 123544 108088 123584 108128
rect 123626 108088 123666 108128
rect 123708 108088 123748 108128
rect 123790 108088 123830 108128
rect 123872 108088 123912 108128
rect 138664 108088 138704 108128
rect 138746 108088 138786 108128
rect 138828 108088 138868 108128
rect 138910 108088 138950 108128
rect 138992 108088 139032 108128
rect 124784 107332 124824 107372
rect 124866 107332 124906 107372
rect 124948 107332 124988 107372
rect 125030 107332 125070 107372
rect 125112 107332 125152 107372
rect 139904 107332 139944 107372
rect 139986 107332 140026 107372
rect 140068 107332 140108 107372
rect 140150 107332 140190 107372
rect 140232 107332 140272 107372
rect 123544 106576 123584 106616
rect 123626 106576 123666 106616
rect 123708 106576 123748 106616
rect 123790 106576 123830 106616
rect 123872 106576 123912 106616
rect 138664 106576 138704 106616
rect 138746 106576 138786 106616
rect 138828 106576 138868 106616
rect 138910 106576 138950 106616
rect 138992 106576 139032 106616
rect 124784 105820 124824 105860
rect 124866 105820 124906 105860
rect 124948 105820 124988 105860
rect 125030 105820 125070 105860
rect 125112 105820 125152 105860
rect 139904 105820 139944 105860
rect 139986 105820 140026 105860
rect 140068 105820 140108 105860
rect 140150 105820 140190 105860
rect 140232 105820 140272 105860
rect 123544 105064 123584 105104
rect 123626 105064 123666 105104
rect 123708 105064 123748 105104
rect 123790 105064 123830 105104
rect 123872 105064 123912 105104
rect 138664 105064 138704 105104
rect 138746 105064 138786 105104
rect 138828 105064 138868 105104
rect 138910 105064 138950 105104
rect 138992 105064 139032 105104
rect 124784 104308 124824 104348
rect 124866 104308 124906 104348
rect 124948 104308 124988 104348
rect 125030 104308 125070 104348
rect 125112 104308 125152 104348
rect 139904 104308 139944 104348
rect 139986 104308 140026 104348
rect 140068 104308 140108 104348
rect 140150 104308 140190 104348
rect 140232 104308 140272 104348
rect 121612 103720 121652 103760
rect 123544 103552 123584 103592
rect 123626 103552 123666 103592
rect 123708 103552 123748 103592
rect 123790 103552 123830 103592
rect 123872 103552 123912 103592
rect 138664 103552 138704 103592
rect 138746 103552 138786 103592
rect 138828 103552 138868 103592
rect 138910 103552 138950 103592
rect 138992 103552 139032 103592
rect 124784 102796 124824 102836
rect 124866 102796 124906 102836
rect 124948 102796 124988 102836
rect 125030 102796 125070 102836
rect 125112 102796 125152 102836
rect 139904 102796 139944 102836
rect 139986 102796 140026 102836
rect 140068 102796 140108 102836
rect 140150 102796 140190 102836
rect 140232 102796 140272 102836
rect 123544 102040 123584 102080
rect 123626 102040 123666 102080
rect 123708 102040 123748 102080
rect 123790 102040 123830 102080
rect 123872 102040 123912 102080
rect 138664 102040 138704 102080
rect 138746 102040 138786 102080
rect 138828 102040 138868 102080
rect 138910 102040 138950 102080
rect 138992 102040 139032 102080
rect 124784 101284 124824 101324
rect 124866 101284 124906 101324
rect 124948 101284 124988 101324
rect 125030 101284 125070 101324
rect 125112 101284 125152 101324
rect 139904 101284 139944 101324
rect 139986 101284 140026 101324
rect 140068 101284 140108 101324
rect 140150 101284 140190 101324
rect 140232 101284 140272 101324
rect 123544 100528 123584 100568
rect 123626 100528 123666 100568
rect 123708 100528 123748 100568
rect 123790 100528 123830 100568
rect 123872 100528 123912 100568
rect 138664 100528 138704 100568
rect 138746 100528 138786 100568
rect 138828 100528 138868 100568
rect 138910 100528 138950 100568
rect 138992 100528 139032 100568
rect 124784 99772 124824 99812
rect 124866 99772 124906 99812
rect 124948 99772 124988 99812
rect 125030 99772 125070 99812
rect 125112 99772 125152 99812
rect 139904 99772 139944 99812
rect 139986 99772 140026 99812
rect 140068 99772 140108 99812
rect 140150 99772 140190 99812
rect 140232 99772 140272 99812
rect 123544 99016 123584 99056
rect 123626 99016 123666 99056
rect 123708 99016 123748 99056
rect 123790 99016 123830 99056
rect 123872 99016 123912 99056
rect 138664 99016 138704 99056
rect 138746 99016 138786 99056
rect 138828 99016 138868 99056
rect 138910 99016 138950 99056
rect 138992 99016 139032 99056
rect 124784 98260 124824 98300
rect 124866 98260 124906 98300
rect 124948 98260 124988 98300
rect 125030 98260 125070 98300
rect 125112 98260 125152 98300
rect 139904 98260 139944 98300
rect 139986 98260 140026 98300
rect 140068 98260 140108 98300
rect 140150 98260 140190 98300
rect 140232 98260 140272 98300
rect 123544 97504 123584 97544
rect 123626 97504 123666 97544
rect 123708 97504 123748 97544
rect 123790 97504 123830 97544
rect 123872 97504 123912 97544
rect 138664 97504 138704 97544
rect 138746 97504 138786 97544
rect 138828 97504 138868 97544
rect 138910 97504 138950 97544
rect 138992 97504 139032 97544
rect 124784 96748 124824 96788
rect 124866 96748 124906 96788
rect 124948 96748 124988 96788
rect 125030 96748 125070 96788
rect 125112 96748 125152 96788
rect 139904 96748 139944 96788
rect 139986 96748 140026 96788
rect 140068 96748 140108 96788
rect 140150 96748 140190 96788
rect 140232 96748 140272 96788
rect 123544 95992 123584 96032
rect 123626 95992 123666 96032
rect 123708 95992 123748 96032
rect 123790 95992 123830 96032
rect 123872 95992 123912 96032
rect 138664 95992 138704 96032
rect 138746 95992 138786 96032
rect 138828 95992 138868 96032
rect 138910 95992 138950 96032
rect 138992 95992 139032 96032
rect 124784 95236 124824 95276
rect 124866 95236 124906 95276
rect 124948 95236 124988 95276
rect 125030 95236 125070 95276
rect 125112 95236 125152 95276
rect 139904 95236 139944 95276
rect 139986 95236 140026 95276
rect 140068 95236 140108 95276
rect 140150 95236 140190 95276
rect 140232 95236 140272 95276
rect 123544 94480 123584 94520
rect 123626 94480 123666 94520
rect 123708 94480 123748 94520
rect 123790 94480 123830 94520
rect 123872 94480 123912 94520
rect 138664 94480 138704 94520
rect 138746 94480 138786 94520
rect 138828 94480 138868 94520
rect 138910 94480 138950 94520
rect 138992 94480 139032 94520
rect 124784 93724 124824 93764
rect 124866 93724 124906 93764
rect 124948 93724 124988 93764
rect 125030 93724 125070 93764
rect 125112 93724 125152 93764
rect 139904 93724 139944 93764
rect 139986 93724 140026 93764
rect 140068 93724 140108 93764
rect 140150 93724 140190 93764
rect 140232 93724 140272 93764
rect 123544 92968 123584 93008
rect 123626 92968 123666 93008
rect 123708 92968 123748 93008
rect 123790 92968 123830 93008
rect 123872 92968 123912 93008
rect 138664 92968 138704 93008
rect 138746 92968 138786 93008
rect 138828 92968 138868 93008
rect 138910 92968 138950 93008
rect 138992 92968 139032 93008
rect 124784 92212 124824 92252
rect 124866 92212 124906 92252
rect 124948 92212 124988 92252
rect 125030 92212 125070 92252
rect 125112 92212 125152 92252
rect 139904 92212 139944 92252
rect 139986 92212 140026 92252
rect 140068 92212 140108 92252
rect 140150 92212 140190 92252
rect 140232 92212 140272 92252
rect 123544 91456 123584 91496
rect 123626 91456 123666 91496
rect 123708 91456 123748 91496
rect 123790 91456 123830 91496
rect 123872 91456 123912 91496
rect 138664 91456 138704 91496
rect 138746 91456 138786 91496
rect 138828 91456 138868 91496
rect 138910 91456 138950 91496
rect 138992 91456 139032 91496
rect 124784 90700 124824 90740
rect 124866 90700 124906 90740
rect 124948 90700 124988 90740
rect 125030 90700 125070 90740
rect 125112 90700 125152 90740
rect 139904 90700 139944 90740
rect 139986 90700 140026 90740
rect 140068 90700 140108 90740
rect 140150 90700 140190 90740
rect 140232 90700 140272 90740
rect 123544 89944 123584 89984
rect 123626 89944 123666 89984
rect 123708 89944 123748 89984
rect 123790 89944 123830 89984
rect 123872 89944 123912 89984
rect 138664 89944 138704 89984
rect 138746 89944 138786 89984
rect 138828 89944 138868 89984
rect 138910 89944 138950 89984
rect 138992 89944 139032 89984
rect 124784 89188 124824 89228
rect 124866 89188 124906 89228
rect 124948 89188 124988 89228
rect 125030 89188 125070 89228
rect 125112 89188 125152 89228
rect 139904 89188 139944 89228
rect 139986 89188 140026 89228
rect 140068 89188 140108 89228
rect 140150 89188 140190 89228
rect 140232 89188 140272 89228
rect 123544 88432 123584 88472
rect 123626 88432 123666 88472
rect 123708 88432 123748 88472
rect 123790 88432 123830 88472
rect 123872 88432 123912 88472
rect 138664 88432 138704 88472
rect 138746 88432 138786 88472
rect 138828 88432 138868 88472
rect 138910 88432 138950 88472
rect 138992 88432 139032 88472
rect 148204 87844 148244 87884
rect 124784 87676 124824 87716
rect 124866 87676 124906 87716
rect 124948 87676 124988 87716
rect 125030 87676 125070 87716
rect 125112 87676 125152 87716
rect 139904 87676 139944 87716
rect 139986 87676 140026 87716
rect 140068 87676 140108 87716
rect 140150 87676 140190 87716
rect 140232 87676 140272 87716
rect 123544 86920 123584 86960
rect 123626 86920 123666 86960
rect 123708 86920 123748 86960
rect 123790 86920 123830 86960
rect 123872 86920 123912 86960
rect 138664 86920 138704 86960
rect 138746 86920 138786 86960
rect 138828 86920 138868 86960
rect 138910 86920 138950 86960
rect 138992 86920 139032 86960
rect 124784 86164 124824 86204
rect 124866 86164 124906 86204
rect 124948 86164 124988 86204
rect 125030 86164 125070 86204
rect 125112 86164 125152 86204
rect 139904 86164 139944 86204
rect 139986 86164 140026 86204
rect 140068 86164 140108 86204
rect 140150 86164 140190 86204
rect 140232 86164 140272 86204
rect 123544 85408 123584 85448
rect 123626 85408 123666 85448
rect 123708 85408 123748 85448
rect 123790 85408 123830 85448
rect 123872 85408 123912 85448
rect 138664 85408 138704 85448
rect 138746 85408 138786 85448
rect 138828 85408 138868 85448
rect 138910 85408 138950 85448
rect 138992 85408 139032 85448
rect 124784 84652 124824 84692
rect 124866 84652 124906 84692
rect 124948 84652 124988 84692
rect 125030 84652 125070 84692
rect 125112 84652 125152 84692
rect 139904 84652 139944 84692
rect 139986 84652 140026 84692
rect 140068 84652 140108 84692
rect 140150 84652 140190 84692
rect 140232 84652 140272 84692
rect 123544 83896 123584 83936
rect 123626 83896 123666 83936
rect 123708 83896 123748 83936
rect 123790 83896 123830 83936
rect 123872 83896 123912 83936
rect 138664 83896 138704 83936
rect 138746 83896 138786 83936
rect 138828 83896 138868 83936
rect 138910 83896 138950 83936
rect 138992 83896 139032 83936
rect 124784 83140 124824 83180
rect 124866 83140 124906 83180
rect 124948 83140 124988 83180
rect 125030 83140 125070 83180
rect 125112 83140 125152 83180
rect 139904 83140 139944 83180
rect 139986 83140 140026 83180
rect 140068 83140 140108 83180
rect 140150 83140 140190 83180
rect 140232 83140 140272 83180
rect 123544 82384 123584 82424
rect 123626 82384 123666 82424
rect 123708 82384 123748 82424
rect 123790 82384 123830 82424
rect 123872 82384 123912 82424
rect 138664 82384 138704 82424
rect 138746 82384 138786 82424
rect 138828 82384 138868 82424
rect 138910 82384 138950 82424
rect 138992 82384 139032 82424
rect 124784 81628 124824 81668
rect 124866 81628 124906 81668
rect 124948 81628 124988 81668
rect 125030 81628 125070 81668
rect 125112 81628 125152 81668
rect 139904 81628 139944 81668
rect 139986 81628 140026 81668
rect 140068 81628 140108 81668
rect 140150 81628 140190 81668
rect 140232 81628 140272 81668
rect 123544 80872 123584 80912
rect 123626 80872 123666 80912
rect 123708 80872 123748 80912
rect 123790 80872 123830 80912
rect 123872 80872 123912 80912
rect 138664 80872 138704 80912
rect 138746 80872 138786 80912
rect 138828 80872 138868 80912
rect 138910 80872 138950 80912
rect 138992 80872 139032 80912
rect 124784 80116 124824 80156
rect 124866 80116 124906 80156
rect 124948 80116 124988 80156
rect 125030 80116 125070 80156
rect 125112 80116 125152 80156
rect 139904 80116 139944 80156
rect 139986 80116 140026 80156
rect 140068 80116 140108 80156
rect 140150 80116 140190 80156
rect 140232 80116 140272 80156
rect 123544 79360 123584 79400
rect 123626 79360 123666 79400
rect 123708 79360 123748 79400
rect 123790 79360 123830 79400
rect 123872 79360 123912 79400
rect 138664 79360 138704 79400
rect 138746 79360 138786 79400
rect 138828 79360 138868 79400
rect 138910 79360 138950 79400
rect 138992 79360 139032 79400
rect 124784 78604 124824 78644
rect 124866 78604 124906 78644
rect 124948 78604 124988 78644
rect 125030 78604 125070 78644
rect 125112 78604 125152 78644
rect 139904 78604 139944 78644
rect 139986 78604 140026 78644
rect 140068 78604 140108 78644
rect 140150 78604 140190 78644
rect 140232 78604 140272 78644
rect 123544 77848 123584 77888
rect 123626 77848 123666 77888
rect 123708 77848 123748 77888
rect 123790 77848 123830 77888
rect 123872 77848 123912 77888
rect 138664 77848 138704 77888
rect 138746 77848 138786 77888
rect 138828 77848 138868 77888
rect 138910 77848 138950 77888
rect 138992 77848 139032 77888
rect 124784 77092 124824 77132
rect 124866 77092 124906 77132
rect 124948 77092 124988 77132
rect 125030 77092 125070 77132
rect 125112 77092 125152 77132
rect 139904 77092 139944 77132
rect 139986 77092 140026 77132
rect 140068 77092 140108 77132
rect 140150 77092 140190 77132
rect 140232 77092 140272 77132
rect 123544 76336 123584 76376
rect 123626 76336 123666 76376
rect 123708 76336 123748 76376
rect 123790 76336 123830 76376
rect 123872 76336 123912 76376
rect 138664 76336 138704 76376
rect 138746 76336 138786 76376
rect 138828 76336 138868 76376
rect 138910 76336 138950 76376
rect 138992 76336 139032 76376
rect 124784 75580 124824 75620
rect 124866 75580 124906 75620
rect 124948 75580 124988 75620
rect 125030 75580 125070 75620
rect 125112 75580 125152 75620
rect 139904 75580 139944 75620
rect 139986 75580 140026 75620
rect 140068 75580 140108 75620
rect 140150 75580 140190 75620
rect 140232 75580 140272 75620
rect 148204 72388 148244 72428
rect 73324 64156 73364 64196
<< metal3 >>
rect 119692 159704 119732 160029
rect 112291 159664 112300 159704
rect 112340 159664 119732 159704
rect 64099 152020 64108 152060
rect 64148 152020 94060 152060
rect 94100 152020 94109 152060
rect 160012 151640 160052 151704
rect 115939 151600 115948 151640
rect 115988 151600 160052 151640
rect 79415 148156 79424 148196
rect 79464 148156 79506 148196
rect 79546 148156 79588 148196
rect 79628 148156 79670 148196
rect 79710 148156 79752 148196
rect 79792 148156 79801 148196
rect 94535 148156 94544 148196
rect 94584 148156 94626 148196
rect 94666 148156 94708 148196
rect 94748 148156 94790 148196
rect 94830 148156 94872 148196
rect 94912 148156 94921 148196
rect 109655 148156 109664 148196
rect 109704 148156 109746 148196
rect 109786 148156 109828 148196
rect 109868 148156 109910 148196
rect 109950 148156 109992 148196
rect 110032 148156 110041 148196
rect 124775 148156 124784 148196
rect 124824 148156 124866 148196
rect 124906 148156 124948 148196
rect 124988 148156 125030 148196
rect 125070 148156 125112 148196
rect 125152 148156 125161 148196
rect 139895 148156 139904 148196
rect 139944 148156 139986 148196
rect 140026 148156 140068 148196
rect 140108 148156 140150 148196
rect 140190 148156 140232 148196
rect 140272 148156 140281 148196
rect 78175 147400 78184 147440
rect 78224 147400 78266 147440
rect 78306 147400 78348 147440
rect 78388 147400 78430 147440
rect 78470 147400 78512 147440
rect 78552 147400 78561 147440
rect 93295 147400 93304 147440
rect 93344 147400 93386 147440
rect 93426 147400 93468 147440
rect 93508 147400 93550 147440
rect 93590 147400 93632 147440
rect 93672 147400 93681 147440
rect 108415 147400 108424 147440
rect 108464 147400 108506 147440
rect 108546 147400 108588 147440
rect 108628 147400 108670 147440
rect 108710 147400 108752 147440
rect 108792 147400 108801 147440
rect 123535 147400 123544 147440
rect 123584 147400 123626 147440
rect 123666 147400 123708 147440
rect 123748 147400 123790 147440
rect 123830 147400 123872 147440
rect 123912 147400 123921 147440
rect 138655 147400 138664 147440
rect 138704 147400 138746 147440
rect 138786 147400 138828 147440
rect 138868 147400 138910 147440
rect 138950 147400 138992 147440
rect 139032 147400 139041 147440
rect 79415 146644 79424 146684
rect 79464 146644 79506 146684
rect 79546 146644 79588 146684
rect 79628 146644 79670 146684
rect 79710 146644 79752 146684
rect 79792 146644 79801 146684
rect 94535 146644 94544 146684
rect 94584 146644 94626 146684
rect 94666 146644 94708 146684
rect 94748 146644 94790 146684
rect 94830 146644 94872 146684
rect 94912 146644 94921 146684
rect 109655 146644 109664 146684
rect 109704 146644 109746 146684
rect 109786 146644 109828 146684
rect 109868 146644 109910 146684
rect 109950 146644 109992 146684
rect 110032 146644 110041 146684
rect 124775 146644 124784 146684
rect 124824 146644 124866 146684
rect 124906 146644 124948 146684
rect 124988 146644 125030 146684
rect 125070 146644 125112 146684
rect 125152 146644 125161 146684
rect 139895 146644 139904 146684
rect 139944 146644 139986 146684
rect 140026 146644 140068 146684
rect 140108 146644 140150 146684
rect 140190 146644 140232 146684
rect 140272 146644 140281 146684
rect 78175 145888 78184 145928
rect 78224 145888 78266 145928
rect 78306 145888 78348 145928
rect 78388 145888 78430 145928
rect 78470 145888 78512 145928
rect 78552 145888 78561 145928
rect 93295 145888 93304 145928
rect 93344 145888 93386 145928
rect 93426 145888 93468 145928
rect 93508 145888 93550 145928
rect 93590 145888 93632 145928
rect 93672 145888 93681 145928
rect 108415 145888 108424 145928
rect 108464 145888 108506 145928
rect 108546 145888 108588 145928
rect 108628 145888 108670 145928
rect 108710 145888 108752 145928
rect 108792 145888 108801 145928
rect 123535 145888 123544 145928
rect 123584 145888 123626 145928
rect 123666 145888 123708 145928
rect 123748 145888 123790 145928
rect 123830 145888 123872 145928
rect 123912 145888 123921 145928
rect 138655 145888 138664 145928
rect 138704 145888 138746 145928
rect 138786 145888 138828 145928
rect 138868 145888 138910 145928
rect 138950 145888 138992 145928
rect 139032 145888 139041 145928
rect 79415 145132 79424 145172
rect 79464 145132 79506 145172
rect 79546 145132 79588 145172
rect 79628 145132 79670 145172
rect 79710 145132 79752 145172
rect 79792 145132 79801 145172
rect 94535 145132 94544 145172
rect 94584 145132 94626 145172
rect 94666 145132 94708 145172
rect 94748 145132 94790 145172
rect 94830 145132 94872 145172
rect 94912 145132 94921 145172
rect 109655 145132 109664 145172
rect 109704 145132 109746 145172
rect 109786 145132 109828 145172
rect 109868 145132 109910 145172
rect 109950 145132 109992 145172
rect 110032 145132 110041 145172
rect 124775 145132 124784 145172
rect 124824 145132 124866 145172
rect 124906 145132 124948 145172
rect 124988 145132 125030 145172
rect 125070 145132 125112 145172
rect 125152 145132 125161 145172
rect 139895 145132 139904 145172
rect 139944 145132 139986 145172
rect 140026 145132 140068 145172
rect 140108 145132 140150 145172
rect 140190 145132 140232 145172
rect 140272 145132 140281 145172
rect 78175 144376 78184 144416
rect 78224 144376 78266 144416
rect 78306 144376 78348 144416
rect 78388 144376 78430 144416
rect 78470 144376 78512 144416
rect 78552 144376 78561 144416
rect 93295 144376 93304 144416
rect 93344 144376 93386 144416
rect 93426 144376 93468 144416
rect 93508 144376 93550 144416
rect 93590 144376 93632 144416
rect 93672 144376 93681 144416
rect 108415 144376 108424 144416
rect 108464 144376 108506 144416
rect 108546 144376 108588 144416
rect 108628 144376 108670 144416
rect 108710 144376 108752 144416
rect 108792 144376 108801 144416
rect 123535 144376 123544 144416
rect 123584 144376 123626 144416
rect 123666 144376 123708 144416
rect 123748 144376 123790 144416
rect 123830 144376 123872 144416
rect 123912 144376 123921 144416
rect 138655 144376 138664 144416
rect 138704 144376 138746 144416
rect 138786 144376 138828 144416
rect 138868 144376 138910 144416
rect 138950 144376 138992 144416
rect 139032 144376 139041 144416
rect 79415 143620 79424 143660
rect 79464 143620 79506 143660
rect 79546 143620 79588 143660
rect 79628 143620 79670 143660
rect 79710 143620 79752 143660
rect 79792 143620 79801 143660
rect 94535 143620 94544 143660
rect 94584 143620 94626 143660
rect 94666 143620 94708 143660
rect 94748 143620 94790 143660
rect 94830 143620 94872 143660
rect 94912 143620 94921 143660
rect 109655 143620 109664 143660
rect 109704 143620 109746 143660
rect 109786 143620 109828 143660
rect 109868 143620 109910 143660
rect 109950 143620 109992 143660
rect 110032 143620 110041 143660
rect 124775 143620 124784 143660
rect 124824 143620 124866 143660
rect 124906 143620 124948 143660
rect 124988 143620 125030 143660
rect 125070 143620 125112 143660
rect 125152 143620 125161 143660
rect 139895 143620 139904 143660
rect 139944 143620 139986 143660
rect 140026 143620 140068 143660
rect 140108 143620 140150 143660
rect 140190 143620 140232 143660
rect 140272 143620 140281 143660
rect 78175 142864 78184 142904
rect 78224 142864 78266 142904
rect 78306 142864 78348 142904
rect 78388 142864 78430 142904
rect 78470 142864 78512 142904
rect 78552 142864 78561 142904
rect 93295 142864 93304 142904
rect 93344 142864 93386 142904
rect 93426 142864 93468 142904
rect 93508 142864 93550 142904
rect 93590 142864 93632 142904
rect 93672 142864 93681 142904
rect 108415 142864 108424 142904
rect 108464 142864 108506 142904
rect 108546 142864 108588 142904
rect 108628 142864 108670 142904
rect 108710 142864 108752 142904
rect 108792 142864 108801 142904
rect 123535 142864 123544 142904
rect 123584 142864 123626 142904
rect 123666 142864 123708 142904
rect 123748 142864 123790 142904
rect 123830 142864 123872 142904
rect 123912 142864 123921 142904
rect 138655 142864 138664 142904
rect 138704 142864 138746 142904
rect 138786 142864 138828 142904
rect 138868 142864 138910 142904
rect 138950 142864 138992 142904
rect 139032 142864 139041 142904
rect 79415 142108 79424 142148
rect 79464 142108 79506 142148
rect 79546 142108 79588 142148
rect 79628 142108 79670 142148
rect 79710 142108 79752 142148
rect 79792 142108 79801 142148
rect 94535 142108 94544 142148
rect 94584 142108 94626 142148
rect 94666 142108 94708 142148
rect 94748 142108 94790 142148
rect 94830 142108 94872 142148
rect 94912 142108 94921 142148
rect 109655 142108 109664 142148
rect 109704 142108 109746 142148
rect 109786 142108 109828 142148
rect 109868 142108 109910 142148
rect 109950 142108 109992 142148
rect 110032 142108 110041 142148
rect 124775 142108 124784 142148
rect 124824 142108 124866 142148
rect 124906 142108 124948 142148
rect 124988 142108 125030 142148
rect 125070 142108 125112 142148
rect 125152 142108 125161 142148
rect 139895 142108 139904 142148
rect 139944 142108 139986 142148
rect 140026 142108 140068 142148
rect 140108 142108 140150 142148
rect 140190 142108 140232 142148
rect 140272 142108 140281 142148
rect 78175 141352 78184 141392
rect 78224 141352 78266 141392
rect 78306 141352 78348 141392
rect 78388 141352 78430 141392
rect 78470 141352 78512 141392
rect 78552 141352 78561 141392
rect 93295 141352 93304 141392
rect 93344 141352 93386 141392
rect 93426 141352 93468 141392
rect 93508 141352 93550 141392
rect 93590 141352 93632 141392
rect 93672 141352 93681 141392
rect 108415 141352 108424 141392
rect 108464 141352 108506 141392
rect 108546 141352 108588 141392
rect 108628 141352 108670 141392
rect 108710 141352 108752 141392
rect 108792 141352 108801 141392
rect 123535 141352 123544 141392
rect 123584 141352 123626 141392
rect 123666 141352 123708 141392
rect 123748 141352 123790 141392
rect 123830 141352 123872 141392
rect 123912 141352 123921 141392
rect 138655 141352 138664 141392
rect 138704 141352 138746 141392
rect 138786 141352 138828 141392
rect 138868 141352 138910 141392
rect 138950 141352 138992 141392
rect 139032 141352 139041 141392
rect 79415 140596 79424 140636
rect 79464 140596 79506 140636
rect 79546 140596 79588 140636
rect 79628 140596 79670 140636
rect 79710 140596 79752 140636
rect 79792 140596 79801 140636
rect 94535 140596 94544 140636
rect 94584 140596 94626 140636
rect 94666 140596 94708 140636
rect 94748 140596 94790 140636
rect 94830 140596 94872 140636
rect 94912 140596 94921 140636
rect 109655 140596 109664 140636
rect 109704 140596 109746 140636
rect 109786 140596 109828 140636
rect 109868 140596 109910 140636
rect 109950 140596 109992 140636
rect 110032 140596 110041 140636
rect 124775 140596 124784 140636
rect 124824 140596 124866 140636
rect 124906 140596 124948 140636
rect 124988 140596 125030 140636
rect 125070 140596 125112 140636
rect 125152 140596 125161 140636
rect 139895 140596 139904 140636
rect 139944 140596 139986 140636
rect 140026 140596 140068 140636
rect 140108 140596 140150 140636
rect 140190 140596 140232 140636
rect 140272 140596 140281 140636
rect 78175 139840 78184 139880
rect 78224 139840 78266 139880
rect 78306 139840 78348 139880
rect 78388 139840 78430 139880
rect 78470 139840 78512 139880
rect 78552 139840 78561 139880
rect 93295 139840 93304 139880
rect 93344 139840 93386 139880
rect 93426 139840 93468 139880
rect 93508 139840 93550 139880
rect 93590 139840 93632 139880
rect 93672 139840 93681 139880
rect 108415 139840 108424 139880
rect 108464 139840 108506 139880
rect 108546 139840 108588 139880
rect 108628 139840 108670 139880
rect 108710 139840 108752 139880
rect 108792 139840 108801 139880
rect 123535 139840 123544 139880
rect 123584 139840 123626 139880
rect 123666 139840 123708 139880
rect 123748 139840 123790 139880
rect 123830 139840 123872 139880
rect 123912 139840 123921 139880
rect 138655 139840 138664 139880
rect 138704 139840 138746 139880
rect 138786 139840 138828 139880
rect 138868 139840 138910 139880
rect 138950 139840 138992 139880
rect 139032 139840 139041 139880
rect 79415 139084 79424 139124
rect 79464 139084 79506 139124
rect 79546 139084 79588 139124
rect 79628 139084 79670 139124
rect 79710 139084 79752 139124
rect 79792 139084 79801 139124
rect 94535 139084 94544 139124
rect 94584 139084 94626 139124
rect 94666 139084 94708 139124
rect 94748 139084 94790 139124
rect 94830 139084 94872 139124
rect 94912 139084 94921 139124
rect 109655 139084 109664 139124
rect 109704 139084 109746 139124
rect 109786 139084 109828 139124
rect 109868 139084 109910 139124
rect 109950 139084 109992 139124
rect 110032 139084 110041 139124
rect 124775 139084 124784 139124
rect 124824 139084 124866 139124
rect 124906 139084 124948 139124
rect 124988 139084 125030 139124
rect 125070 139084 125112 139124
rect 125152 139084 125161 139124
rect 139895 139084 139904 139124
rect 139944 139084 139986 139124
rect 140026 139084 140068 139124
rect 140108 139084 140150 139124
rect 140190 139084 140232 139124
rect 140272 139084 140281 139124
rect 78175 138328 78184 138368
rect 78224 138328 78266 138368
rect 78306 138328 78348 138368
rect 78388 138328 78430 138368
rect 78470 138328 78512 138368
rect 78552 138328 78561 138368
rect 93295 138328 93304 138368
rect 93344 138328 93386 138368
rect 93426 138328 93468 138368
rect 93508 138328 93550 138368
rect 93590 138328 93632 138368
rect 93672 138328 93681 138368
rect 108415 138328 108424 138368
rect 108464 138328 108506 138368
rect 108546 138328 108588 138368
rect 108628 138328 108670 138368
rect 108710 138328 108752 138368
rect 108792 138328 108801 138368
rect 123535 138328 123544 138368
rect 123584 138328 123626 138368
rect 123666 138328 123708 138368
rect 123748 138328 123790 138368
rect 123830 138328 123872 138368
rect 123912 138328 123921 138368
rect 138655 138328 138664 138368
rect 138704 138328 138746 138368
rect 138786 138328 138828 138368
rect 138868 138328 138910 138368
rect 138950 138328 138992 138368
rect 139032 138328 139041 138368
rect 79415 137572 79424 137612
rect 79464 137572 79506 137612
rect 79546 137572 79588 137612
rect 79628 137572 79670 137612
rect 79710 137572 79752 137612
rect 79792 137572 79801 137612
rect 94535 137572 94544 137612
rect 94584 137572 94626 137612
rect 94666 137572 94708 137612
rect 94748 137572 94790 137612
rect 94830 137572 94872 137612
rect 94912 137572 94921 137612
rect 109655 137572 109664 137612
rect 109704 137572 109746 137612
rect 109786 137572 109828 137612
rect 109868 137572 109910 137612
rect 109950 137572 109992 137612
rect 110032 137572 110041 137612
rect 124775 137572 124784 137612
rect 124824 137572 124866 137612
rect 124906 137572 124948 137612
rect 124988 137572 125030 137612
rect 125070 137572 125112 137612
rect 125152 137572 125161 137612
rect 139895 137572 139904 137612
rect 139944 137572 139986 137612
rect 140026 137572 140068 137612
rect 140108 137572 140150 137612
rect 140190 137572 140232 137612
rect 140272 137572 140281 137612
rect 78175 136816 78184 136856
rect 78224 136816 78266 136856
rect 78306 136816 78348 136856
rect 78388 136816 78430 136856
rect 78470 136816 78512 136856
rect 78552 136816 78561 136856
rect 93295 136816 93304 136856
rect 93344 136816 93386 136856
rect 93426 136816 93468 136856
rect 93508 136816 93550 136856
rect 93590 136816 93632 136856
rect 93672 136816 93681 136856
rect 108415 136816 108424 136856
rect 108464 136816 108506 136856
rect 108546 136816 108588 136856
rect 108628 136816 108670 136856
rect 108710 136816 108752 136856
rect 108792 136816 108801 136856
rect 123535 136816 123544 136856
rect 123584 136816 123626 136856
rect 123666 136816 123708 136856
rect 123748 136816 123790 136856
rect 123830 136816 123872 136856
rect 123912 136816 123921 136856
rect 138655 136816 138664 136856
rect 138704 136816 138746 136856
rect 138786 136816 138828 136856
rect 138868 136816 138910 136856
rect 138950 136816 138992 136856
rect 139032 136816 139041 136856
rect 79415 136060 79424 136100
rect 79464 136060 79506 136100
rect 79546 136060 79588 136100
rect 79628 136060 79670 136100
rect 79710 136060 79752 136100
rect 79792 136060 79801 136100
rect 94535 136060 94544 136100
rect 94584 136060 94626 136100
rect 94666 136060 94708 136100
rect 94748 136060 94790 136100
rect 94830 136060 94872 136100
rect 94912 136060 94921 136100
rect 109655 136060 109664 136100
rect 109704 136060 109746 136100
rect 109786 136060 109828 136100
rect 109868 136060 109910 136100
rect 109950 136060 109992 136100
rect 110032 136060 110041 136100
rect 124775 136060 124784 136100
rect 124824 136060 124866 136100
rect 124906 136060 124948 136100
rect 124988 136060 125030 136100
rect 125070 136060 125112 136100
rect 125152 136060 125161 136100
rect 139895 136060 139904 136100
rect 139944 136060 139986 136100
rect 140026 136060 140068 136100
rect 140108 136060 140150 136100
rect 140190 136060 140232 136100
rect 140272 136060 140281 136100
rect 148300 135640 160032 135680
rect 148300 135596 148340 135640
rect 121795 135556 121804 135596
rect 121844 135556 148340 135596
rect 67660 135472 78604 135512
rect 78644 135472 78653 135512
rect 67660 135428 67700 135472
rect 64099 135388 64108 135428
rect 64148 135388 67700 135428
rect 78175 135304 78184 135344
rect 78224 135304 78266 135344
rect 78306 135304 78348 135344
rect 78388 135304 78430 135344
rect 78470 135304 78512 135344
rect 78552 135304 78561 135344
rect 93295 135304 93304 135344
rect 93344 135304 93386 135344
rect 93426 135304 93468 135344
rect 93508 135304 93550 135344
rect 93590 135304 93632 135344
rect 93672 135304 93681 135344
rect 108415 135304 108424 135344
rect 108464 135304 108506 135344
rect 108546 135304 108588 135344
rect 108628 135304 108670 135344
rect 108710 135304 108752 135344
rect 108792 135304 108801 135344
rect 123535 135304 123544 135344
rect 123584 135304 123626 135344
rect 123666 135304 123708 135344
rect 123748 135304 123790 135344
rect 123830 135304 123872 135344
rect 123912 135304 123921 135344
rect 138655 135304 138664 135344
rect 138704 135304 138746 135344
rect 138786 135304 138828 135344
rect 138868 135304 138910 135344
rect 138950 135304 138992 135344
rect 139032 135304 139041 135344
rect 79415 134548 79424 134588
rect 79464 134548 79506 134588
rect 79546 134548 79588 134588
rect 79628 134548 79670 134588
rect 79710 134548 79752 134588
rect 79792 134548 79801 134588
rect 94535 134548 94544 134588
rect 94584 134548 94626 134588
rect 94666 134548 94708 134588
rect 94748 134548 94790 134588
rect 94830 134548 94872 134588
rect 94912 134548 94921 134588
rect 109655 134548 109664 134588
rect 109704 134548 109746 134588
rect 109786 134548 109828 134588
rect 109868 134548 109910 134588
rect 109950 134548 109992 134588
rect 110032 134548 110041 134588
rect 124775 134548 124784 134588
rect 124824 134548 124866 134588
rect 124906 134548 124948 134588
rect 124988 134548 125030 134588
rect 125070 134548 125112 134588
rect 125152 134548 125161 134588
rect 139895 134548 139904 134588
rect 139944 134548 139986 134588
rect 140026 134548 140068 134588
rect 140108 134548 140150 134588
rect 140190 134548 140232 134588
rect 140272 134548 140281 134588
rect 97411 134212 97420 134252
rect 97460 134212 98188 134252
rect 98228 134212 98237 134252
rect 98659 134212 98668 134252
rect 98708 134212 105100 134252
rect 105140 134212 105149 134252
rect 99811 134044 99820 134084
rect 99860 134044 100012 134084
rect 100052 134044 151660 134084
rect 151700 134044 151709 134084
rect 115075 133960 115084 134000
rect 115124 133960 115948 134000
rect 115988 133960 115997 134000
rect 78175 133792 78184 133832
rect 78224 133792 78266 133832
rect 78306 133792 78348 133832
rect 78388 133792 78430 133832
rect 78470 133792 78512 133832
rect 78552 133792 78561 133832
rect 93295 133792 93304 133832
rect 93344 133792 93386 133832
rect 93426 133792 93468 133832
rect 93508 133792 93550 133832
rect 93590 133792 93632 133832
rect 93672 133792 93681 133832
rect 108415 133792 108424 133832
rect 108464 133792 108506 133832
rect 108546 133792 108588 133832
rect 108628 133792 108670 133832
rect 108710 133792 108752 133832
rect 108792 133792 108801 133832
rect 123535 133792 123544 133832
rect 123584 133792 123626 133832
rect 123666 133792 123708 133832
rect 123748 133792 123790 133832
rect 123830 133792 123872 133832
rect 123912 133792 123921 133832
rect 138655 133792 138664 133832
rect 138704 133792 138746 133832
rect 138786 133792 138828 133832
rect 138868 133792 138910 133832
rect 138950 133792 138992 133832
rect 139032 133792 139041 133832
rect 114787 133372 114796 133412
rect 114836 133372 120460 133412
rect 120500 133372 120652 133412
rect 120692 133372 120701 133412
rect 112867 133204 112876 133244
rect 112916 133204 114412 133244
rect 114452 133204 114461 133244
rect 79415 133036 79424 133076
rect 79464 133036 79506 133076
rect 79546 133036 79588 133076
rect 79628 133036 79670 133076
rect 79710 133036 79752 133076
rect 79792 133036 79801 133076
rect 94535 133036 94544 133076
rect 94584 133036 94626 133076
rect 94666 133036 94708 133076
rect 94748 133036 94790 133076
rect 94830 133036 94872 133076
rect 94912 133036 94921 133076
rect 109655 133036 109664 133076
rect 109704 133036 109746 133076
rect 109786 133036 109828 133076
rect 109868 133036 109910 133076
rect 109950 133036 109992 133076
rect 110032 133036 110041 133076
rect 124775 133036 124784 133076
rect 124824 133036 124866 133076
rect 124906 133036 124948 133076
rect 124988 133036 125030 133076
rect 125070 133036 125112 133076
rect 125152 133036 125161 133076
rect 139895 133036 139904 133076
rect 139944 133036 139986 133076
rect 140026 133036 140068 133076
rect 140108 133036 140150 133076
rect 140190 133036 140232 133076
rect 140272 133036 140281 133076
rect 115171 132784 115180 132824
rect 115220 132784 120980 132824
rect 120940 132740 120980 132784
rect 98755 132700 98764 132740
rect 98804 132700 100012 132740
rect 100052 132700 100061 132740
rect 102211 132700 102220 132740
rect 102260 132700 102988 132740
rect 103028 132700 103037 132740
rect 119299 132700 119308 132740
rect 119348 132700 120076 132740
rect 120116 132700 120125 132740
rect 120931 132700 120940 132740
rect 120980 132700 121804 132740
rect 121844 132700 121853 132740
rect 101347 132616 101356 132656
rect 101396 132616 106252 132656
rect 106292 132616 135724 132656
rect 135764 132616 135773 132656
rect 79267 132532 79276 132572
rect 79316 132532 94252 132572
rect 94292 132532 94301 132572
rect 118531 132532 118540 132572
rect 118580 132532 120268 132572
rect 120308 132532 120317 132572
rect 78175 132280 78184 132320
rect 78224 132280 78266 132320
rect 78306 132280 78348 132320
rect 78388 132280 78430 132320
rect 78470 132280 78512 132320
rect 78552 132280 78561 132320
rect 93295 132280 93304 132320
rect 93344 132280 93386 132320
rect 93426 132280 93468 132320
rect 93508 132280 93550 132320
rect 93590 132280 93632 132320
rect 93672 132280 93681 132320
rect 108415 132280 108424 132320
rect 108464 132280 108506 132320
rect 108546 132280 108588 132320
rect 108628 132280 108670 132320
rect 108710 132280 108752 132320
rect 108792 132280 108801 132320
rect 123535 132280 123544 132320
rect 123584 132280 123626 132320
rect 123666 132280 123708 132320
rect 123748 132280 123790 132320
rect 123830 132280 123872 132320
rect 123912 132280 123921 132320
rect 138655 132280 138664 132320
rect 138704 132280 138746 132320
rect 138786 132280 138828 132320
rect 138868 132280 138910 132320
rect 138950 132280 138992 132320
rect 139032 132280 139041 132320
rect 98851 132028 98860 132068
rect 98900 132028 99052 132068
rect 99092 132028 99436 132068
rect 99476 132028 101068 132068
rect 101108 132028 101117 132068
rect 99523 131944 99532 131984
rect 99572 131944 100012 131984
rect 100052 131944 101164 131984
rect 101204 131944 101213 131984
rect 100195 131860 100204 131900
rect 100244 131860 101356 131900
rect 101396 131860 101405 131900
rect 110755 131776 110764 131816
rect 110804 131776 112396 131816
rect 112436 131776 112445 131816
rect 99235 131692 99244 131732
rect 99284 131692 101548 131732
rect 101588 131692 101597 131732
rect 112579 131692 112588 131732
rect 112628 131692 113164 131732
rect 113204 131692 113213 131732
rect 108739 131608 108748 131648
rect 108788 131608 113068 131648
rect 113108 131608 113117 131648
rect 79415 131524 79424 131564
rect 79464 131524 79506 131564
rect 79546 131524 79588 131564
rect 79628 131524 79670 131564
rect 79710 131524 79752 131564
rect 79792 131524 79801 131564
rect 94535 131524 94544 131564
rect 94584 131524 94626 131564
rect 94666 131524 94708 131564
rect 94748 131524 94790 131564
rect 94830 131524 94872 131564
rect 94912 131524 94921 131564
rect 109655 131524 109664 131564
rect 109704 131524 109746 131564
rect 109786 131524 109828 131564
rect 109868 131524 109910 131564
rect 109950 131524 109992 131564
rect 110032 131524 110041 131564
rect 112483 131524 112492 131564
rect 112532 131524 115084 131564
rect 115124 131524 115133 131564
rect 124775 131524 124784 131564
rect 124824 131524 124866 131564
rect 124906 131524 124948 131564
rect 124988 131524 125030 131564
rect 125070 131524 125112 131564
rect 125152 131524 125161 131564
rect 139895 131524 139904 131564
rect 139944 131524 139986 131564
rect 140026 131524 140068 131564
rect 140108 131524 140150 131564
rect 140190 131524 140232 131564
rect 140272 131524 140281 131564
rect 103939 131440 103948 131480
rect 103988 131440 111436 131480
rect 111476 131440 111820 131480
rect 111860 131440 114988 131480
rect 115028 131440 115037 131480
rect 109411 131356 109420 131396
rect 109460 131356 109804 131396
rect 109844 131356 109853 131396
rect 110371 131356 110380 131396
rect 110420 131356 110764 131396
rect 110804 131356 110813 131396
rect 112291 131356 112300 131396
rect 112340 131356 112780 131396
rect 112820 131356 112829 131396
rect 101251 131272 101260 131312
rect 101300 131272 102124 131312
rect 102164 131272 102173 131312
rect 109036 131272 114932 131312
rect 118243 131272 118252 131312
rect 118292 131272 119116 131312
rect 119156 131272 119165 131312
rect 109036 131228 109076 131272
rect 114892 131228 114932 131272
rect 100579 131188 100588 131228
rect 100628 131188 102028 131228
rect 102068 131188 102077 131228
rect 103459 131188 103468 131228
rect 103508 131188 109036 131228
rect 109076 131188 109085 131228
rect 109411 131188 109420 131228
rect 109460 131188 110476 131228
rect 110516 131188 110525 131228
rect 113155 131188 113164 131228
rect 113204 131188 113213 131228
rect 114883 131188 114892 131228
rect 114932 131188 114941 131228
rect 117571 131188 117580 131228
rect 117620 131188 119404 131228
rect 119444 131188 119453 131228
rect 113164 131144 113204 131188
rect 102220 131104 104332 131144
rect 104372 131104 108748 131144
rect 108788 131104 108940 131144
rect 108980 131104 108989 131144
rect 109123 131104 109132 131144
rect 109172 131104 110380 131144
rect 110420 131104 110429 131144
rect 113164 131104 118252 131144
rect 118292 131104 118301 131144
rect 102220 131060 102260 131104
rect 99331 131020 99340 131060
rect 99380 131020 102220 131060
rect 102260 131020 102269 131060
rect 103555 131020 103564 131060
rect 103604 131020 104044 131060
rect 104084 131020 104093 131060
rect 109603 131020 109612 131060
rect 109652 131020 110572 131060
rect 110612 131020 112492 131060
rect 112532 131020 112541 131060
rect 110755 130936 110764 130976
rect 110804 130936 112204 130976
rect 112244 130936 112253 130976
rect 78175 130768 78184 130808
rect 78224 130768 78266 130808
rect 78306 130768 78348 130808
rect 78388 130768 78430 130808
rect 78470 130768 78512 130808
rect 78552 130768 78561 130808
rect 93295 130768 93304 130808
rect 93344 130768 93386 130808
rect 93426 130768 93468 130808
rect 93508 130768 93550 130808
rect 93590 130768 93632 130808
rect 93672 130768 93681 130808
rect 108415 130768 108424 130808
rect 108464 130768 108506 130808
rect 108546 130768 108588 130808
rect 108628 130768 108670 130808
rect 108710 130768 108752 130808
rect 108792 130768 108801 130808
rect 123535 130768 123544 130808
rect 123584 130768 123626 130808
rect 123666 130768 123708 130808
rect 123748 130768 123790 130808
rect 123830 130768 123872 130808
rect 123912 130768 123921 130808
rect 138655 130768 138664 130808
rect 138704 130768 138746 130808
rect 138786 130768 138828 130808
rect 138868 130768 138910 130808
rect 138950 130768 138992 130808
rect 139032 130768 139041 130808
rect 105091 130684 105100 130724
rect 105140 130684 108020 130724
rect 107980 130640 108020 130684
rect 107980 130600 108748 130640
rect 108788 130600 110668 130640
rect 110708 130600 110717 130640
rect 112963 130432 112972 130472
rect 113012 130432 117676 130472
rect 117716 130432 119212 130472
rect 119252 130432 119261 130472
rect 96835 130348 96844 130388
rect 96884 130348 98092 130388
rect 98132 130348 99052 130388
rect 99092 130348 99101 130388
rect 101635 130348 101644 130388
rect 101684 130348 105388 130388
rect 105428 130348 105964 130388
rect 106004 130348 106013 130388
rect 110179 130348 110188 130388
rect 110228 130348 112012 130388
rect 112052 130348 112061 130388
rect 115171 130348 115180 130388
rect 115220 130348 117484 130388
rect 117524 130348 119116 130388
rect 119156 130348 119165 130388
rect 99139 130264 99148 130304
rect 99188 130264 103084 130304
rect 103124 130264 103468 130304
rect 103508 130264 103517 130304
rect 103267 130180 103276 130220
rect 103316 130180 104716 130220
rect 104756 130180 104765 130220
rect 105955 130180 105964 130220
rect 106004 130180 110668 130220
rect 110708 130180 112396 130220
rect 112436 130180 112445 130220
rect 97219 130096 97228 130136
rect 97268 130096 99916 130136
rect 99956 130096 99965 130136
rect 79415 130012 79424 130052
rect 79464 130012 79506 130052
rect 79546 130012 79588 130052
rect 79628 130012 79670 130052
rect 79710 130012 79752 130052
rect 79792 130012 79801 130052
rect 94535 130012 94544 130052
rect 94584 130012 94626 130052
rect 94666 130012 94708 130052
rect 94748 130012 94790 130052
rect 94830 130012 94872 130052
rect 94912 130012 94921 130052
rect 109655 130012 109664 130052
rect 109704 130012 109746 130052
rect 109786 130012 109828 130052
rect 109868 130012 109910 130052
rect 109950 130012 109992 130052
rect 110032 130012 110041 130052
rect 124775 130012 124784 130052
rect 124824 130012 124866 130052
rect 124906 130012 124948 130052
rect 124988 130012 125030 130052
rect 125070 130012 125112 130052
rect 125152 130012 125161 130052
rect 139895 130012 139904 130052
rect 139944 130012 139986 130052
rect 140026 130012 140068 130052
rect 140108 130012 140150 130052
rect 140190 130012 140232 130052
rect 140272 130012 140281 130052
rect 95011 129928 95020 129968
rect 95060 129928 97132 129968
rect 97172 129928 97181 129968
rect 99907 129928 99916 129968
rect 99956 129928 103124 129968
rect 103084 129884 103124 129928
rect 94147 129844 94156 129884
rect 94196 129844 96172 129884
rect 96212 129844 96221 129884
rect 97411 129844 97420 129884
rect 97460 129844 98956 129884
rect 98996 129844 100108 129884
rect 100148 129844 100157 129884
rect 103075 129844 103084 129884
rect 103124 129844 110764 129884
rect 110804 129844 110813 129884
rect 73315 129676 73324 129716
rect 73364 129676 110572 129716
rect 110612 129676 110621 129716
rect 112003 129676 112012 129716
rect 112052 129676 113932 129716
rect 113972 129676 113981 129716
rect 78175 129256 78184 129296
rect 78224 129256 78266 129296
rect 78306 129256 78348 129296
rect 78388 129256 78430 129296
rect 78470 129256 78512 129296
rect 78552 129256 78561 129296
rect 93295 129256 93304 129296
rect 93344 129256 93386 129296
rect 93426 129256 93468 129296
rect 93508 129256 93550 129296
rect 93590 129256 93632 129296
rect 93672 129256 93681 129296
rect 108415 129256 108424 129296
rect 108464 129256 108506 129296
rect 108546 129256 108588 129296
rect 108628 129256 108670 129296
rect 108710 129256 108752 129296
rect 108792 129256 108801 129296
rect 123535 129256 123544 129296
rect 123584 129256 123626 129296
rect 123666 129256 123708 129296
rect 123748 129256 123790 129296
rect 123830 129256 123872 129296
rect 123912 129256 123921 129296
rect 138655 129256 138664 129296
rect 138704 129256 138746 129296
rect 138786 129256 138828 129296
rect 138868 129256 138910 129296
rect 138950 129256 138992 129296
rect 139032 129256 139041 129296
rect 121987 128836 121996 128876
rect 122036 128836 123148 128876
rect 123188 128836 123197 128876
rect 119683 128668 119692 128708
rect 119732 128668 121900 128708
rect 121940 128668 121949 128708
rect 79415 128500 79424 128540
rect 79464 128500 79506 128540
rect 79546 128500 79588 128540
rect 79628 128500 79670 128540
rect 79710 128500 79752 128540
rect 79792 128500 79801 128540
rect 94535 128500 94544 128540
rect 94584 128500 94626 128540
rect 94666 128500 94708 128540
rect 94748 128500 94790 128540
rect 94830 128500 94872 128540
rect 94912 128500 94921 128540
rect 109655 128500 109664 128540
rect 109704 128500 109746 128540
rect 109786 128500 109828 128540
rect 109868 128500 109910 128540
rect 109950 128500 109992 128540
rect 110032 128500 110041 128540
rect 124775 128500 124784 128540
rect 124824 128500 124866 128540
rect 124906 128500 124948 128540
rect 124988 128500 125030 128540
rect 125070 128500 125112 128540
rect 125152 128500 125161 128540
rect 139895 128500 139904 128540
rect 139944 128500 139986 128540
rect 140026 128500 140068 128540
rect 140108 128500 140150 128540
rect 140190 128500 140232 128540
rect 140272 128500 140281 128540
rect 94819 128332 94828 128372
rect 94868 128332 96076 128372
rect 96116 128332 96125 128372
rect 95491 128248 95500 128288
rect 95540 128248 97996 128288
rect 98036 128248 99188 128288
rect 118531 128248 118540 128288
rect 118580 128248 118732 128288
rect 118772 128248 119020 128288
rect 119060 128248 119692 128288
rect 119732 128248 119741 128288
rect 99148 128180 99188 128248
rect 99139 128140 99148 128180
rect 99188 128140 99197 128180
rect 119107 128164 119116 128204
rect 119156 128164 119596 128204
rect 119636 128164 119645 128204
rect 120451 128164 120460 128204
rect 120500 128164 121996 128204
rect 122036 128164 122045 128204
rect 118819 127912 118828 127952
rect 118868 127912 119212 127952
rect 119252 127912 119261 127952
rect 78175 127744 78184 127784
rect 78224 127744 78266 127784
rect 78306 127744 78348 127784
rect 78388 127744 78430 127784
rect 78470 127744 78512 127784
rect 78552 127744 78561 127784
rect 93295 127744 93304 127784
rect 93344 127744 93386 127784
rect 93426 127744 93468 127784
rect 93508 127744 93550 127784
rect 93590 127744 93632 127784
rect 93672 127744 93681 127784
rect 108415 127744 108424 127784
rect 108464 127744 108506 127784
rect 108546 127744 108588 127784
rect 108628 127744 108670 127784
rect 108710 127744 108752 127784
rect 108792 127744 108801 127784
rect 123535 127744 123544 127784
rect 123584 127744 123626 127784
rect 123666 127744 123708 127784
rect 123748 127744 123790 127784
rect 123830 127744 123872 127784
rect 123912 127744 123921 127784
rect 138655 127744 138664 127784
rect 138704 127744 138746 127784
rect 138786 127744 138828 127784
rect 138868 127744 138910 127784
rect 138950 127744 138992 127784
rect 139032 127744 139041 127784
rect 87820 127324 94732 127364
rect 94772 127324 94781 127364
rect 87820 127280 87860 127324
rect 79843 127240 79852 127280
rect 79892 127240 87860 127280
rect 79415 126988 79424 127028
rect 79464 126988 79506 127028
rect 79546 126988 79588 127028
rect 79628 126988 79670 127028
rect 79710 126988 79752 127028
rect 79792 126988 79801 127028
rect 94535 126988 94544 127028
rect 94584 126988 94626 127028
rect 94666 126988 94708 127028
rect 94748 126988 94790 127028
rect 94830 126988 94872 127028
rect 94912 126988 94921 127028
rect 109655 126988 109664 127028
rect 109704 126988 109746 127028
rect 109786 126988 109828 127028
rect 109868 126988 109910 127028
rect 109950 126988 109992 127028
rect 110032 126988 110041 127028
rect 124775 126988 124784 127028
rect 124824 126988 124866 127028
rect 124906 126988 124948 127028
rect 124988 126988 125030 127028
rect 125070 126988 125112 127028
rect 125152 126988 125161 127028
rect 139895 126988 139904 127028
rect 139944 126988 139986 127028
rect 140026 126988 140068 127028
rect 140108 126988 140150 127028
rect 140190 126988 140232 127028
rect 140272 126988 140281 127028
rect 94051 126820 94060 126860
rect 94100 126820 94636 126860
rect 94676 126820 94685 126860
rect 93955 126736 93964 126776
rect 94004 126736 94732 126776
rect 94772 126736 94781 126776
rect 94915 126652 94924 126692
rect 94964 126652 95884 126692
rect 95924 126652 119980 126692
rect 120020 126652 120029 126692
rect 93763 126568 93772 126608
rect 93812 126568 94828 126608
rect 94868 126568 94877 126608
rect 95011 126568 95020 126608
rect 95060 126568 95788 126608
rect 95828 126568 104044 126608
rect 104084 126568 104093 126608
rect 94828 126524 94868 126568
rect 94828 126484 95596 126524
rect 95636 126484 95645 126524
rect 94243 126400 94252 126440
rect 94292 126400 95692 126440
rect 95732 126400 95741 126440
rect 78175 126232 78184 126272
rect 78224 126232 78266 126272
rect 78306 126232 78348 126272
rect 78388 126232 78430 126272
rect 78470 126232 78512 126272
rect 78552 126232 78561 126272
rect 93295 126232 93304 126272
rect 93344 126232 93386 126272
rect 93426 126232 93468 126272
rect 93508 126232 93550 126272
rect 93590 126232 93632 126272
rect 93672 126232 93681 126272
rect 108415 126232 108424 126272
rect 108464 126232 108506 126272
rect 108546 126232 108588 126272
rect 108628 126232 108670 126272
rect 108710 126232 108752 126272
rect 108792 126232 108801 126272
rect 123535 126232 123544 126272
rect 123584 126232 123626 126272
rect 123666 126232 123708 126272
rect 123748 126232 123790 126272
rect 123830 126232 123872 126272
rect 123912 126232 123921 126272
rect 138655 126232 138664 126272
rect 138704 126232 138746 126272
rect 138786 126232 138828 126272
rect 138868 126232 138910 126272
rect 138950 126232 138992 126272
rect 139032 126232 139041 126272
rect 79415 125476 79424 125516
rect 79464 125476 79506 125516
rect 79546 125476 79588 125516
rect 79628 125476 79670 125516
rect 79710 125476 79752 125516
rect 79792 125476 79801 125516
rect 94535 125476 94544 125516
rect 94584 125476 94626 125516
rect 94666 125476 94708 125516
rect 94748 125476 94790 125516
rect 94830 125476 94872 125516
rect 94912 125476 94921 125516
rect 109655 125476 109664 125516
rect 109704 125476 109746 125516
rect 109786 125476 109828 125516
rect 109868 125476 109910 125516
rect 109950 125476 109992 125516
rect 110032 125476 110041 125516
rect 124775 125476 124784 125516
rect 124824 125476 124866 125516
rect 124906 125476 124948 125516
rect 124988 125476 125030 125516
rect 125070 125476 125112 125516
rect 125152 125476 125161 125516
rect 139895 125476 139904 125516
rect 139944 125476 139986 125516
rect 140026 125476 140068 125516
rect 140108 125476 140150 125516
rect 140190 125476 140232 125516
rect 140272 125476 140281 125516
rect 119011 125308 119020 125348
rect 119060 125308 121036 125348
rect 121076 125308 121085 125348
rect 93763 125264 93821 125265
rect 93678 125224 93772 125264
rect 93812 125224 93821 125264
rect 93763 125223 93821 125224
rect 78175 124720 78184 124760
rect 78224 124720 78266 124760
rect 78306 124720 78348 124760
rect 78388 124720 78430 124760
rect 78470 124720 78512 124760
rect 78552 124720 78561 124760
rect 93295 124720 93304 124760
rect 93344 124720 93386 124760
rect 93426 124720 93468 124760
rect 93508 124720 93550 124760
rect 93590 124720 93632 124760
rect 93672 124720 93681 124760
rect 108415 124720 108424 124760
rect 108464 124720 108506 124760
rect 108546 124720 108588 124760
rect 108628 124720 108670 124760
rect 108710 124720 108752 124760
rect 108792 124720 108801 124760
rect 123535 124720 123544 124760
rect 123584 124720 123626 124760
rect 123666 124720 123708 124760
rect 123748 124720 123790 124760
rect 123830 124720 123872 124760
rect 123912 124720 123921 124760
rect 138655 124720 138664 124760
rect 138704 124720 138746 124760
rect 138786 124720 138828 124760
rect 138868 124720 138910 124760
rect 138950 124720 138992 124760
rect 139032 124720 139041 124760
rect 78883 124300 78892 124340
rect 78932 124300 93868 124340
rect 93908 124300 93917 124340
rect 79415 123964 79424 124004
rect 79464 123964 79506 124004
rect 79546 123964 79588 124004
rect 79628 123964 79670 124004
rect 79710 123964 79752 124004
rect 79792 123964 79801 124004
rect 94535 123964 94544 124004
rect 94584 123964 94626 124004
rect 94666 123964 94708 124004
rect 94748 123964 94790 124004
rect 94830 123964 94872 124004
rect 94912 123964 94921 124004
rect 109655 123964 109664 124004
rect 109704 123964 109746 124004
rect 109786 123964 109828 124004
rect 109868 123964 109910 124004
rect 109950 123964 109992 124004
rect 110032 123964 110041 124004
rect 124775 123964 124784 124004
rect 124824 123964 124866 124004
rect 124906 123964 124948 124004
rect 124988 123964 125030 124004
rect 125070 123964 125112 124004
rect 125152 123964 125161 124004
rect 139895 123964 139904 124004
rect 139944 123964 139986 124004
rect 140026 123964 140068 124004
rect 140108 123964 140150 124004
rect 140190 123964 140232 124004
rect 140272 123964 140281 124004
rect 78175 123208 78184 123248
rect 78224 123208 78266 123248
rect 78306 123208 78348 123248
rect 78388 123208 78430 123248
rect 78470 123208 78512 123248
rect 78552 123208 78561 123248
rect 93295 123208 93304 123248
rect 93344 123208 93386 123248
rect 93426 123208 93468 123248
rect 93508 123208 93550 123248
rect 93590 123208 93632 123248
rect 93672 123208 93681 123248
rect 108415 123208 108424 123248
rect 108464 123208 108506 123248
rect 108546 123208 108588 123248
rect 108628 123208 108670 123248
rect 108710 123208 108752 123248
rect 108792 123208 108801 123248
rect 123535 123208 123544 123248
rect 123584 123208 123626 123248
rect 123666 123208 123708 123248
rect 123748 123208 123790 123248
rect 123830 123208 123872 123248
rect 123912 123208 123921 123248
rect 138655 123208 138664 123248
rect 138704 123208 138746 123248
rect 138786 123208 138828 123248
rect 138868 123208 138910 123248
rect 138950 123208 138992 123248
rect 139032 123208 139041 123248
rect 79415 122452 79424 122492
rect 79464 122452 79506 122492
rect 79546 122452 79588 122492
rect 79628 122452 79670 122492
rect 79710 122452 79752 122492
rect 79792 122452 79801 122492
rect 94535 122452 94544 122492
rect 94584 122452 94626 122492
rect 94666 122452 94708 122492
rect 94748 122452 94790 122492
rect 94830 122452 94872 122492
rect 94912 122452 94921 122492
rect 109655 122452 109664 122492
rect 109704 122452 109746 122492
rect 109786 122452 109828 122492
rect 109868 122452 109910 122492
rect 109950 122452 109992 122492
rect 110032 122452 110041 122492
rect 124775 122452 124784 122492
rect 124824 122452 124866 122492
rect 124906 122452 124948 122492
rect 124988 122452 125030 122492
rect 125070 122452 125112 122492
rect 125152 122452 125161 122492
rect 139895 122452 139904 122492
rect 139944 122452 139986 122492
rect 140026 122452 140068 122492
rect 140108 122452 140150 122492
rect 140190 122452 140232 122492
rect 140272 122452 140281 122492
rect 93763 122408 93821 122409
rect 93678 122368 93772 122408
rect 93812 122368 93821 122408
rect 93763 122367 93821 122368
rect 78175 121696 78184 121736
rect 78224 121696 78266 121736
rect 78306 121696 78348 121736
rect 78388 121696 78430 121736
rect 78470 121696 78512 121736
rect 78552 121696 78561 121736
rect 93295 121696 93304 121736
rect 93344 121696 93386 121736
rect 93426 121696 93468 121736
rect 93508 121696 93550 121736
rect 93590 121696 93632 121736
rect 93672 121696 93681 121736
rect 108415 121696 108424 121736
rect 108464 121696 108506 121736
rect 108546 121696 108588 121736
rect 108628 121696 108670 121736
rect 108710 121696 108752 121736
rect 108792 121696 108801 121736
rect 123535 121696 123544 121736
rect 123584 121696 123626 121736
rect 123666 121696 123708 121736
rect 123748 121696 123790 121736
rect 123830 121696 123872 121736
rect 123912 121696 123921 121736
rect 138655 121696 138664 121736
rect 138704 121696 138746 121736
rect 138786 121696 138828 121736
rect 138868 121696 138910 121736
rect 138950 121696 138992 121736
rect 139032 121696 139041 121736
rect 79415 120940 79424 120980
rect 79464 120940 79506 120980
rect 79546 120940 79588 120980
rect 79628 120940 79670 120980
rect 79710 120940 79752 120980
rect 79792 120940 79801 120980
rect 94535 120940 94544 120980
rect 94584 120940 94626 120980
rect 94666 120940 94708 120980
rect 94748 120940 94790 120980
rect 94830 120940 94872 120980
rect 94912 120940 94921 120980
rect 109655 120940 109664 120980
rect 109704 120940 109746 120980
rect 109786 120940 109828 120980
rect 109868 120940 109910 120980
rect 109950 120940 109992 120980
rect 110032 120940 110041 120980
rect 124775 120940 124784 120980
rect 124824 120940 124866 120980
rect 124906 120940 124948 120980
rect 124988 120940 125030 120980
rect 125070 120940 125112 120980
rect 125152 120940 125161 120980
rect 139895 120940 139904 120980
rect 139944 120940 139986 120980
rect 140026 120940 140068 120980
rect 140108 120940 140150 120980
rect 140190 120940 140232 120980
rect 140272 120940 140281 120980
rect 64099 120856 64108 120896
rect 64148 120856 78892 120896
rect 78932 120856 78941 120896
rect 78175 120184 78184 120224
rect 78224 120184 78266 120224
rect 78306 120184 78348 120224
rect 78388 120184 78430 120224
rect 78470 120184 78512 120224
rect 78552 120184 78561 120224
rect 93295 120184 93304 120224
rect 93344 120184 93386 120224
rect 93426 120184 93468 120224
rect 93508 120184 93550 120224
rect 93590 120184 93632 120224
rect 93672 120184 93681 120224
rect 108415 120184 108424 120224
rect 108464 120184 108506 120224
rect 108546 120184 108588 120224
rect 108628 120184 108670 120224
rect 108710 120184 108752 120224
rect 108792 120184 108801 120224
rect 123535 120184 123544 120224
rect 123584 120184 123626 120224
rect 123666 120184 123708 120224
rect 123748 120184 123790 120224
rect 123830 120184 123872 120224
rect 123912 120184 123921 120224
rect 138655 120184 138664 120224
rect 138704 120184 138746 120224
rect 138786 120184 138828 120224
rect 138868 120184 138910 120224
rect 138950 120184 138992 120224
rect 139032 120184 139041 120224
rect 160012 119636 160052 119700
rect 123139 119596 123148 119636
rect 123188 119596 160052 119636
rect 79415 119428 79424 119468
rect 79464 119428 79506 119468
rect 79546 119428 79588 119468
rect 79628 119428 79670 119468
rect 79710 119428 79752 119468
rect 79792 119428 79801 119468
rect 94535 119428 94544 119468
rect 94584 119428 94626 119468
rect 94666 119428 94708 119468
rect 94748 119428 94790 119468
rect 94830 119428 94872 119468
rect 94912 119428 94921 119468
rect 109655 119428 109664 119468
rect 109704 119428 109746 119468
rect 109786 119428 109828 119468
rect 109868 119428 109910 119468
rect 109950 119428 109992 119468
rect 110032 119428 110041 119468
rect 124775 119428 124784 119468
rect 124824 119428 124866 119468
rect 124906 119428 124948 119468
rect 124988 119428 125030 119468
rect 125070 119428 125112 119468
rect 125152 119428 125161 119468
rect 139895 119428 139904 119468
rect 139944 119428 139986 119468
rect 140026 119428 140068 119468
rect 140108 119428 140150 119468
rect 140190 119428 140232 119468
rect 140272 119428 140281 119468
rect 78175 118672 78184 118712
rect 78224 118672 78266 118712
rect 78306 118672 78348 118712
rect 78388 118672 78430 118712
rect 78470 118672 78512 118712
rect 78552 118672 78561 118712
rect 93295 118672 93304 118712
rect 93344 118672 93386 118712
rect 93426 118672 93468 118712
rect 93508 118672 93550 118712
rect 93590 118672 93632 118712
rect 93672 118672 93681 118712
rect 108415 118672 108424 118712
rect 108464 118672 108506 118712
rect 108546 118672 108588 118712
rect 108628 118672 108670 118712
rect 108710 118672 108752 118712
rect 108792 118672 108801 118712
rect 123535 118672 123544 118712
rect 123584 118672 123626 118712
rect 123666 118672 123708 118712
rect 123748 118672 123790 118712
rect 123830 118672 123872 118712
rect 123912 118672 123921 118712
rect 138655 118672 138664 118712
rect 138704 118672 138746 118712
rect 138786 118672 138828 118712
rect 138868 118672 138910 118712
rect 138950 118672 138992 118712
rect 139032 118672 139041 118712
rect 79415 117916 79424 117956
rect 79464 117916 79506 117956
rect 79546 117916 79588 117956
rect 79628 117916 79670 117956
rect 79710 117916 79752 117956
rect 79792 117916 79801 117956
rect 94535 117916 94544 117956
rect 94584 117916 94626 117956
rect 94666 117916 94708 117956
rect 94748 117916 94790 117956
rect 94830 117916 94872 117956
rect 94912 117916 94921 117956
rect 109655 117916 109664 117956
rect 109704 117916 109746 117956
rect 109786 117916 109828 117956
rect 109868 117916 109910 117956
rect 109950 117916 109992 117956
rect 110032 117916 110041 117956
rect 124775 117916 124784 117956
rect 124824 117916 124866 117956
rect 124906 117916 124948 117956
rect 124988 117916 125030 117956
rect 125070 117916 125112 117956
rect 125152 117916 125161 117956
rect 139895 117916 139904 117956
rect 139944 117916 139986 117956
rect 140026 117916 140068 117956
rect 140108 117916 140150 117956
rect 140190 117916 140232 117956
rect 140272 117916 140281 117956
rect 78175 117160 78184 117200
rect 78224 117160 78266 117200
rect 78306 117160 78348 117200
rect 78388 117160 78430 117200
rect 78470 117160 78512 117200
rect 78552 117160 78561 117200
rect 93295 117160 93304 117200
rect 93344 117160 93386 117200
rect 93426 117160 93468 117200
rect 93508 117160 93550 117200
rect 93590 117160 93632 117200
rect 93672 117160 93681 117200
rect 108415 117160 108424 117200
rect 108464 117160 108506 117200
rect 108546 117160 108588 117200
rect 108628 117160 108670 117200
rect 108710 117160 108752 117200
rect 108792 117160 108801 117200
rect 123535 117160 123544 117200
rect 123584 117160 123626 117200
rect 123666 117160 123708 117200
rect 123748 117160 123790 117200
rect 123830 117160 123872 117200
rect 123912 117160 123921 117200
rect 138655 117160 138664 117200
rect 138704 117160 138746 117200
rect 138786 117160 138828 117200
rect 138868 117160 138910 117200
rect 138950 117160 138992 117200
rect 139032 117160 139041 117200
rect 79415 116404 79424 116444
rect 79464 116404 79506 116444
rect 79546 116404 79588 116444
rect 79628 116404 79670 116444
rect 79710 116404 79752 116444
rect 79792 116404 79801 116444
rect 94535 116404 94544 116444
rect 94584 116404 94626 116444
rect 94666 116404 94708 116444
rect 94748 116404 94790 116444
rect 94830 116404 94872 116444
rect 94912 116404 94921 116444
rect 109655 116404 109664 116444
rect 109704 116404 109746 116444
rect 109786 116404 109828 116444
rect 109868 116404 109910 116444
rect 109950 116404 109992 116444
rect 110032 116404 110041 116444
rect 124775 116404 124784 116444
rect 124824 116404 124866 116444
rect 124906 116404 124948 116444
rect 124988 116404 125030 116444
rect 125070 116404 125112 116444
rect 125152 116404 125161 116444
rect 139895 116404 139904 116444
rect 139944 116404 139986 116444
rect 140026 116404 140068 116444
rect 140108 116404 140150 116444
rect 140190 116404 140232 116444
rect 140272 116404 140281 116444
rect 78175 115648 78184 115688
rect 78224 115648 78266 115688
rect 78306 115648 78348 115688
rect 78388 115648 78430 115688
rect 78470 115648 78512 115688
rect 78552 115648 78561 115688
rect 93295 115648 93304 115688
rect 93344 115648 93386 115688
rect 93426 115648 93468 115688
rect 93508 115648 93550 115688
rect 93590 115648 93632 115688
rect 93672 115648 93681 115688
rect 108415 115648 108424 115688
rect 108464 115648 108506 115688
rect 108546 115648 108588 115688
rect 108628 115648 108670 115688
rect 108710 115648 108752 115688
rect 108792 115648 108801 115688
rect 123535 115648 123544 115688
rect 123584 115648 123626 115688
rect 123666 115648 123708 115688
rect 123748 115648 123790 115688
rect 123830 115648 123872 115688
rect 123912 115648 123921 115688
rect 138655 115648 138664 115688
rect 138704 115648 138746 115688
rect 138786 115648 138828 115688
rect 138868 115648 138910 115688
rect 138950 115648 138992 115688
rect 139032 115648 139041 115688
rect 79415 114892 79424 114932
rect 79464 114892 79506 114932
rect 79546 114892 79588 114932
rect 79628 114892 79670 114932
rect 79710 114892 79752 114932
rect 79792 114892 79801 114932
rect 94535 114892 94544 114932
rect 94584 114892 94626 114932
rect 94666 114892 94708 114932
rect 94748 114892 94790 114932
rect 94830 114892 94872 114932
rect 94912 114892 94921 114932
rect 109655 114892 109664 114932
rect 109704 114892 109746 114932
rect 109786 114892 109828 114932
rect 109868 114892 109910 114932
rect 109950 114892 109992 114932
rect 110032 114892 110041 114932
rect 124775 114892 124784 114932
rect 124824 114892 124866 114932
rect 124906 114892 124948 114932
rect 124988 114892 125030 114932
rect 125070 114892 125112 114932
rect 125152 114892 125161 114932
rect 139895 114892 139904 114932
rect 139944 114892 139986 114932
rect 140026 114892 140068 114932
rect 140108 114892 140150 114932
rect 140190 114892 140232 114932
rect 140272 114892 140281 114932
rect 78175 114136 78184 114176
rect 78224 114136 78266 114176
rect 78306 114136 78348 114176
rect 78388 114136 78430 114176
rect 78470 114136 78512 114176
rect 78552 114136 78561 114176
rect 93295 114136 93304 114176
rect 93344 114136 93386 114176
rect 93426 114136 93468 114176
rect 93508 114136 93550 114176
rect 93590 114136 93632 114176
rect 93672 114136 93681 114176
rect 108415 114136 108424 114176
rect 108464 114136 108506 114176
rect 108546 114136 108588 114176
rect 108628 114136 108670 114176
rect 108710 114136 108752 114176
rect 108792 114136 108801 114176
rect 123535 114136 123544 114176
rect 123584 114136 123626 114176
rect 123666 114136 123708 114176
rect 123748 114136 123790 114176
rect 123830 114136 123872 114176
rect 123912 114136 123921 114176
rect 138655 114136 138664 114176
rect 138704 114136 138746 114176
rect 138786 114136 138828 114176
rect 138868 114136 138910 114176
rect 138950 114136 138992 114176
rect 139032 114136 139041 114176
rect 79415 113380 79424 113420
rect 79464 113380 79506 113420
rect 79546 113380 79588 113420
rect 79628 113380 79670 113420
rect 79710 113380 79752 113420
rect 79792 113380 79801 113420
rect 94535 113380 94544 113420
rect 94584 113380 94626 113420
rect 94666 113380 94708 113420
rect 94748 113380 94790 113420
rect 94830 113380 94872 113420
rect 94912 113380 94921 113420
rect 109655 113380 109664 113420
rect 109704 113380 109746 113420
rect 109786 113380 109828 113420
rect 109868 113380 109910 113420
rect 109950 113380 109992 113420
rect 110032 113380 110041 113420
rect 124775 113380 124784 113420
rect 124824 113380 124866 113420
rect 124906 113380 124948 113420
rect 124988 113380 125030 113420
rect 125070 113380 125112 113420
rect 125152 113380 125161 113420
rect 139895 113380 139904 113420
rect 139944 113380 139986 113420
rect 140026 113380 140068 113420
rect 140108 113380 140150 113420
rect 140190 113380 140232 113420
rect 140272 113380 140281 113420
rect 78175 112624 78184 112664
rect 78224 112624 78266 112664
rect 78306 112624 78348 112664
rect 78388 112624 78430 112664
rect 78470 112624 78512 112664
rect 78552 112624 78561 112664
rect 93295 112624 93304 112664
rect 93344 112624 93386 112664
rect 93426 112624 93468 112664
rect 93508 112624 93550 112664
rect 93590 112624 93632 112664
rect 93672 112624 93681 112664
rect 108415 112624 108424 112664
rect 108464 112624 108506 112664
rect 108546 112624 108588 112664
rect 108628 112624 108670 112664
rect 108710 112624 108752 112664
rect 108792 112624 108801 112664
rect 123535 112624 123544 112664
rect 123584 112624 123626 112664
rect 123666 112624 123708 112664
rect 123748 112624 123790 112664
rect 123830 112624 123872 112664
rect 123912 112624 123921 112664
rect 138655 112624 138664 112664
rect 138704 112624 138746 112664
rect 138786 112624 138828 112664
rect 138868 112624 138910 112664
rect 138950 112624 138992 112664
rect 139032 112624 139041 112664
rect 79415 111868 79424 111908
rect 79464 111868 79506 111908
rect 79546 111868 79588 111908
rect 79628 111868 79670 111908
rect 79710 111868 79752 111908
rect 79792 111868 79801 111908
rect 94535 111868 94544 111908
rect 94584 111868 94626 111908
rect 94666 111868 94708 111908
rect 94748 111868 94790 111908
rect 94830 111868 94872 111908
rect 94912 111868 94921 111908
rect 109655 111868 109664 111908
rect 109704 111868 109746 111908
rect 109786 111868 109828 111908
rect 109868 111868 109910 111908
rect 109950 111868 109992 111908
rect 110032 111868 110041 111908
rect 124775 111868 124784 111908
rect 124824 111868 124866 111908
rect 124906 111868 124948 111908
rect 124988 111868 125030 111908
rect 125070 111868 125112 111908
rect 125152 111868 125161 111908
rect 139895 111868 139904 111908
rect 139944 111868 139986 111908
rect 140026 111868 140068 111908
rect 140108 111868 140150 111908
rect 140190 111868 140232 111908
rect 140272 111868 140281 111908
rect 78175 111112 78184 111152
rect 78224 111112 78266 111152
rect 78306 111112 78348 111152
rect 78388 111112 78430 111152
rect 78470 111112 78512 111152
rect 78552 111112 78561 111152
rect 93295 111112 93304 111152
rect 93344 111112 93386 111152
rect 93426 111112 93468 111152
rect 93508 111112 93550 111152
rect 93590 111112 93632 111152
rect 93672 111112 93681 111152
rect 108415 111112 108424 111152
rect 108464 111112 108506 111152
rect 108546 111112 108588 111152
rect 108628 111112 108670 111152
rect 108710 111112 108752 111152
rect 108792 111112 108801 111152
rect 123535 111112 123544 111152
rect 123584 111112 123626 111152
rect 123666 111112 123708 111152
rect 123748 111112 123790 111152
rect 123830 111112 123872 111152
rect 123912 111112 123921 111152
rect 138655 111112 138664 111152
rect 138704 111112 138746 111152
rect 138786 111112 138828 111152
rect 138868 111112 138910 111152
rect 138950 111112 138992 111152
rect 139032 111112 139041 111152
rect 79415 110356 79424 110396
rect 79464 110356 79506 110396
rect 79546 110356 79588 110396
rect 79628 110356 79670 110396
rect 79710 110356 79752 110396
rect 79792 110356 79801 110396
rect 94535 110356 94544 110396
rect 94584 110356 94626 110396
rect 94666 110356 94708 110396
rect 94748 110356 94790 110396
rect 94830 110356 94872 110396
rect 94912 110356 94921 110396
rect 109655 110356 109664 110396
rect 109704 110356 109746 110396
rect 109786 110356 109828 110396
rect 109868 110356 109910 110396
rect 109950 110356 109992 110396
rect 110032 110356 110041 110396
rect 124775 110356 124784 110396
rect 124824 110356 124866 110396
rect 124906 110356 124948 110396
rect 124988 110356 125030 110396
rect 125070 110356 125112 110396
rect 125152 110356 125161 110396
rect 139895 110356 139904 110396
rect 139944 110356 139986 110396
rect 140026 110356 140068 110396
rect 140108 110356 140150 110396
rect 140190 110356 140232 110396
rect 140272 110356 140281 110396
rect 78175 109600 78184 109640
rect 78224 109600 78266 109640
rect 78306 109600 78348 109640
rect 78388 109600 78430 109640
rect 78470 109600 78512 109640
rect 78552 109600 78561 109640
rect 93295 109600 93304 109640
rect 93344 109600 93386 109640
rect 93426 109600 93468 109640
rect 93508 109600 93550 109640
rect 93590 109600 93632 109640
rect 93672 109600 93681 109640
rect 108415 109600 108424 109640
rect 108464 109600 108506 109640
rect 108546 109600 108588 109640
rect 108628 109600 108670 109640
rect 108710 109600 108752 109640
rect 108792 109600 108801 109640
rect 123535 109600 123544 109640
rect 123584 109600 123626 109640
rect 123666 109600 123708 109640
rect 123748 109600 123790 109640
rect 123830 109600 123872 109640
rect 123912 109600 123921 109640
rect 138655 109600 138664 109640
rect 138704 109600 138746 109640
rect 138786 109600 138828 109640
rect 138868 109600 138910 109640
rect 138950 109600 138992 109640
rect 139032 109600 139041 109640
rect 79415 108844 79424 108884
rect 79464 108844 79506 108884
rect 79546 108844 79588 108884
rect 79628 108844 79670 108884
rect 79710 108844 79752 108884
rect 79792 108844 79801 108884
rect 94535 108844 94544 108884
rect 94584 108844 94626 108884
rect 94666 108844 94708 108884
rect 94748 108844 94790 108884
rect 94830 108844 94872 108884
rect 94912 108844 94921 108884
rect 109655 108844 109664 108884
rect 109704 108844 109746 108884
rect 109786 108844 109828 108884
rect 109868 108844 109910 108884
rect 109950 108844 109992 108884
rect 110032 108844 110041 108884
rect 124775 108844 124784 108884
rect 124824 108844 124866 108884
rect 124906 108844 124948 108884
rect 124988 108844 125030 108884
rect 125070 108844 125112 108884
rect 125152 108844 125161 108884
rect 139895 108844 139904 108884
rect 139944 108844 139986 108884
rect 140026 108844 140068 108884
rect 140108 108844 140150 108884
rect 140190 108844 140232 108884
rect 140272 108844 140281 108884
rect 78175 108088 78184 108128
rect 78224 108088 78266 108128
rect 78306 108088 78348 108128
rect 78388 108088 78430 108128
rect 78470 108088 78512 108128
rect 78552 108088 78561 108128
rect 93295 108088 93304 108128
rect 93344 108088 93386 108128
rect 93426 108088 93468 108128
rect 93508 108088 93550 108128
rect 93590 108088 93632 108128
rect 93672 108088 93681 108128
rect 108415 108088 108424 108128
rect 108464 108088 108506 108128
rect 108546 108088 108588 108128
rect 108628 108088 108670 108128
rect 108710 108088 108752 108128
rect 108792 108088 108801 108128
rect 123535 108088 123544 108128
rect 123584 108088 123626 108128
rect 123666 108088 123708 108128
rect 123748 108088 123790 108128
rect 123830 108088 123872 108128
rect 123912 108088 123921 108128
rect 138655 108088 138664 108128
rect 138704 108088 138746 108128
rect 138786 108088 138828 108128
rect 138868 108088 138910 108128
rect 138950 108088 138992 108128
rect 139032 108088 139041 108128
rect 79415 107332 79424 107372
rect 79464 107332 79506 107372
rect 79546 107332 79588 107372
rect 79628 107332 79670 107372
rect 79710 107332 79752 107372
rect 79792 107332 79801 107372
rect 94535 107332 94544 107372
rect 94584 107332 94626 107372
rect 94666 107332 94708 107372
rect 94748 107332 94790 107372
rect 94830 107332 94872 107372
rect 94912 107332 94921 107372
rect 109655 107332 109664 107372
rect 109704 107332 109746 107372
rect 109786 107332 109828 107372
rect 109868 107332 109910 107372
rect 109950 107332 109992 107372
rect 110032 107332 110041 107372
rect 124775 107332 124784 107372
rect 124824 107332 124866 107372
rect 124906 107332 124948 107372
rect 124988 107332 125030 107372
rect 125070 107332 125112 107372
rect 125152 107332 125161 107372
rect 139895 107332 139904 107372
rect 139944 107332 139986 107372
rect 140026 107332 140068 107372
rect 140108 107332 140150 107372
rect 140190 107332 140232 107372
rect 140272 107332 140281 107372
rect 78175 106576 78184 106616
rect 78224 106576 78266 106616
rect 78306 106576 78348 106616
rect 78388 106576 78430 106616
rect 78470 106576 78512 106616
rect 78552 106576 78561 106616
rect 93295 106576 93304 106616
rect 93344 106576 93386 106616
rect 93426 106576 93468 106616
rect 93508 106576 93550 106616
rect 93590 106576 93632 106616
rect 93672 106576 93681 106616
rect 108415 106576 108424 106616
rect 108464 106576 108506 106616
rect 108546 106576 108588 106616
rect 108628 106576 108670 106616
rect 108710 106576 108752 106616
rect 108792 106576 108801 106616
rect 123535 106576 123544 106616
rect 123584 106576 123626 106616
rect 123666 106576 123708 106616
rect 123748 106576 123790 106616
rect 123830 106576 123872 106616
rect 123912 106576 123921 106616
rect 138655 106576 138664 106616
rect 138704 106576 138746 106616
rect 138786 106576 138828 106616
rect 138868 106576 138910 106616
rect 138950 106576 138992 106616
rect 139032 106576 139041 106616
rect 79415 105820 79424 105860
rect 79464 105820 79506 105860
rect 79546 105820 79588 105860
rect 79628 105820 79670 105860
rect 79710 105820 79752 105860
rect 79792 105820 79801 105860
rect 94535 105820 94544 105860
rect 94584 105820 94626 105860
rect 94666 105820 94708 105860
rect 94748 105820 94790 105860
rect 94830 105820 94872 105860
rect 94912 105820 94921 105860
rect 109655 105820 109664 105860
rect 109704 105820 109746 105860
rect 109786 105820 109828 105860
rect 109868 105820 109910 105860
rect 109950 105820 109992 105860
rect 110032 105820 110041 105860
rect 124775 105820 124784 105860
rect 124824 105820 124866 105860
rect 124906 105820 124948 105860
rect 124988 105820 125030 105860
rect 125070 105820 125112 105860
rect 125152 105820 125161 105860
rect 139895 105820 139904 105860
rect 139944 105820 139986 105860
rect 140026 105820 140068 105860
rect 140108 105820 140150 105860
rect 140190 105820 140232 105860
rect 140272 105820 140281 105860
rect 78175 105064 78184 105104
rect 78224 105064 78266 105104
rect 78306 105064 78348 105104
rect 78388 105064 78430 105104
rect 78470 105064 78512 105104
rect 78552 105064 78561 105104
rect 93295 105064 93304 105104
rect 93344 105064 93386 105104
rect 93426 105064 93468 105104
rect 93508 105064 93550 105104
rect 93590 105064 93632 105104
rect 93672 105064 93681 105104
rect 108415 105064 108424 105104
rect 108464 105064 108506 105104
rect 108546 105064 108588 105104
rect 108628 105064 108670 105104
rect 108710 105064 108752 105104
rect 108792 105064 108801 105104
rect 123535 105064 123544 105104
rect 123584 105064 123626 105104
rect 123666 105064 123708 105104
rect 123748 105064 123790 105104
rect 123830 105064 123872 105104
rect 123912 105064 123921 105104
rect 138655 105064 138664 105104
rect 138704 105064 138746 105104
rect 138786 105064 138828 105104
rect 138868 105064 138910 105104
rect 138950 105064 138992 105104
rect 139032 105064 139041 105104
rect 64099 104980 64108 105020
rect 64148 104980 94444 105020
rect 94484 104980 94493 105020
rect 79415 104308 79424 104348
rect 79464 104308 79506 104348
rect 79546 104308 79588 104348
rect 79628 104308 79670 104348
rect 79710 104308 79752 104348
rect 79792 104308 79801 104348
rect 94535 104308 94544 104348
rect 94584 104308 94626 104348
rect 94666 104308 94708 104348
rect 94748 104308 94790 104348
rect 94830 104308 94872 104348
rect 94912 104308 94921 104348
rect 109655 104308 109664 104348
rect 109704 104308 109746 104348
rect 109786 104308 109828 104348
rect 109868 104308 109910 104348
rect 109950 104308 109992 104348
rect 110032 104308 110041 104348
rect 124775 104308 124784 104348
rect 124824 104308 124866 104348
rect 124906 104308 124948 104348
rect 124988 104308 125030 104348
rect 125070 104308 125112 104348
rect 125152 104308 125161 104348
rect 139895 104308 139904 104348
rect 139944 104308 139986 104348
rect 140026 104308 140068 104348
rect 140108 104308 140150 104348
rect 140190 104308 140232 104348
rect 140272 104308 140281 104348
rect 121603 103720 121612 103760
rect 121652 103720 160032 103760
rect 78175 103552 78184 103592
rect 78224 103552 78266 103592
rect 78306 103552 78348 103592
rect 78388 103552 78430 103592
rect 78470 103552 78512 103592
rect 78552 103552 78561 103592
rect 93295 103552 93304 103592
rect 93344 103552 93386 103592
rect 93426 103552 93468 103592
rect 93508 103552 93550 103592
rect 93590 103552 93632 103592
rect 93672 103552 93681 103592
rect 108415 103552 108424 103592
rect 108464 103552 108506 103592
rect 108546 103552 108588 103592
rect 108628 103552 108670 103592
rect 108710 103552 108752 103592
rect 108792 103552 108801 103592
rect 123535 103552 123544 103592
rect 123584 103552 123626 103592
rect 123666 103552 123708 103592
rect 123748 103552 123790 103592
rect 123830 103552 123872 103592
rect 123912 103552 123921 103592
rect 138655 103552 138664 103592
rect 138704 103552 138746 103592
rect 138786 103552 138828 103592
rect 138868 103552 138910 103592
rect 138950 103552 138992 103592
rect 139032 103552 139041 103592
rect 79415 102796 79424 102836
rect 79464 102796 79506 102836
rect 79546 102796 79588 102836
rect 79628 102796 79670 102836
rect 79710 102796 79752 102836
rect 79792 102796 79801 102836
rect 94535 102796 94544 102836
rect 94584 102796 94626 102836
rect 94666 102796 94708 102836
rect 94748 102796 94790 102836
rect 94830 102796 94872 102836
rect 94912 102796 94921 102836
rect 109655 102796 109664 102836
rect 109704 102796 109746 102836
rect 109786 102796 109828 102836
rect 109868 102796 109910 102836
rect 109950 102796 109992 102836
rect 110032 102796 110041 102836
rect 124775 102796 124784 102836
rect 124824 102796 124866 102836
rect 124906 102796 124948 102836
rect 124988 102796 125030 102836
rect 125070 102796 125112 102836
rect 125152 102796 125161 102836
rect 139895 102796 139904 102836
rect 139944 102796 139986 102836
rect 140026 102796 140068 102836
rect 140108 102796 140150 102836
rect 140190 102796 140232 102836
rect 140272 102796 140281 102836
rect 78175 102040 78184 102080
rect 78224 102040 78266 102080
rect 78306 102040 78348 102080
rect 78388 102040 78430 102080
rect 78470 102040 78512 102080
rect 78552 102040 78561 102080
rect 93295 102040 93304 102080
rect 93344 102040 93386 102080
rect 93426 102040 93468 102080
rect 93508 102040 93550 102080
rect 93590 102040 93632 102080
rect 93672 102040 93681 102080
rect 108415 102040 108424 102080
rect 108464 102040 108506 102080
rect 108546 102040 108588 102080
rect 108628 102040 108670 102080
rect 108710 102040 108752 102080
rect 108792 102040 108801 102080
rect 123535 102040 123544 102080
rect 123584 102040 123626 102080
rect 123666 102040 123708 102080
rect 123748 102040 123790 102080
rect 123830 102040 123872 102080
rect 123912 102040 123921 102080
rect 138655 102040 138664 102080
rect 138704 102040 138746 102080
rect 138786 102040 138828 102080
rect 138868 102040 138910 102080
rect 138950 102040 138992 102080
rect 139032 102040 139041 102080
rect 79415 101284 79424 101324
rect 79464 101284 79506 101324
rect 79546 101284 79588 101324
rect 79628 101284 79670 101324
rect 79710 101284 79752 101324
rect 79792 101284 79801 101324
rect 94535 101284 94544 101324
rect 94584 101284 94626 101324
rect 94666 101284 94708 101324
rect 94748 101284 94790 101324
rect 94830 101284 94872 101324
rect 94912 101284 94921 101324
rect 109655 101284 109664 101324
rect 109704 101284 109746 101324
rect 109786 101284 109828 101324
rect 109868 101284 109910 101324
rect 109950 101284 109992 101324
rect 110032 101284 110041 101324
rect 124775 101284 124784 101324
rect 124824 101284 124866 101324
rect 124906 101284 124948 101324
rect 124988 101284 125030 101324
rect 125070 101284 125112 101324
rect 125152 101284 125161 101324
rect 139895 101284 139904 101324
rect 139944 101284 139986 101324
rect 140026 101284 140068 101324
rect 140108 101284 140150 101324
rect 140190 101284 140232 101324
rect 140272 101284 140281 101324
rect 78175 100528 78184 100568
rect 78224 100528 78266 100568
rect 78306 100528 78348 100568
rect 78388 100528 78430 100568
rect 78470 100528 78512 100568
rect 78552 100528 78561 100568
rect 93295 100528 93304 100568
rect 93344 100528 93386 100568
rect 93426 100528 93468 100568
rect 93508 100528 93550 100568
rect 93590 100528 93632 100568
rect 93672 100528 93681 100568
rect 108415 100528 108424 100568
rect 108464 100528 108506 100568
rect 108546 100528 108588 100568
rect 108628 100528 108670 100568
rect 108710 100528 108752 100568
rect 108792 100528 108801 100568
rect 123535 100528 123544 100568
rect 123584 100528 123626 100568
rect 123666 100528 123708 100568
rect 123748 100528 123790 100568
rect 123830 100528 123872 100568
rect 123912 100528 123921 100568
rect 138655 100528 138664 100568
rect 138704 100528 138746 100568
rect 138786 100528 138828 100568
rect 138868 100528 138910 100568
rect 138950 100528 138992 100568
rect 139032 100528 139041 100568
rect 79415 99772 79424 99812
rect 79464 99772 79506 99812
rect 79546 99772 79588 99812
rect 79628 99772 79670 99812
rect 79710 99772 79752 99812
rect 79792 99772 79801 99812
rect 94535 99772 94544 99812
rect 94584 99772 94626 99812
rect 94666 99772 94708 99812
rect 94748 99772 94790 99812
rect 94830 99772 94872 99812
rect 94912 99772 94921 99812
rect 109655 99772 109664 99812
rect 109704 99772 109746 99812
rect 109786 99772 109828 99812
rect 109868 99772 109910 99812
rect 109950 99772 109992 99812
rect 110032 99772 110041 99812
rect 124775 99772 124784 99812
rect 124824 99772 124866 99812
rect 124906 99772 124948 99812
rect 124988 99772 125030 99812
rect 125070 99772 125112 99812
rect 125152 99772 125161 99812
rect 139895 99772 139904 99812
rect 139944 99772 139986 99812
rect 140026 99772 140068 99812
rect 140108 99772 140150 99812
rect 140190 99772 140232 99812
rect 140272 99772 140281 99812
rect 78175 99016 78184 99056
rect 78224 99016 78266 99056
rect 78306 99016 78348 99056
rect 78388 99016 78430 99056
rect 78470 99016 78512 99056
rect 78552 99016 78561 99056
rect 93295 99016 93304 99056
rect 93344 99016 93386 99056
rect 93426 99016 93468 99056
rect 93508 99016 93550 99056
rect 93590 99016 93632 99056
rect 93672 99016 93681 99056
rect 108415 99016 108424 99056
rect 108464 99016 108506 99056
rect 108546 99016 108588 99056
rect 108628 99016 108670 99056
rect 108710 99016 108752 99056
rect 108792 99016 108801 99056
rect 123535 99016 123544 99056
rect 123584 99016 123626 99056
rect 123666 99016 123708 99056
rect 123748 99016 123790 99056
rect 123830 99016 123872 99056
rect 123912 99016 123921 99056
rect 138655 99016 138664 99056
rect 138704 99016 138746 99056
rect 138786 99016 138828 99056
rect 138868 99016 138910 99056
rect 138950 99016 138992 99056
rect 139032 99016 139041 99056
rect 79415 98260 79424 98300
rect 79464 98260 79506 98300
rect 79546 98260 79588 98300
rect 79628 98260 79670 98300
rect 79710 98260 79752 98300
rect 79792 98260 79801 98300
rect 94535 98260 94544 98300
rect 94584 98260 94626 98300
rect 94666 98260 94708 98300
rect 94748 98260 94790 98300
rect 94830 98260 94872 98300
rect 94912 98260 94921 98300
rect 109655 98260 109664 98300
rect 109704 98260 109746 98300
rect 109786 98260 109828 98300
rect 109868 98260 109910 98300
rect 109950 98260 109992 98300
rect 110032 98260 110041 98300
rect 124775 98260 124784 98300
rect 124824 98260 124866 98300
rect 124906 98260 124948 98300
rect 124988 98260 125030 98300
rect 125070 98260 125112 98300
rect 125152 98260 125161 98300
rect 139895 98260 139904 98300
rect 139944 98260 139986 98300
rect 140026 98260 140068 98300
rect 140108 98260 140150 98300
rect 140190 98260 140232 98300
rect 140272 98260 140281 98300
rect 78175 97504 78184 97544
rect 78224 97504 78266 97544
rect 78306 97504 78348 97544
rect 78388 97504 78430 97544
rect 78470 97504 78512 97544
rect 78552 97504 78561 97544
rect 93295 97504 93304 97544
rect 93344 97504 93386 97544
rect 93426 97504 93468 97544
rect 93508 97504 93550 97544
rect 93590 97504 93632 97544
rect 93672 97504 93681 97544
rect 108415 97504 108424 97544
rect 108464 97504 108506 97544
rect 108546 97504 108588 97544
rect 108628 97504 108670 97544
rect 108710 97504 108752 97544
rect 108792 97504 108801 97544
rect 123535 97504 123544 97544
rect 123584 97504 123626 97544
rect 123666 97504 123708 97544
rect 123748 97504 123790 97544
rect 123830 97504 123872 97544
rect 123912 97504 123921 97544
rect 138655 97504 138664 97544
rect 138704 97504 138746 97544
rect 138786 97504 138828 97544
rect 138868 97504 138910 97544
rect 138950 97504 138992 97544
rect 139032 97504 139041 97544
rect 79415 96748 79424 96788
rect 79464 96748 79506 96788
rect 79546 96748 79588 96788
rect 79628 96748 79670 96788
rect 79710 96748 79752 96788
rect 79792 96748 79801 96788
rect 94535 96748 94544 96788
rect 94584 96748 94626 96788
rect 94666 96748 94708 96788
rect 94748 96748 94790 96788
rect 94830 96748 94872 96788
rect 94912 96748 94921 96788
rect 109655 96748 109664 96788
rect 109704 96748 109746 96788
rect 109786 96748 109828 96788
rect 109868 96748 109910 96788
rect 109950 96748 109992 96788
rect 110032 96748 110041 96788
rect 124775 96748 124784 96788
rect 124824 96748 124866 96788
rect 124906 96748 124948 96788
rect 124988 96748 125030 96788
rect 125070 96748 125112 96788
rect 125152 96748 125161 96788
rect 139895 96748 139904 96788
rect 139944 96748 139986 96788
rect 140026 96748 140068 96788
rect 140108 96748 140150 96788
rect 140190 96748 140232 96788
rect 140272 96748 140281 96788
rect 78175 95992 78184 96032
rect 78224 95992 78266 96032
rect 78306 95992 78348 96032
rect 78388 95992 78430 96032
rect 78470 95992 78512 96032
rect 78552 95992 78561 96032
rect 93295 95992 93304 96032
rect 93344 95992 93386 96032
rect 93426 95992 93468 96032
rect 93508 95992 93550 96032
rect 93590 95992 93632 96032
rect 93672 95992 93681 96032
rect 108415 95992 108424 96032
rect 108464 95992 108506 96032
rect 108546 95992 108588 96032
rect 108628 95992 108670 96032
rect 108710 95992 108752 96032
rect 108792 95992 108801 96032
rect 123535 95992 123544 96032
rect 123584 95992 123626 96032
rect 123666 95992 123708 96032
rect 123748 95992 123790 96032
rect 123830 95992 123872 96032
rect 123912 95992 123921 96032
rect 138655 95992 138664 96032
rect 138704 95992 138746 96032
rect 138786 95992 138828 96032
rect 138868 95992 138910 96032
rect 138950 95992 138992 96032
rect 139032 95992 139041 96032
rect 88003 95572 88012 95612
rect 88052 95572 103660 95612
rect 103700 95572 103709 95612
rect 79415 95236 79424 95276
rect 79464 95236 79506 95276
rect 79546 95236 79588 95276
rect 79628 95236 79670 95276
rect 79710 95236 79752 95276
rect 79792 95236 79801 95276
rect 94535 95236 94544 95276
rect 94584 95236 94626 95276
rect 94666 95236 94708 95276
rect 94748 95236 94790 95276
rect 94830 95236 94872 95276
rect 94912 95236 94921 95276
rect 109655 95236 109664 95276
rect 109704 95236 109746 95276
rect 109786 95236 109828 95276
rect 109868 95236 109910 95276
rect 109950 95236 109992 95276
rect 110032 95236 110041 95276
rect 124775 95236 124784 95276
rect 124824 95236 124866 95276
rect 124906 95236 124948 95276
rect 124988 95236 125030 95276
rect 125070 95236 125112 95276
rect 125152 95236 125161 95276
rect 139895 95236 139904 95276
rect 139944 95236 139986 95276
rect 140026 95236 140068 95276
rect 140108 95236 140150 95276
rect 140190 95236 140232 95276
rect 140272 95236 140281 95276
rect 78175 94480 78184 94520
rect 78224 94480 78266 94520
rect 78306 94480 78348 94520
rect 78388 94480 78430 94520
rect 78470 94480 78512 94520
rect 78552 94480 78561 94520
rect 93295 94480 93304 94520
rect 93344 94480 93386 94520
rect 93426 94480 93468 94520
rect 93508 94480 93550 94520
rect 93590 94480 93632 94520
rect 93672 94480 93681 94520
rect 108415 94480 108424 94520
rect 108464 94480 108506 94520
rect 108546 94480 108588 94520
rect 108628 94480 108670 94520
rect 108710 94480 108752 94520
rect 108792 94480 108801 94520
rect 123535 94480 123544 94520
rect 123584 94480 123626 94520
rect 123666 94480 123708 94520
rect 123748 94480 123790 94520
rect 123830 94480 123872 94520
rect 123912 94480 123921 94520
rect 138655 94480 138664 94520
rect 138704 94480 138746 94520
rect 138786 94480 138828 94520
rect 138868 94480 138910 94520
rect 138950 94480 138992 94520
rect 139032 94480 139041 94520
rect 79415 93724 79424 93764
rect 79464 93724 79506 93764
rect 79546 93724 79588 93764
rect 79628 93724 79670 93764
rect 79710 93724 79752 93764
rect 79792 93724 79801 93764
rect 94535 93724 94544 93764
rect 94584 93724 94626 93764
rect 94666 93724 94708 93764
rect 94748 93724 94790 93764
rect 94830 93724 94872 93764
rect 94912 93724 94921 93764
rect 109655 93724 109664 93764
rect 109704 93724 109746 93764
rect 109786 93724 109828 93764
rect 109868 93724 109910 93764
rect 109950 93724 109992 93764
rect 110032 93724 110041 93764
rect 124775 93724 124784 93764
rect 124824 93724 124866 93764
rect 124906 93724 124948 93764
rect 124988 93724 125030 93764
rect 125070 93724 125112 93764
rect 125152 93724 125161 93764
rect 139895 93724 139904 93764
rect 139944 93724 139986 93764
rect 140026 93724 140068 93764
rect 140108 93724 140150 93764
rect 140190 93724 140232 93764
rect 140272 93724 140281 93764
rect 78175 92968 78184 93008
rect 78224 92968 78266 93008
rect 78306 92968 78348 93008
rect 78388 92968 78430 93008
rect 78470 92968 78512 93008
rect 78552 92968 78561 93008
rect 93295 92968 93304 93008
rect 93344 92968 93386 93008
rect 93426 92968 93468 93008
rect 93508 92968 93550 93008
rect 93590 92968 93632 93008
rect 93672 92968 93681 93008
rect 108415 92968 108424 93008
rect 108464 92968 108506 93008
rect 108546 92968 108588 93008
rect 108628 92968 108670 93008
rect 108710 92968 108752 93008
rect 108792 92968 108801 93008
rect 123535 92968 123544 93008
rect 123584 92968 123626 93008
rect 123666 92968 123708 93008
rect 123748 92968 123790 93008
rect 123830 92968 123872 93008
rect 123912 92968 123921 93008
rect 138655 92968 138664 93008
rect 138704 92968 138746 93008
rect 138786 92968 138828 93008
rect 138868 92968 138910 93008
rect 138950 92968 138992 93008
rect 139032 92968 139041 93008
rect 79415 92212 79424 92252
rect 79464 92212 79506 92252
rect 79546 92212 79588 92252
rect 79628 92212 79670 92252
rect 79710 92212 79752 92252
rect 79792 92212 79801 92252
rect 94535 92212 94544 92252
rect 94584 92212 94626 92252
rect 94666 92212 94708 92252
rect 94748 92212 94790 92252
rect 94830 92212 94872 92252
rect 94912 92212 94921 92252
rect 109655 92212 109664 92252
rect 109704 92212 109746 92252
rect 109786 92212 109828 92252
rect 109868 92212 109910 92252
rect 109950 92212 109992 92252
rect 110032 92212 110041 92252
rect 124775 92212 124784 92252
rect 124824 92212 124866 92252
rect 124906 92212 124948 92252
rect 124988 92212 125030 92252
rect 125070 92212 125112 92252
rect 125152 92212 125161 92252
rect 139895 92212 139904 92252
rect 139944 92212 139986 92252
rect 140026 92212 140068 92252
rect 140108 92212 140150 92252
rect 140190 92212 140232 92252
rect 140272 92212 140281 92252
rect 78175 91456 78184 91496
rect 78224 91456 78266 91496
rect 78306 91456 78348 91496
rect 78388 91456 78430 91496
rect 78470 91456 78512 91496
rect 78552 91456 78561 91496
rect 93295 91456 93304 91496
rect 93344 91456 93386 91496
rect 93426 91456 93468 91496
rect 93508 91456 93550 91496
rect 93590 91456 93632 91496
rect 93672 91456 93681 91496
rect 108415 91456 108424 91496
rect 108464 91456 108506 91496
rect 108546 91456 108588 91496
rect 108628 91456 108670 91496
rect 108710 91456 108752 91496
rect 108792 91456 108801 91496
rect 123535 91456 123544 91496
rect 123584 91456 123626 91496
rect 123666 91456 123708 91496
rect 123748 91456 123790 91496
rect 123830 91456 123872 91496
rect 123912 91456 123921 91496
rect 138655 91456 138664 91496
rect 138704 91456 138746 91496
rect 138786 91456 138828 91496
rect 138868 91456 138910 91496
rect 138950 91456 138992 91496
rect 139032 91456 139041 91496
rect 79415 90700 79424 90740
rect 79464 90700 79506 90740
rect 79546 90700 79588 90740
rect 79628 90700 79670 90740
rect 79710 90700 79752 90740
rect 79792 90700 79801 90740
rect 94535 90700 94544 90740
rect 94584 90700 94626 90740
rect 94666 90700 94708 90740
rect 94748 90700 94790 90740
rect 94830 90700 94872 90740
rect 94912 90700 94921 90740
rect 109655 90700 109664 90740
rect 109704 90700 109746 90740
rect 109786 90700 109828 90740
rect 109868 90700 109910 90740
rect 109950 90700 109992 90740
rect 110032 90700 110041 90740
rect 124775 90700 124784 90740
rect 124824 90700 124866 90740
rect 124906 90700 124948 90740
rect 124988 90700 125030 90740
rect 125070 90700 125112 90740
rect 125152 90700 125161 90740
rect 139895 90700 139904 90740
rect 139944 90700 139986 90740
rect 140026 90700 140068 90740
rect 140108 90700 140150 90740
rect 140190 90700 140232 90740
rect 140272 90700 140281 90740
rect 78175 89944 78184 89984
rect 78224 89944 78266 89984
rect 78306 89944 78348 89984
rect 78388 89944 78430 89984
rect 78470 89944 78512 89984
rect 78552 89944 78561 89984
rect 93295 89944 93304 89984
rect 93344 89944 93386 89984
rect 93426 89944 93468 89984
rect 93508 89944 93550 89984
rect 93590 89944 93632 89984
rect 93672 89944 93681 89984
rect 108415 89944 108424 89984
rect 108464 89944 108506 89984
rect 108546 89944 108588 89984
rect 108628 89944 108670 89984
rect 108710 89944 108752 89984
rect 108792 89944 108801 89984
rect 123535 89944 123544 89984
rect 123584 89944 123626 89984
rect 123666 89944 123708 89984
rect 123748 89944 123790 89984
rect 123830 89944 123872 89984
rect 123912 89944 123921 89984
rect 138655 89944 138664 89984
rect 138704 89944 138746 89984
rect 138786 89944 138828 89984
rect 138868 89944 138910 89984
rect 138950 89944 138992 89984
rect 139032 89944 139041 89984
rect 79415 89188 79424 89228
rect 79464 89188 79506 89228
rect 79546 89188 79588 89228
rect 79628 89188 79670 89228
rect 79710 89188 79752 89228
rect 79792 89188 79801 89228
rect 94535 89188 94544 89228
rect 94584 89188 94626 89228
rect 94666 89188 94708 89228
rect 94748 89188 94790 89228
rect 94830 89188 94872 89228
rect 94912 89188 94921 89228
rect 109655 89188 109664 89228
rect 109704 89188 109746 89228
rect 109786 89188 109828 89228
rect 109868 89188 109910 89228
rect 109950 89188 109992 89228
rect 110032 89188 110041 89228
rect 124775 89188 124784 89228
rect 124824 89188 124866 89228
rect 124906 89188 124948 89228
rect 124988 89188 125030 89228
rect 125070 89188 125112 89228
rect 125152 89188 125161 89228
rect 139895 89188 139904 89228
rect 139944 89188 139986 89228
rect 140026 89188 140068 89228
rect 140108 89188 140150 89228
rect 140190 89188 140232 89228
rect 140272 89188 140281 89228
rect 90691 89144 90749 89145
rect 64108 89104 90700 89144
rect 90740 89104 90749 89144
rect 64108 88010 64148 89104
rect 90691 89103 90749 89104
rect 92131 89144 92189 89145
rect 92131 89104 92140 89144
rect 92180 89104 94252 89144
rect 94292 89104 94301 89144
rect 92131 89103 92189 89104
rect 78175 88432 78184 88472
rect 78224 88432 78266 88472
rect 78306 88432 78348 88472
rect 78388 88432 78430 88472
rect 78470 88432 78512 88472
rect 78552 88432 78561 88472
rect 93295 88432 93304 88472
rect 93344 88432 93386 88472
rect 93426 88432 93468 88472
rect 93508 88432 93550 88472
rect 93590 88432 93632 88472
rect 93672 88432 93681 88472
rect 108415 88432 108424 88472
rect 108464 88432 108506 88472
rect 108546 88432 108588 88472
rect 108628 88432 108670 88472
rect 108710 88432 108752 88472
rect 108792 88432 108801 88472
rect 123535 88432 123544 88472
rect 123584 88432 123626 88472
rect 123666 88432 123708 88472
rect 123748 88432 123790 88472
rect 123830 88432 123872 88472
rect 123912 88432 123921 88472
rect 138655 88432 138664 88472
rect 138704 88432 138746 88472
rect 138786 88432 138828 88472
rect 138868 88432 138910 88472
rect 138950 88432 138992 88472
rect 139032 88432 139041 88472
rect 64099 87970 64108 88010
rect 64148 87970 64157 88010
rect 148195 87844 148204 87884
rect 148244 87844 160032 87884
rect 79415 87676 79424 87716
rect 79464 87676 79506 87716
rect 79546 87676 79588 87716
rect 79628 87676 79670 87716
rect 79710 87676 79752 87716
rect 79792 87676 79801 87716
rect 94535 87676 94544 87716
rect 94584 87676 94626 87716
rect 94666 87676 94708 87716
rect 94748 87676 94790 87716
rect 94830 87676 94872 87716
rect 94912 87676 94921 87716
rect 109655 87676 109664 87716
rect 109704 87676 109746 87716
rect 109786 87676 109828 87716
rect 109868 87676 109910 87716
rect 109950 87676 109992 87716
rect 110032 87676 110041 87716
rect 124775 87676 124784 87716
rect 124824 87676 124866 87716
rect 124906 87676 124948 87716
rect 124988 87676 125030 87716
rect 125070 87676 125112 87716
rect 125152 87676 125161 87716
rect 139895 87676 139904 87716
rect 139944 87676 139986 87716
rect 140026 87676 140068 87716
rect 140108 87676 140150 87716
rect 140190 87676 140232 87716
rect 140272 87676 140281 87716
rect 78175 86920 78184 86960
rect 78224 86920 78266 86960
rect 78306 86920 78348 86960
rect 78388 86920 78430 86960
rect 78470 86920 78512 86960
rect 78552 86920 78561 86960
rect 93295 86920 93304 86960
rect 93344 86920 93386 86960
rect 93426 86920 93468 86960
rect 93508 86920 93550 86960
rect 93590 86920 93632 86960
rect 93672 86920 93681 86960
rect 108415 86920 108424 86960
rect 108464 86920 108506 86960
rect 108546 86920 108588 86960
rect 108628 86920 108670 86960
rect 108710 86920 108752 86960
rect 108792 86920 108801 86960
rect 123535 86920 123544 86960
rect 123584 86920 123626 86960
rect 123666 86920 123708 86960
rect 123748 86920 123790 86960
rect 123830 86920 123872 86960
rect 123912 86920 123921 86960
rect 138655 86920 138664 86960
rect 138704 86920 138746 86960
rect 138786 86920 138828 86960
rect 138868 86920 138910 86960
rect 138950 86920 138992 86960
rect 139032 86920 139041 86960
rect 79415 86164 79424 86204
rect 79464 86164 79506 86204
rect 79546 86164 79588 86204
rect 79628 86164 79670 86204
rect 79710 86164 79752 86204
rect 79792 86164 79801 86204
rect 94535 86164 94544 86204
rect 94584 86164 94626 86204
rect 94666 86164 94708 86204
rect 94748 86164 94790 86204
rect 94830 86164 94872 86204
rect 94912 86164 94921 86204
rect 109655 86164 109664 86204
rect 109704 86164 109746 86204
rect 109786 86164 109828 86204
rect 109868 86164 109910 86204
rect 109950 86164 109992 86204
rect 110032 86164 110041 86204
rect 124775 86164 124784 86204
rect 124824 86164 124866 86204
rect 124906 86164 124948 86204
rect 124988 86164 125030 86204
rect 125070 86164 125112 86204
rect 125152 86164 125161 86204
rect 139895 86164 139904 86204
rect 139944 86164 139986 86204
rect 140026 86164 140068 86204
rect 140108 86164 140150 86204
rect 140190 86164 140232 86204
rect 140272 86164 140281 86204
rect 78175 85408 78184 85448
rect 78224 85408 78266 85448
rect 78306 85408 78348 85448
rect 78388 85408 78430 85448
rect 78470 85408 78512 85448
rect 78552 85408 78561 85448
rect 93295 85408 93304 85448
rect 93344 85408 93386 85448
rect 93426 85408 93468 85448
rect 93508 85408 93550 85448
rect 93590 85408 93632 85448
rect 93672 85408 93681 85448
rect 108415 85408 108424 85448
rect 108464 85408 108506 85448
rect 108546 85408 108588 85448
rect 108628 85408 108670 85448
rect 108710 85408 108752 85448
rect 108792 85408 108801 85448
rect 123535 85408 123544 85448
rect 123584 85408 123626 85448
rect 123666 85408 123708 85448
rect 123748 85408 123790 85448
rect 123830 85408 123872 85448
rect 123912 85408 123921 85448
rect 138655 85408 138664 85448
rect 138704 85408 138746 85448
rect 138786 85408 138828 85448
rect 138868 85408 138910 85448
rect 138950 85408 138992 85448
rect 139032 85408 139041 85448
rect 79415 84652 79424 84692
rect 79464 84652 79506 84692
rect 79546 84652 79588 84692
rect 79628 84652 79670 84692
rect 79710 84652 79752 84692
rect 79792 84652 79801 84692
rect 94535 84652 94544 84692
rect 94584 84652 94626 84692
rect 94666 84652 94708 84692
rect 94748 84652 94790 84692
rect 94830 84652 94872 84692
rect 94912 84652 94921 84692
rect 109655 84652 109664 84692
rect 109704 84652 109746 84692
rect 109786 84652 109828 84692
rect 109868 84652 109910 84692
rect 109950 84652 109992 84692
rect 110032 84652 110041 84692
rect 124775 84652 124784 84692
rect 124824 84652 124866 84692
rect 124906 84652 124948 84692
rect 124988 84652 125030 84692
rect 125070 84652 125112 84692
rect 125152 84652 125161 84692
rect 139895 84652 139904 84692
rect 139944 84652 139986 84692
rect 140026 84652 140068 84692
rect 140108 84652 140150 84692
rect 140190 84652 140232 84692
rect 140272 84652 140281 84692
rect 78175 83896 78184 83936
rect 78224 83896 78266 83936
rect 78306 83896 78348 83936
rect 78388 83896 78430 83936
rect 78470 83896 78512 83936
rect 78552 83896 78561 83936
rect 93295 83896 93304 83936
rect 93344 83896 93386 83936
rect 93426 83896 93468 83936
rect 93508 83896 93550 83936
rect 93590 83896 93632 83936
rect 93672 83896 93681 83936
rect 108415 83896 108424 83936
rect 108464 83896 108506 83936
rect 108546 83896 108588 83936
rect 108628 83896 108670 83936
rect 108710 83896 108752 83936
rect 108792 83896 108801 83936
rect 123535 83896 123544 83936
rect 123584 83896 123626 83936
rect 123666 83896 123708 83936
rect 123748 83896 123790 83936
rect 123830 83896 123872 83936
rect 123912 83896 123921 83936
rect 138655 83896 138664 83936
rect 138704 83896 138746 83936
rect 138786 83896 138828 83936
rect 138868 83896 138910 83936
rect 138950 83896 138992 83936
rect 139032 83896 139041 83936
rect 79415 83140 79424 83180
rect 79464 83140 79506 83180
rect 79546 83140 79588 83180
rect 79628 83140 79670 83180
rect 79710 83140 79752 83180
rect 79792 83140 79801 83180
rect 94535 83140 94544 83180
rect 94584 83140 94626 83180
rect 94666 83140 94708 83180
rect 94748 83140 94790 83180
rect 94830 83140 94872 83180
rect 94912 83140 94921 83180
rect 109655 83140 109664 83180
rect 109704 83140 109746 83180
rect 109786 83140 109828 83180
rect 109868 83140 109910 83180
rect 109950 83140 109992 83180
rect 110032 83140 110041 83180
rect 124775 83140 124784 83180
rect 124824 83140 124866 83180
rect 124906 83140 124948 83180
rect 124988 83140 125030 83180
rect 125070 83140 125112 83180
rect 125152 83140 125161 83180
rect 139895 83140 139904 83180
rect 139944 83140 139986 83180
rect 140026 83140 140068 83180
rect 140108 83140 140150 83180
rect 140190 83140 140232 83180
rect 140272 83140 140281 83180
rect 78175 82384 78184 82424
rect 78224 82384 78266 82424
rect 78306 82384 78348 82424
rect 78388 82384 78430 82424
rect 78470 82384 78512 82424
rect 78552 82384 78561 82424
rect 93295 82384 93304 82424
rect 93344 82384 93386 82424
rect 93426 82384 93468 82424
rect 93508 82384 93550 82424
rect 93590 82384 93632 82424
rect 93672 82384 93681 82424
rect 108415 82384 108424 82424
rect 108464 82384 108506 82424
rect 108546 82384 108588 82424
rect 108628 82384 108670 82424
rect 108710 82384 108752 82424
rect 108792 82384 108801 82424
rect 123535 82384 123544 82424
rect 123584 82384 123626 82424
rect 123666 82384 123708 82424
rect 123748 82384 123790 82424
rect 123830 82384 123872 82424
rect 123912 82384 123921 82424
rect 138655 82384 138664 82424
rect 138704 82384 138746 82424
rect 138786 82384 138828 82424
rect 138868 82384 138910 82424
rect 138950 82384 138992 82424
rect 139032 82384 139041 82424
rect 79415 81628 79424 81668
rect 79464 81628 79506 81668
rect 79546 81628 79588 81668
rect 79628 81628 79670 81668
rect 79710 81628 79752 81668
rect 79792 81628 79801 81668
rect 94535 81628 94544 81668
rect 94584 81628 94626 81668
rect 94666 81628 94708 81668
rect 94748 81628 94790 81668
rect 94830 81628 94872 81668
rect 94912 81628 94921 81668
rect 109655 81628 109664 81668
rect 109704 81628 109746 81668
rect 109786 81628 109828 81668
rect 109868 81628 109910 81668
rect 109950 81628 109992 81668
rect 110032 81628 110041 81668
rect 124775 81628 124784 81668
rect 124824 81628 124866 81668
rect 124906 81628 124948 81668
rect 124988 81628 125030 81668
rect 125070 81628 125112 81668
rect 125152 81628 125161 81668
rect 139895 81628 139904 81668
rect 139944 81628 139986 81668
rect 140026 81628 140068 81668
rect 140108 81628 140150 81668
rect 140190 81628 140232 81668
rect 140272 81628 140281 81668
rect 78175 80872 78184 80912
rect 78224 80872 78266 80912
rect 78306 80872 78348 80912
rect 78388 80872 78430 80912
rect 78470 80872 78512 80912
rect 78552 80872 78561 80912
rect 93295 80872 93304 80912
rect 93344 80872 93386 80912
rect 93426 80872 93468 80912
rect 93508 80872 93550 80912
rect 93590 80872 93632 80912
rect 93672 80872 93681 80912
rect 108415 80872 108424 80912
rect 108464 80872 108506 80912
rect 108546 80872 108588 80912
rect 108628 80872 108670 80912
rect 108710 80872 108752 80912
rect 108792 80872 108801 80912
rect 123535 80872 123544 80912
rect 123584 80872 123626 80912
rect 123666 80872 123708 80912
rect 123748 80872 123790 80912
rect 123830 80872 123872 80912
rect 123912 80872 123921 80912
rect 138655 80872 138664 80912
rect 138704 80872 138746 80912
rect 138786 80872 138828 80912
rect 138868 80872 138910 80912
rect 138950 80872 138992 80912
rect 139032 80872 139041 80912
rect 79415 80116 79424 80156
rect 79464 80116 79506 80156
rect 79546 80116 79588 80156
rect 79628 80116 79670 80156
rect 79710 80116 79752 80156
rect 79792 80116 79801 80156
rect 94535 80116 94544 80156
rect 94584 80116 94626 80156
rect 94666 80116 94708 80156
rect 94748 80116 94790 80156
rect 94830 80116 94872 80156
rect 94912 80116 94921 80156
rect 109655 80116 109664 80156
rect 109704 80116 109746 80156
rect 109786 80116 109828 80156
rect 109868 80116 109910 80156
rect 109950 80116 109992 80156
rect 110032 80116 110041 80156
rect 124775 80116 124784 80156
rect 124824 80116 124866 80156
rect 124906 80116 124948 80156
rect 124988 80116 125030 80156
rect 125070 80116 125112 80156
rect 125152 80116 125161 80156
rect 139895 80116 139904 80156
rect 139944 80116 139986 80156
rect 140026 80116 140068 80156
rect 140108 80116 140150 80156
rect 140190 80116 140232 80156
rect 140272 80116 140281 80156
rect 78175 79360 78184 79400
rect 78224 79360 78266 79400
rect 78306 79360 78348 79400
rect 78388 79360 78430 79400
rect 78470 79360 78512 79400
rect 78552 79360 78561 79400
rect 93295 79360 93304 79400
rect 93344 79360 93386 79400
rect 93426 79360 93468 79400
rect 93508 79360 93550 79400
rect 93590 79360 93632 79400
rect 93672 79360 93681 79400
rect 108415 79360 108424 79400
rect 108464 79360 108506 79400
rect 108546 79360 108588 79400
rect 108628 79360 108670 79400
rect 108710 79360 108752 79400
rect 108792 79360 108801 79400
rect 123535 79360 123544 79400
rect 123584 79360 123626 79400
rect 123666 79360 123708 79400
rect 123748 79360 123790 79400
rect 123830 79360 123872 79400
rect 123912 79360 123921 79400
rect 138655 79360 138664 79400
rect 138704 79360 138746 79400
rect 138786 79360 138828 79400
rect 138868 79360 138910 79400
rect 138950 79360 138992 79400
rect 139032 79360 139041 79400
rect 79415 78604 79424 78644
rect 79464 78604 79506 78644
rect 79546 78604 79588 78644
rect 79628 78604 79670 78644
rect 79710 78604 79752 78644
rect 79792 78604 79801 78644
rect 94535 78604 94544 78644
rect 94584 78604 94626 78644
rect 94666 78604 94708 78644
rect 94748 78604 94790 78644
rect 94830 78604 94872 78644
rect 94912 78604 94921 78644
rect 109655 78604 109664 78644
rect 109704 78604 109746 78644
rect 109786 78604 109828 78644
rect 109868 78604 109910 78644
rect 109950 78604 109992 78644
rect 110032 78604 110041 78644
rect 124775 78604 124784 78644
rect 124824 78604 124866 78644
rect 124906 78604 124948 78644
rect 124988 78604 125030 78644
rect 125070 78604 125112 78644
rect 125152 78604 125161 78644
rect 139895 78604 139904 78644
rect 139944 78604 139986 78644
rect 140026 78604 140068 78644
rect 140108 78604 140150 78644
rect 140190 78604 140232 78644
rect 140272 78604 140281 78644
rect 78175 77848 78184 77888
rect 78224 77848 78266 77888
rect 78306 77848 78348 77888
rect 78388 77848 78430 77888
rect 78470 77848 78512 77888
rect 78552 77848 78561 77888
rect 93295 77848 93304 77888
rect 93344 77848 93386 77888
rect 93426 77848 93468 77888
rect 93508 77848 93550 77888
rect 93590 77848 93632 77888
rect 93672 77848 93681 77888
rect 108415 77848 108424 77888
rect 108464 77848 108506 77888
rect 108546 77848 108588 77888
rect 108628 77848 108670 77888
rect 108710 77848 108752 77888
rect 108792 77848 108801 77888
rect 123535 77848 123544 77888
rect 123584 77848 123626 77888
rect 123666 77848 123708 77888
rect 123748 77848 123790 77888
rect 123830 77848 123872 77888
rect 123912 77848 123921 77888
rect 138655 77848 138664 77888
rect 138704 77848 138746 77888
rect 138786 77848 138828 77888
rect 138868 77848 138910 77888
rect 138950 77848 138992 77888
rect 139032 77848 139041 77888
rect 79415 77092 79424 77132
rect 79464 77092 79506 77132
rect 79546 77092 79588 77132
rect 79628 77092 79670 77132
rect 79710 77092 79752 77132
rect 79792 77092 79801 77132
rect 94535 77092 94544 77132
rect 94584 77092 94626 77132
rect 94666 77092 94708 77132
rect 94748 77092 94790 77132
rect 94830 77092 94872 77132
rect 94912 77092 94921 77132
rect 109655 77092 109664 77132
rect 109704 77092 109746 77132
rect 109786 77092 109828 77132
rect 109868 77092 109910 77132
rect 109950 77092 109992 77132
rect 110032 77092 110041 77132
rect 124775 77092 124784 77132
rect 124824 77092 124866 77132
rect 124906 77092 124948 77132
rect 124988 77092 125030 77132
rect 125070 77092 125112 77132
rect 125152 77092 125161 77132
rect 139895 77092 139904 77132
rect 139944 77092 139986 77132
rect 140026 77092 140068 77132
rect 140108 77092 140150 77132
rect 140190 77092 140232 77132
rect 140272 77092 140281 77132
rect 78175 76336 78184 76376
rect 78224 76336 78266 76376
rect 78306 76336 78348 76376
rect 78388 76336 78430 76376
rect 78470 76336 78512 76376
rect 78552 76336 78561 76376
rect 93295 76336 93304 76376
rect 93344 76336 93386 76376
rect 93426 76336 93468 76376
rect 93508 76336 93550 76376
rect 93590 76336 93632 76376
rect 93672 76336 93681 76376
rect 108415 76336 108424 76376
rect 108464 76336 108506 76376
rect 108546 76336 108588 76376
rect 108628 76336 108670 76376
rect 108710 76336 108752 76376
rect 108792 76336 108801 76376
rect 123535 76336 123544 76376
rect 123584 76336 123626 76376
rect 123666 76336 123708 76376
rect 123748 76336 123790 76376
rect 123830 76336 123872 76376
rect 123912 76336 123921 76376
rect 138655 76336 138664 76376
rect 138704 76336 138746 76376
rect 138786 76336 138828 76376
rect 138868 76336 138910 76376
rect 138950 76336 138992 76376
rect 139032 76336 139041 76376
rect 79415 75580 79424 75620
rect 79464 75580 79506 75620
rect 79546 75580 79588 75620
rect 79628 75580 79670 75620
rect 79710 75580 79752 75620
rect 79792 75580 79801 75620
rect 94535 75580 94544 75620
rect 94584 75580 94626 75620
rect 94666 75580 94708 75620
rect 94748 75580 94790 75620
rect 94830 75580 94872 75620
rect 94912 75580 94921 75620
rect 109655 75580 109664 75620
rect 109704 75580 109746 75620
rect 109786 75580 109828 75620
rect 109868 75580 109910 75620
rect 109950 75580 109992 75620
rect 110032 75580 110041 75620
rect 124775 75580 124784 75620
rect 124824 75580 124866 75620
rect 124906 75580 124948 75620
rect 124988 75580 125030 75620
rect 125070 75580 125112 75620
rect 125152 75580 125161 75620
rect 139895 75580 139904 75620
rect 139944 75580 139986 75620
rect 140026 75580 140068 75620
rect 140108 75580 140150 75620
rect 140190 75580 140232 75620
rect 140272 75580 140281 75620
rect 148195 72388 148204 72428
rect 148244 72388 148340 72428
rect 148300 72344 148340 72388
rect 148300 72304 160032 72344
rect 64099 71968 64108 72008
rect 64148 71968 67700 72008
rect 67660 71252 67700 71968
rect 90691 71252 90749 71253
rect 67660 71212 90700 71252
rect 90740 71212 90749 71252
rect 90691 71211 90749 71212
rect 92131 71252 92189 71253
rect 92131 71212 92140 71252
rect 92180 71212 93772 71252
rect 93812 71212 93821 71252
rect 92131 71211 92189 71212
rect 71980 64156 73324 64196
rect 73364 64156 73373 64196
rect 71980 63971 72020 64156
<< via3 >>
rect 79424 148156 79464 148196
rect 79506 148156 79546 148196
rect 79588 148156 79628 148196
rect 79670 148156 79710 148196
rect 79752 148156 79792 148196
rect 94544 148156 94584 148196
rect 94626 148156 94666 148196
rect 94708 148156 94748 148196
rect 94790 148156 94830 148196
rect 94872 148156 94912 148196
rect 109664 148156 109704 148196
rect 109746 148156 109786 148196
rect 109828 148156 109868 148196
rect 109910 148156 109950 148196
rect 109992 148156 110032 148196
rect 124784 148156 124824 148196
rect 124866 148156 124906 148196
rect 124948 148156 124988 148196
rect 125030 148156 125070 148196
rect 125112 148156 125152 148196
rect 139904 148156 139944 148196
rect 139986 148156 140026 148196
rect 140068 148156 140108 148196
rect 140150 148156 140190 148196
rect 140232 148156 140272 148196
rect 78184 147400 78224 147440
rect 78266 147400 78306 147440
rect 78348 147400 78388 147440
rect 78430 147400 78470 147440
rect 78512 147400 78552 147440
rect 93304 147400 93344 147440
rect 93386 147400 93426 147440
rect 93468 147400 93508 147440
rect 93550 147400 93590 147440
rect 93632 147400 93672 147440
rect 108424 147400 108464 147440
rect 108506 147400 108546 147440
rect 108588 147400 108628 147440
rect 108670 147400 108710 147440
rect 108752 147400 108792 147440
rect 123544 147400 123584 147440
rect 123626 147400 123666 147440
rect 123708 147400 123748 147440
rect 123790 147400 123830 147440
rect 123872 147400 123912 147440
rect 138664 147400 138704 147440
rect 138746 147400 138786 147440
rect 138828 147400 138868 147440
rect 138910 147400 138950 147440
rect 138992 147400 139032 147440
rect 79424 146644 79464 146684
rect 79506 146644 79546 146684
rect 79588 146644 79628 146684
rect 79670 146644 79710 146684
rect 79752 146644 79792 146684
rect 94544 146644 94584 146684
rect 94626 146644 94666 146684
rect 94708 146644 94748 146684
rect 94790 146644 94830 146684
rect 94872 146644 94912 146684
rect 109664 146644 109704 146684
rect 109746 146644 109786 146684
rect 109828 146644 109868 146684
rect 109910 146644 109950 146684
rect 109992 146644 110032 146684
rect 124784 146644 124824 146684
rect 124866 146644 124906 146684
rect 124948 146644 124988 146684
rect 125030 146644 125070 146684
rect 125112 146644 125152 146684
rect 139904 146644 139944 146684
rect 139986 146644 140026 146684
rect 140068 146644 140108 146684
rect 140150 146644 140190 146684
rect 140232 146644 140272 146684
rect 78184 145888 78224 145928
rect 78266 145888 78306 145928
rect 78348 145888 78388 145928
rect 78430 145888 78470 145928
rect 78512 145888 78552 145928
rect 93304 145888 93344 145928
rect 93386 145888 93426 145928
rect 93468 145888 93508 145928
rect 93550 145888 93590 145928
rect 93632 145888 93672 145928
rect 108424 145888 108464 145928
rect 108506 145888 108546 145928
rect 108588 145888 108628 145928
rect 108670 145888 108710 145928
rect 108752 145888 108792 145928
rect 123544 145888 123584 145928
rect 123626 145888 123666 145928
rect 123708 145888 123748 145928
rect 123790 145888 123830 145928
rect 123872 145888 123912 145928
rect 138664 145888 138704 145928
rect 138746 145888 138786 145928
rect 138828 145888 138868 145928
rect 138910 145888 138950 145928
rect 138992 145888 139032 145928
rect 79424 145132 79464 145172
rect 79506 145132 79546 145172
rect 79588 145132 79628 145172
rect 79670 145132 79710 145172
rect 79752 145132 79792 145172
rect 94544 145132 94584 145172
rect 94626 145132 94666 145172
rect 94708 145132 94748 145172
rect 94790 145132 94830 145172
rect 94872 145132 94912 145172
rect 109664 145132 109704 145172
rect 109746 145132 109786 145172
rect 109828 145132 109868 145172
rect 109910 145132 109950 145172
rect 109992 145132 110032 145172
rect 124784 145132 124824 145172
rect 124866 145132 124906 145172
rect 124948 145132 124988 145172
rect 125030 145132 125070 145172
rect 125112 145132 125152 145172
rect 139904 145132 139944 145172
rect 139986 145132 140026 145172
rect 140068 145132 140108 145172
rect 140150 145132 140190 145172
rect 140232 145132 140272 145172
rect 78184 144376 78224 144416
rect 78266 144376 78306 144416
rect 78348 144376 78388 144416
rect 78430 144376 78470 144416
rect 78512 144376 78552 144416
rect 93304 144376 93344 144416
rect 93386 144376 93426 144416
rect 93468 144376 93508 144416
rect 93550 144376 93590 144416
rect 93632 144376 93672 144416
rect 108424 144376 108464 144416
rect 108506 144376 108546 144416
rect 108588 144376 108628 144416
rect 108670 144376 108710 144416
rect 108752 144376 108792 144416
rect 123544 144376 123584 144416
rect 123626 144376 123666 144416
rect 123708 144376 123748 144416
rect 123790 144376 123830 144416
rect 123872 144376 123912 144416
rect 138664 144376 138704 144416
rect 138746 144376 138786 144416
rect 138828 144376 138868 144416
rect 138910 144376 138950 144416
rect 138992 144376 139032 144416
rect 79424 143620 79464 143660
rect 79506 143620 79546 143660
rect 79588 143620 79628 143660
rect 79670 143620 79710 143660
rect 79752 143620 79792 143660
rect 94544 143620 94584 143660
rect 94626 143620 94666 143660
rect 94708 143620 94748 143660
rect 94790 143620 94830 143660
rect 94872 143620 94912 143660
rect 109664 143620 109704 143660
rect 109746 143620 109786 143660
rect 109828 143620 109868 143660
rect 109910 143620 109950 143660
rect 109992 143620 110032 143660
rect 124784 143620 124824 143660
rect 124866 143620 124906 143660
rect 124948 143620 124988 143660
rect 125030 143620 125070 143660
rect 125112 143620 125152 143660
rect 139904 143620 139944 143660
rect 139986 143620 140026 143660
rect 140068 143620 140108 143660
rect 140150 143620 140190 143660
rect 140232 143620 140272 143660
rect 78184 142864 78224 142904
rect 78266 142864 78306 142904
rect 78348 142864 78388 142904
rect 78430 142864 78470 142904
rect 78512 142864 78552 142904
rect 93304 142864 93344 142904
rect 93386 142864 93426 142904
rect 93468 142864 93508 142904
rect 93550 142864 93590 142904
rect 93632 142864 93672 142904
rect 108424 142864 108464 142904
rect 108506 142864 108546 142904
rect 108588 142864 108628 142904
rect 108670 142864 108710 142904
rect 108752 142864 108792 142904
rect 123544 142864 123584 142904
rect 123626 142864 123666 142904
rect 123708 142864 123748 142904
rect 123790 142864 123830 142904
rect 123872 142864 123912 142904
rect 138664 142864 138704 142904
rect 138746 142864 138786 142904
rect 138828 142864 138868 142904
rect 138910 142864 138950 142904
rect 138992 142864 139032 142904
rect 79424 142108 79464 142148
rect 79506 142108 79546 142148
rect 79588 142108 79628 142148
rect 79670 142108 79710 142148
rect 79752 142108 79792 142148
rect 94544 142108 94584 142148
rect 94626 142108 94666 142148
rect 94708 142108 94748 142148
rect 94790 142108 94830 142148
rect 94872 142108 94912 142148
rect 109664 142108 109704 142148
rect 109746 142108 109786 142148
rect 109828 142108 109868 142148
rect 109910 142108 109950 142148
rect 109992 142108 110032 142148
rect 124784 142108 124824 142148
rect 124866 142108 124906 142148
rect 124948 142108 124988 142148
rect 125030 142108 125070 142148
rect 125112 142108 125152 142148
rect 139904 142108 139944 142148
rect 139986 142108 140026 142148
rect 140068 142108 140108 142148
rect 140150 142108 140190 142148
rect 140232 142108 140272 142148
rect 78184 141352 78224 141392
rect 78266 141352 78306 141392
rect 78348 141352 78388 141392
rect 78430 141352 78470 141392
rect 78512 141352 78552 141392
rect 93304 141352 93344 141392
rect 93386 141352 93426 141392
rect 93468 141352 93508 141392
rect 93550 141352 93590 141392
rect 93632 141352 93672 141392
rect 108424 141352 108464 141392
rect 108506 141352 108546 141392
rect 108588 141352 108628 141392
rect 108670 141352 108710 141392
rect 108752 141352 108792 141392
rect 123544 141352 123584 141392
rect 123626 141352 123666 141392
rect 123708 141352 123748 141392
rect 123790 141352 123830 141392
rect 123872 141352 123912 141392
rect 138664 141352 138704 141392
rect 138746 141352 138786 141392
rect 138828 141352 138868 141392
rect 138910 141352 138950 141392
rect 138992 141352 139032 141392
rect 79424 140596 79464 140636
rect 79506 140596 79546 140636
rect 79588 140596 79628 140636
rect 79670 140596 79710 140636
rect 79752 140596 79792 140636
rect 94544 140596 94584 140636
rect 94626 140596 94666 140636
rect 94708 140596 94748 140636
rect 94790 140596 94830 140636
rect 94872 140596 94912 140636
rect 109664 140596 109704 140636
rect 109746 140596 109786 140636
rect 109828 140596 109868 140636
rect 109910 140596 109950 140636
rect 109992 140596 110032 140636
rect 124784 140596 124824 140636
rect 124866 140596 124906 140636
rect 124948 140596 124988 140636
rect 125030 140596 125070 140636
rect 125112 140596 125152 140636
rect 139904 140596 139944 140636
rect 139986 140596 140026 140636
rect 140068 140596 140108 140636
rect 140150 140596 140190 140636
rect 140232 140596 140272 140636
rect 78184 139840 78224 139880
rect 78266 139840 78306 139880
rect 78348 139840 78388 139880
rect 78430 139840 78470 139880
rect 78512 139840 78552 139880
rect 93304 139840 93344 139880
rect 93386 139840 93426 139880
rect 93468 139840 93508 139880
rect 93550 139840 93590 139880
rect 93632 139840 93672 139880
rect 108424 139840 108464 139880
rect 108506 139840 108546 139880
rect 108588 139840 108628 139880
rect 108670 139840 108710 139880
rect 108752 139840 108792 139880
rect 123544 139840 123584 139880
rect 123626 139840 123666 139880
rect 123708 139840 123748 139880
rect 123790 139840 123830 139880
rect 123872 139840 123912 139880
rect 138664 139840 138704 139880
rect 138746 139840 138786 139880
rect 138828 139840 138868 139880
rect 138910 139840 138950 139880
rect 138992 139840 139032 139880
rect 79424 139084 79464 139124
rect 79506 139084 79546 139124
rect 79588 139084 79628 139124
rect 79670 139084 79710 139124
rect 79752 139084 79792 139124
rect 94544 139084 94584 139124
rect 94626 139084 94666 139124
rect 94708 139084 94748 139124
rect 94790 139084 94830 139124
rect 94872 139084 94912 139124
rect 109664 139084 109704 139124
rect 109746 139084 109786 139124
rect 109828 139084 109868 139124
rect 109910 139084 109950 139124
rect 109992 139084 110032 139124
rect 124784 139084 124824 139124
rect 124866 139084 124906 139124
rect 124948 139084 124988 139124
rect 125030 139084 125070 139124
rect 125112 139084 125152 139124
rect 139904 139084 139944 139124
rect 139986 139084 140026 139124
rect 140068 139084 140108 139124
rect 140150 139084 140190 139124
rect 140232 139084 140272 139124
rect 78184 138328 78224 138368
rect 78266 138328 78306 138368
rect 78348 138328 78388 138368
rect 78430 138328 78470 138368
rect 78512 138328 78552 138368
rect 93304 138328 93344 138368
rect 93386 138328 93426 138368
rect 93468 138328 93508 138368
rect 93550 138328 93590 138368
rect 93632 138328 93672 138368
rect 108424 138328 108464 138368
rect 108506 138328 108546 138368
rect 108588 138328 108628 138368
rect 108670 138328 108710 138368
rect 108752 138328 108792 138368
rect 123544 138328 123584 138368
rect 123626 138328 123666 138368
rect 123708 138328 123748 138368
rect 123790 138328 123830 138368
rect 123872 138328 123912 138368
rect 138664 138328 138704 138368
rect 138746 138328 138786 138368
rect 138828 138328 138868 138368
rect 138910 138328 138950 138368
rect 138992 138328 139032 138368
rect 79424 137572 79464 137612
rect 79506 137572 79546 137612
rect 79588 137572 79628 137612
rect 79670 137572 79710 137612
rect 79752 137572 79792 137612
rect 94544 137572 94584 137612
rect 94626 137572 94666 137612
rect 94708 137572 94748 137612
rect 94790 137572 94830 137612
rect 94872 137572 94912 137612
rect 109664 137572 109704 137612
rect 109746 137572 109786 137612
rect 109828 137572 109868 137612
rect 109910 137572 109950 137612
rect 109992 137572 110032 137612
rect 124784 137572 124824 137612
rect 124866 137572 124906 137612
rect 124948 137572 124988 137612
rect 125030 137572 125070 137612
rect 125112 137572 125152 137612
rect 139904 137572 139944 137612
rect 139986 137572 140026 137612
rect 140068 137572 140108 137612
rect 140150 137572 140190 137612
rect 140232 137572 140272 137612
rect 78184 136816 78224 136856
rect 78266 136816 78306 136856
rect 78348 136816 78388 136856
rect 78430 136816 78470 136856
rect 78512 136816 78552 136856
rect 93304 136816 93344 136856
rect 93386 136816 93426 136856
rect 93468 136816 93508 136856
rect 93550 136816 93590 136856
rect 93632 136816 93672 136856
rect 108424 136816 108464 136856
rect 108506 136816 108546 136856
rect 108588 136816 108628 136856
rect 108670 136816 108710 136856
rect 108752 136816 108792 136856
rect 123544 136816 123584 136856
rect 123626 136816 123666 136856
rect 123708 136816 123748 136856
rect 123790 136816 123830 136856
rect 123872 136816 123912 136856
rect 138664 136816 138704 136856
rect 138746 136816 138786 136856
rect 138828 136816 138868 136856
rect 138910 136816 138950 136856
rect 138992 136816 139032 136856
rect 79424 136060 79464 136100
rect 79506 136060 79546 136100
rect 79588 136060 79628 136100
rect 79670 136060 79710 136100
rect 79752 136060 79792 136100
rect 94544 136060 94584 136100
rect 94626 136060 94666 136100
rect 94708 136060 94748 136100
rect 94790 136060 94830 136100
rect 94872 136060 94912 136100
rect 109664 136060 109704 136100
rect 109746 136060 109786 136100
rect 109828 136060 109868 136100
rect 109910 136060 109950 136100
rect 109992 136060 110032 136100
rect 124784 136060 124824 136100
rect 124866 136060 124906 136100
rect 124948 136060 124988 136100
rect 125030 136060 125070 136100
rect 125112 136060 125152 136100
rect 139904 136060 139944 136100
rect 139986 136060 140026 136100
rect 140068 136060 140108 136100
rect 140150 136060 140190 136100
rect 140232 136060 140272 136100
rect 78184 135304 78224 135344
rect 78266 135304 78306 135344
rect 78348 135304 78388 135344
rect 78430 135304 78470 135344
rect 78512 135304 78552 135344
rect 93304 135304 93344 135344
rect 93386 135304 93426 135344
rect 93468 135304 93508 135344
rect 93550 135304 93590 135344
rect 93632 135304 93672 135344
rect 108424 135304 108464 135344
rect 108506 135304 108546 135344
rect 108588 135304 108628 135344
rect 108670 135304 108710 135344
rect 108752 135304 108792 135344
rect 123544 135304 123584 135344
rect 123626 135304 123666 135344
rect 123708 135304 123748 135344
rect 123790 135304 123830 135344
rect 123872 135304 123912 135344
rect 138664 135304 138704 135344
rect 138746 135304 138786 135344
rect 138828 135304 138868 135344
rect 138910 135304 138950 135344
rect 138992 135304 139032 135344
rect 79424 134548 79464 134588
rect 79506 134548 79546 134588
rect 79588 134548 79628 134588
rect 79670 134548 79710 134588
rect 79752 134548 79792 134588
rect 94544 134548 94584 134588
rect 94626 134548 94666 134588
rect 94708 134548 94748 134588
rect 94790 134548 94830 134588
rect 94872 134548 94912 134588
rect 109664 134548 109704 134588
rect 109746 134548 109786 134588
rect 109828 134548 109868 134588
rect 109910 134548 109950 134588
rect 109992 134548 110032 134588
rect 124784 134548 124824 134588
rect 124866 134548 124906 134588
rect 124948 134548 124988 134588
rect 125030 134548 125070 134588
rect 125112 134548 125152 134588
rect 139904 134548 139944 134588
rect 139986 134548 140026 134588
rect 140068 134548 140108 134588
rect 140150 134548 140190 134588
rect 140232 134548 140272 134588
rect 78184 133792 78224 133832
rect 78266 133792 78306 133832
rect 78348 133792 78388 133832
rect 78430 133792 78470 133832
rect 78512 133792 78552 133832
rect 93304 133792 93344 133832
rect 93386 133792 93426 133832
rect 93468 133792 93508 133832
rect 93550 133792 93590 133832
rect 93632 133792 93672 133832
rect 108424 133792 108464 133832
rect 108506 133792 108546 133832
rect 108588 133792 108628 133832
rect 108670 133792 108710 133832
rect 108752 133792 108792 133832
rect 123544 133792 123584 133832
rect 123626 133792 123666 133832
rect 123708 133792 123748 133832
rect 123790 133792 123830 133832
rect 123872 133792 123912 133832
rect 138664 133792 138704 133832
rect 138746 133792 138786 133832
rect 138828 133792 138868 133832
rect 138910 133792 138950 133832
rect 138992 133792 139032 133832
rect 79424 133036 79464 133076
rect 79506 133036 79546 133076
rect 79588 133036 79628 133076
rect 79670 133036 79710 133076
rect 79752 133036 79792 133076
rect 94544 133036 94584 133076
rect 94626 133036 94666 133076
rect 94708 133036 94748 133076
rect 94790 133036 94830 133076
rect 94872 133036 94912 133076
rect 109664 133036 109704 133076
rect 109746 133036 109786 133076
rect 109828 133036 109868 133076
rect 109910 133036 109950 133076
rect 109992 133036 110032 133076
rect 124784 133036 124824 133076
rect 124866 133036 124906 133076
rect 124948 133036 124988 133076
rect 125030 133036 125070 133076
rect 125112 133036 125152 133076
rect 139904 133036 139944 133076
rect 139986 133036 140026 133076
rect 140068 133036 140108 133076
rect 140150 133036 140190 133076
rect 140232 133036 140272 133076
rect 78184 132280 78224 132320
rect 78266 132280 78306 132320
rect 78348 132280 78388 132320
rect 78430 132280 78470 132320
rect 78512 132280 78552 132320
rect 93304 132280 93344 132320
rect 93386 132280 93426 132320
rect 93468 132280 93508 132320
rect 93550 132280 93590 132320
rect 93632 132280 93672 132320
rect 108424 132280 108464 132320
rect 108506 132280 108546 132320
rect 108588 132280 108628 132320
rect 108670 132280 108710 132320
rect 108752 132280 108792 132320
rect 123544 132280 123584 132320
rect 123626 132280 123666 132320
rect 123708 132280 123748 132320
rect 123790 132280 123830 132320
rect 123872 132280 123912 132320
rect 138664 132280 138704 132320
rect 138746 132280 138786 132320
rect 138828 132280 138868 132320
rect 138910 132280 138950 132320
rect 138992 132280 139032 132320
rect 79424 131524 79464 131564
rect 79506 131524 79546 131564
rect 79588 131524 79628 131564
rect 79670 131524 79710 131564
rect 79752 131524 79792 131564
rect 94544 131524 94584 131564
rect 94626 131524 94666 131564
rect 94708 131524 94748 131564
rect 94790 131524 94830 131564
rect 94872 131524 94912 131564
rect 109664 131524 109704 131564
rect 109746 131524 109786 131564
rect 109828 131524 109868 131564
rect 109910 131524 109950 131564
rect 109992 131524 110032 131564
rect 124784 131524 124824 131564
rect 124866 131524 124906 131564
rect 124948 131524 124988 131564
rect 125030 131524 125070 131564
rect 125112 131524 125152 131564
rect 139904 131524 139944 131564
rect 139986 131524 140026 131564
rect 140068 131524 140108 131564
rect 140150 131524 140190 131564
rect 140232 131524 140272 131564
rect 78184 130768 78224 130808
rect 78266 130768 78306 130808
rect 78348 130768 78388 130808
rect 78430 130768 78470 130808
rect 78512 130768 78552 130808
rect 93304 130768 93344 130808
rect 93386 130768 93426 130808
rect 93468 130768 93508 130808
rect 93550 130768 93590 130808
rect 93632 130768 93672 130808
rect 108424 130768 108464 130808
rect 108506 130768 108546 130808
rect 108588 130768 108628 130808
rect 108670 130768 108710 130808
rect 108752 130768 108792 130808
rect 123544 130768 123584 130808
rect 123626 130768 123666 130808
rect 123708 130768 123748 130808
rect 123790 130768 123830 130808
rect 123872 130768 123912 130808
rect 138664 130768 138704 130808
rect 138746 130768 138786 130808
rect 138828 130768 138868 130808
rect 138910 130768 138950 130808
rect 138992 130768 139032 130808
rect 79424 130012 79464 130052
rect 79506 130012 79546 130052
rect 79588 130012 79628 130052
rect 79670 130012 79710 130052
rect 79752 130012 79792 130052
rect 94544 130012 94584 130052
rect 94626 130012 94666 130052
rect 94708 130012 94748 130052
rect 94790 130012 94830 130052
rect 94872 130012 94912 130052
rect 109664 130012 109704 130052
rect 109746 130012 109786 130052
rect 109828 130012 109868 130052
rect 109910 130012 109950 130052
rect 109992 130012 110032 130052
rect 124784 130012 124824 130052
rect 124866 130012 124906 130052
rect 124948 130012 124988 130052
rect 125030 130012 125070 130052
rect 125112 130012 125152 130052
rect 139904 130012 139944 130052
rect 139986 130012 140026 130052
rect 140068 130012 140108 130052
rect 140150 130012 140190 130052
rect 140232 130012 140272 130052
rect 78184 129256 78224 129296
rect 78266 129256 78306 129296
rect 78348 129256 78388 129296
rect 78430 129256 78470 129296
rect 78512 129256 78552 129296
rect 93304 129256 93344 129296
rect 93386 129256 93426 129296
rect 93468 129256 93508 129296
rect 93550 129256 93590 129296
rect 93632 129256 93672 129296
rect 108424 129256 108464 129296
rect 108506 129256 108546 129296
rect 108588 129256 108628 129296
rect 108670 129256 108710 129296
rect 108752 129256 108792 129296
rect 123544 129256 123584 129296
rect 123626 129256 123666 129296
rect 123708 129256 123748 129296
rect 123790 129256 123830 129296
rect 123872 129256 123912 129296
rect 138664 129256 138704 129296
rect 138746 129256 138786 129296
rect 138828 129256 138868 129296
rect 138910 129256 138950 129296
rect 138992 129256 139032 129296
rect 79424 128500 79464 128540
rect 79506 128500 79546 128540
rect 79588 128500 79628 128540
rect 79670 128500 79710 128540
rect 79752 128500 79792 128540
rect 94544 128500 94584 128540
rect 94626 128500 94666 128540
rect 94708 128500 94748 128540
rect 94790 128500 94830 128540
rect 94872 128500 94912 128540
rect 109664 128500 109704 128540
rect 109746 128500 109786 128540
rect 109828 128500 109868 128540
rect 109910 128500 109950 128540
rect 109992 128500 110032 128540
rect 124784 128500 124824 128540
rect 124866 128500 124906 128540
rect 124948 128500 124988 128540
rect 125030 128500 125070 128540
rect 125112 128500 125152 128540
rect 139904 128500 139944 128540
rect 139986 128500 140026 128540
rect 140068 128500 140108 128540
rect 140150 128500 140190 128540
rect 140232 128500 140272 128540
rect 78184 127744 78224 127784
rect 78266 127744 78306 127784
rect 78348 127744 78388 127784
rect 78430 127744 78470 127784
rect 78512 127744 78552 127784
rect 93304 127744 93344 127784
rect 93386 127744 93426 127784
rect 93468 127744 93508 127784
rect 93550 127744 93590 127784
rect 93632 127744 93672 127784
rect 108424 127744 108464 127784
rect 108506 127744 108546 127784
rect 108588 127744 108628 127784
rect 108670 127744 108710 127784
rect 108752 127744 108792 127784
rect 123544 127744 123584 127784
rect 123626 127744 123666 127784
rect 123708 127744 123748 127784
rect 123790 127744 123830 127784
rect 123872 127744 123912 127784
rect 138664 127744 138704 127784
rect 138746 127744 138786 127784
rect 138828 127744 138868 127784
rect 138910 127744 138950 127784
rect 138992 127744 139032 127784
rect 79424 126988 79464 127028
rect 79506 126988 79546 127028
rect 79588 126988 79628 127028
rect 79670 126988 79710 127028
rect 79752 126988 79792 127028
rect 94544 126988 94584 127028
rect 94626 126988 94666 127028
rect 94708 126988 94748 127028
rect 94790 126988 94830 127028
rect 94872 126988 94912 127028
rect 109664 126988 109704 127028
rect 109746 126988 109786 127028
rect 109828 126988 109868 127028
rect 109910 126988 109950 127028
rect 109992 126988 110032 127028
rect 124784 126988 124824 127028
rect 124866 126988 124906 127028
rect 124948 126988 124988 127028
rect 125030 126988 125070 127028
rect 125112 126988 125152 127028
rect 139904 126988 139944 127028
rect 139986 126988 140026 127028
rect 140068 126988 140108 127028
rect 140150 126988 140190 127028
rect 140232 126988 140272 127028
rect 78184 126232 78224 126272
rect 78266 126232 78306 126272
rect 78348 126232 78388 126272
rect 78430 126232 78470 126272
rect 78512 126232 78552 126272
rect 93304 126232 93344 126272
rect 93386 126232 93426 126272
rect 93468 126232 93508 126272
rect 93550 126232 93590 126272
rect 93632 126232 93672 126272
rect 108424 126232 108464 126272
rect 108506 126232 108546 126272
rect 108588 126232 108628 126272
rect 108670 126232 108710 126272
rect 108752 126232 108792 126272
rect 123544 126232 123584 126272
rect 123626 126232 123666 126272
rect 123708 126232 123748 126272
rect 123790 126232 123830 126272
rect 123872 126232 123912 126272
rect 138664 126232 138704 126272
rect 138746 126232 138786 126272
rect 138828 126232 138868 126272
rect 138910 126232 138950 126272
rect 138992 126232 139032 126272
rect 79424 125476 79464 125516
rect 79506 125476 79546 125516
rect 79588 125476 79628 125516
rect 79670 125476 79710 125516
rect 79752 125476 79792 125516
rect 94544 125476 94584 125516
rect 94626 125476 94666 125516
rect 94708 125476 94748 125516
rect 94790 125476 94830 125516
rect 94872 125476 94912 125516
rect 109664 125476 109704 125516
rect 109746 125476 109786 125516
rect 109828 125476 109868 125516
rect 109910 125476 109950 125516
rect 109992 125476 110032 125516
rect 124784 125476 124824 125516
rect 124866 125476 124906 125516
rect 124948 125476 124988 125516
rect 125030 125476 125070 125516
rect 125112 125476 125152 125516
rect 139904 125476 139944 125516
rect 139986 125476 140026 125516
rect 140068 125476 140108 125516
rect 140150 125476 140190 125516
rect 140232 125476 140272 125516
rect 93772 125224 93812 125264
rect 78184 124720 78224 124760
rect 78266 124720 78306 124760
rect 78348 124720 78388 124760
rect 78430 124720 78470 124760
rect 78512 124720 78552 124760
rect 93304 124720 93344 124760
rect 93386 124720 93426 124760
rect 93468 124720 93508 124760
rect 93550 124720 93590 124760
rect 93632 124720 93672 124760
rect 108424 124720 108464 124760
rect 108506 124720 108546 124760
rect 108588 124720 108628 124760
rect 108670 124720 108710 124760
rect 108752 124720 108792 124760
rect 123544 124720 123584 124760
rect 123626 124720 123666 124760
rect 123708 124720 123748 124760
rect 123790 124720 123830 124760
rect 123872 124720 123912 124760
rect 138664 124720 138704 124760
rect 138746 124720 138786 124760
rect 138828 124720 138868 124760
rect 138910 124720 138950 124760
rect 138992 124720 139032 124760
rect 79424 123964 79464 124004
rect 79506 123964 79546 124004
rect 79588 123964 79628 124004
rect 79670 123964 79710 124004
rect 79752 123964 79792 124004
rect 94544 123964 94584 124004
rect 94626 123964 94666 124004
rect 94708 123964 94748 124004
rect 94790 123964 94830 124004
rect 94872 123964 94912 124004
rect 109664 123964 109704 124004
rect 109746 123964 109786 124004
rect 109828 123964 109868 124004
rect 109910 123964 109950 124004
rect 109992 123964 110032 124004
rect 124784 123964 124824 124004
rect 124866 123964 124906 124004
rect 124948 123964 124988 124004
rect 125030 123964 125070 124004
rect 125112 123964 125152 124004
rect 139904 123964 139944 124004
rect 139986 123964 140026 124004
rect 140068 123964 140108 124004
rect 140150 123964 140190 124004
rect 140232 123964 140272 124004
rect 78184 123208 78224 123248
rect 78266 123208 78306 123248
rect 78348 123208 78388 123248
rect 78430 123208 78470 123248
rect 78512 123208 78552 123248
rect 93304 123208 93344 123248
rect 93386 123208 93426 123248
rect 93468 123208 93508 123248
rect 93550 123208 93590 123248
rect 93632 123208 93672 123248
rect 108424 123208 108464 123248
rect 108506 123208 108546 123248
rect 108588 123208 108628 123248
rect 108670 123208 108710 123248
rect 108752 123208 108792 123248
rect 123544 123208 123584 123248
rect 123626 123208 123666 123248
rect 123708 123208 123748 123248
rect 123790 123208 123830 123248
rect 123872 123208 123912 123248
rect 138664 123208 138704 123248
rect 138746 123208 138786 123248
rect 138828 123208 138868 123248
rect 138910 123208 138950 123248
rect 138992 123208 139032 123248
rect 79424 122452 79464 122492
rect 79506 122452 79546 122492
rect 79588 122452 79628 122492
rect 79670 122452 79710 122492
rect 79752 122452 79792 122492
rect 94544 122452 94584 122492
rect 94626 122452 94666 122492
rect 94708 122452 94748 122492
rect 94790 122452 94830 122492
rect 94872 122452 94912 122492
rect 109664 122452 109704 122492
rect 109746 122452 109786 122492
rect 109828 122452 109868 122492
rect 109910 122452 109950 122492
rect 109992 122452 110032 122492
rect 124784 122452 124824 122492
rect 124866 122452 124906 122492
rect 124948 122452 124988 122492
rect 125030 122452 125070 122492
rect 125112 122452 125152 122492
rect 139904 122452 139944 122492
rect 139986 122452 140026 122492
rect 140068 122452 140108 122492
rect 140150 122452 140190 122492
rect 140232 122452 140272 122492
rect 93772 122368 93812 122408
rect 78184 121696 78224 121736
rect 78266 121696 78306 121736
rect 78348 121696 78388 121736
rect 78430 121696 78470 121736
rect 78512 121696 78552 121736
rect 93304 121696 93344 121736
rect 93386 121696 93426 121736
rect 93468 121696 93508 121736
rect 93550 121696 93590 121736
rect 93632 121696 93672 121736
rect 108424 121696 108464 121736
rect 108506 121696 108546 121736
rect 108588 121696 108628 121736
rect 108670 121696 108710 121736
rect 108752 121696 108792 121736
rect 123544 121696 123584 121736
rect 123626 121696 123666 121736
rect 123708 121696 123748 121736
rect 123790 121696 123830 121736
rect 123872 121696 123912 121736
rect 138664 121696 138704 121736
rect 138746 121696 138786 121736
rect 138828 121696 138868 121736
rect 138910 121696 138950 121736
rect 138992 121696 139032 121736
rect 79424 120940 79464 120980
rect 79506 120940 79546 120980
rect 79588 120940 79628 120980
rect 79670 120940 79710 120980
rect 79752 120940 79792 120980
rect 94544 120940 94584 120980
rect 94626 120940 94666 120980
rect 94708 120940 94748 120980
rect 94790 120940 94830 120980
rect 94872 120940 94912 120980
rect 109664 120940 109704 120980
rect 109746 120940 109786 120980
rect 109828 120940 109868 120980
rect 109910 120940 109950 120980
rect 109992 120940 110032 120980
rect 124784 120940 124824 120980
rect 124866 120940 124906 120980
rect 124948 120940 124988 120980
rect 125030 120940 125070 120980
rect 125112 120940 125152 120980
rect 139904 120940 139944 120980
rect 139986 120940 140026 120980
rect 140068 120940 140108 120980
rect 140150 120940 140190 120980
rect 140232 120940 140272 120980
rect 78184 120184 78224 120224
rect 78266 120184 78306 120224
rect 78348 120184 78388 120224
rect 78430 120184 78470 120224
rect 78512 120184 78552 120224
rect 93304 120184 93344 120224
rect 93386 120184 93426 120224
rect 93468 120184 93508 120224
rect 93550 120184 93590 120224
rect 93632 120184 93672 120224
rect 108424 120184 108464 120224
rect 108506 120184 108546 120224
rect 108588 120184 108628 120224
rect 108670 120184 108710 120224
rect 108752 120184 108792 120224
rect 123544 120184 123584 120224
rect 123626 120184 123666 120224
rect 123708 120184 123748 120224
rect 123790 120184 123830 120224
rect 123872 120184 123912 120224
rect 138664 120184 138704 120224
rect 138746 120184 138786 120224
rect 138828 120184 138868 120224
rect 138910 120184 138950 120224
rect 138992 120184 139032 120224
rect 79424 119428 79464 119468
rect 79506 119428 79546 119468
rect 79588 119428 79628 119468
rect 79670 119428 79710 119468
rect 79752 119428 79792 119468
rect 94544 119428 94584 119468
rect 94626 119428 94666 119468
rect 94708 119428 94748 119468
rect 94790 119428 94830 119468
rect 94872 119428 94912 119468
rect 109664 119428 109704 119468
rect 109746 119428 109786 119468
rect 109828 119428 109868 119468
rect 109910 119428 109950 119468
rect 109992 119428 110032 119468
rect 124784 119428 124824 119468
rect 124866 119428 124906 119468
rect 124948 119428 124988 119468
rect 125030 119428 125070 119468
rect 125112 119428 125152 119468
rect 139904 119428 139944 119468
rect 139986 119428 140026 119468
rect 140068 119428 140108 119468
rect 140150 119428 140190 119468
rect 140232 119428 140272 119468
rect 78184 118672 78224 118712
rect 78266 118672 78306 118712
rect 78348 118672 78388 118712
rect 78430 118672 78470 118712
rect 78512 118672 78552 118712
rect 93304 118672 93344 118712
rect 93386 118672 93426 118712
rect 93468 118672 93508 118712
rect 93550 118672 93590 118712
rect 93632 118672 93672 118712
rect 108424 118672 108464 118712
rect 108506 118672 108546 118712
rect 108588 118672 108628 118712
rect 108670 118672 108710 118712
rect 108752 118672 108792 118712
rect 123544 118672 123584 118712
rect 123626 118672 123666 118712
rect 123708 118672 123748 118712
rect 123790 118672 123830 118712
rect 123872 118672 123912 118712
rect 138664 118672 138704 118712
rect 138746 118672 138786 118712
rect 138828 118672 138868 118712
rect 138910 118672 138950 118712
rect 138992 118672 139032 118712
rect 79424 117916 79464 117956
rect 79506 117916 79546 117956
rect 79588 117916 79628 117956
rect 79670 117916 79710 117956
rect 79752 117916 79792 117956
rect 94544 117916 94584 117956
rect 94626 117916 94666 117956
rect 94708 117916 94748 117956
rect 94790 117916 94830 117956
rect 94872 117916 94912 117956
rect 109664 117916 109704 117956
rect 109746 117916 109786 117956
rect 109828 117916 109868 117956
rect 109910 117916 109950 117956
rect 109992 117916 110032 117956
rect 124784 117916 124824 117956
rect 124866 117916 124906 117956
rect 124948 117916 124988 117956
rect 125030 117916 125070 117956
rect 125112 117916 125152 117956
rect 139904 117916 139944 117956
rect 139986 117916 140026 117956
rect 140068 117916 140108 117956
rect 140150 117916 140190 117956
rect 140232 117916 140272 117956
rect 78184 117160 78224 117200
rect 78266 117160 78306 117200
rect 78348 117160 78388 117200
rect 78430 117160 78470 117200
rect 78512 117160 78552 117200
rect 93304 117160 93344 117200
rect 93386 117160 93426 117200
rect 93468 117160 93508 117200
rect 93550 117160 93590 117200
rect 93632 117160 93672 117200
rect 108424 117160 108464 117200
rect 108506 117160 108546 117200
rect 108588 117160 108628 117200
rect 108670 117160 108710 117200
rect 108752 117160 108792 117200
rect 123544 117160 123584 117200
rect 123626 117160 123666 117200
rect 123708 117160 123748 117200
rect 123790 117160 123830 117200
rect 123872 117160 123912 117200
rect 138664 117160 138704 117200
rect 138746 117160 138786 117200
rect 138828 117160 138868 117200
rect 138910 117160 138950 117200
rect 138992 117160 139032 117200
rect 79424 116404 79464 116444
rect 79506 116404 79546 116444
rect 79588 116404 79628 116444
rect 79670 116404 79710 116444
rect 79752 116404 79792 116444
rect 94544 116404 94584 116444
rect 94626 116404 94666 116444
rect 94708 116404 94748 116444
rect 94790 116404 94830 116444
rect 94872 116404 94912 116444
rect 109664 116404 109704 116444
rect 109746 116404 109786 116444
rect 109828 116404 109868 116444
rect 109910 116404 109950 116444
rect 109992 116404 110032 116444
rect 124784 116404 124824 116444
rect 124866 116404 124906 116444
rect 124948 116404 124988 116444
rect 125030 116404 125070 116444
rect 125112 116404 125152 116444
rect 139904 116404 139944 116444
rect 139986 116404 140026 116444
rect 140068 116404 140108 116444
rect 140150 116404 140190 116444
rect 140232 116404 140272 116444
rect 78184 115648 78224 115688
rect 78266 115648 78306 115688
rect 78348 115648 78388 115688
rect 78430 115648 78470 115688
rect 78512 115648 78552 115688
rect 93304 115648 93344 115688
rect 93386 115648 93426 115688
rect 93468 115648 93508 115688
rect 93550 115648 93590 115688
rect 93632 115648 93672 115688
rect 108424 115648 108464 115688
rect 108506 115648 108546 115688
rect 108588 115648 108628 115688
rect 108670 115648 108710 115688
rect 108752 115648 108792 115688
rect 123544 115648 123584 115688
rect 123626 115648 123666 115688
rect 123708 115648 123748 115688
rect 123790 115648 123830 115688
rect 123872 115648 123912 115688
rect 138664 115648 138704 115688
rect 138746 115648 138786 115688
rect 138828 115648 138868 115688
rect 138910 115648 138950 115688
rect 138992 115648 139032 115688
rect 79424 114892 79464 114932
rect 79506 114892 79546 114932
rect 79588 114892 79628 114932
rect 79670 114892 79710 114932
rect 79752 114892 79792 114932
rect 94544 114892 94584 114932
rect 94626 114892 94666 114932
rect 94708 114892 94748 114932
rect 94790 114892 94830 114932
rect 94872 114892 94912 114932
rect 109664 114892 109704 114932
rect 109746 114892 109786 114932
rect 109828 114892 109868 114932
rect 109910 114892 109950 114932
rect 109992 114892 110032 114932
rect 124784 114892 124824 114932
rect 124866 114892 124906 114932
rect 124948 114892 124988 114932
rect 125030 114892 125070 114932
rect 125112 114892 125152 114932
rect 139904 114892 139944 114932
rect 139986 114892 140026 114932
rect 140068 114892 140108 114932
rect 140150 114892 140190 114932
rect 140232 114892 140272 114932
rect 78184 114136 78224 114176
rect 78266 114136 78306 114176
rect 78348 114136 78388 114176
rect 78430 114136 78470 114176
rect 78512 114136 78552 114176
rect 93304 114136 93344 114176
rect 93386 114136 93426 114176
rect 93468 114136 93508 114176
rect 93550 114136 93590 114176
rect 93632 114136 93672 114176
rect 108424 114136 108464 114176
rect 108506 114136 108546 114176
rect 108588 114136 108628 114176
rect 108670 114136 108710 114176
rect 108752 114136 108792 114176
rect 123544 114136 123584 114176
rect 123626 114136 123666 114176
rect 123708 114136 123748 114176
rect 123790 114136 123830 114176
rect 123872 114136 123912 114176
rect 138664 114136 138704 114176
rect 138746 114136 138786 114176
rect 138828 114136 138868 114176
rect 138910 114136 138950 114176
rect 138992 114136 139032 114176
rect 79424 113380 79464 113420
rect 79506 113380 79546 113420
rect 79588 113380 79628 113420
rect 79670 113380 79710 113420
rect 79752 113380 79792 113420
rect 94544 113380 94584 113420
rect 94626 113380 94666 113420
rect 94708 113380 94748 113420
rect 94790 113380 94830 113420
rect 94872 113380 94912 113420
rect 109664 113380 109704 113420
rect 109746 113380 109786 113420
rect 109828 113380 109868 113420
rect 109910 113380 109950 113420
rect 109992 113380 110032 113420
rect 124784 113380 124824 113420
rect 124866 113380 124906 113420
rect 124948 113380 124988 113420
rect 125030 113380 125070 113420
rect 125112 113380 125152 113420
rect 139904 113380 139944 113420
rect 139986 113380 140026 113420
rect 140068 113380 140108 113420
rect 140150 113380 140190 113420
rect 140232 113380 140272 113420
rect 78184 112624 78224 112664
rect 78266 112624 78306 112664
rect 78348 112624 78388 112664
rect 78430 112624 78470 112664
rect 78512 112624 78552 112664
rect 93304 112624 93344 112664
rect 93386 112624 93426 112664
rect 93468 112624 93508 112664
rect 93550 112624 93590 112664
rect 93632 112624 93672 112664
rect 108424 112624 108464 112664
rect 108506 112624 108546 112664
rect 108588 112624 108628 112664
rect 108670 112624 108710 112664
rect 108752 112624 108792 112664
rect 123544 112624 123584 112664
rect 123626 112624 123666 112664
rect 123708 112624 123748 112664
rect 123790 112624 123830 112664
rect 123872 112624 123912 112664
rect 138664 112624 138704 112664
rect 138746 112624 138786 112664
rect 138828 112624 138868 112664
rect 138910 112624 138950 112664
rect 138992 112624 139032 112664
rect 79424 111868 79464 111908
rect 79506 111868 79546 111908
rect 79588 111868 79628 111908
rect 79670 111868 79710 111908
rect 79752 111868 79792 111908
rect 94544 111868 94584 111908
rect 94626 111868 94666 111908
rect 94708 111868 94748 111908
rect 94790 111868 94830 111908
rect 94872 111868 94912 111908
rect 109664 111868 109704 111908
rect 109746 111868 109786 111908
rect 109828 111868 109868 111908
rect 109910 111868 109950 111908
rect 109992 111868 110032 111908
rect 124784 111868 124824 111908
rect 124866 111868 124906 111908
rect 124948 111868 124988 111908
rect 125030 111868 125070 111908
rect 125112 111868 125152 111908
rect 139904 111868 139944 111908
rect 139986 111868 140026 111908
rect 140068 111868 140108 111908
rect 140150 111868 140190 111908
rect 140232 111868 140272 111908
rect 78184 111112 78224 111152
rect 78266 111112 78306 111152
rect 78348 111112 78388 111152
rect 78430 111112 78470 111152
rect 78512 111112 78552 111152
rect 93304 111112 93344 111152
rect 93386 111112 93426 111152
rect 93468 111112 93508 111152
rect 93550 111112 93590 111152
rect 93632 111112 93672 111152
rect 108424 111112 108464 111152
rect 108506 111112 108546 111152
rect 108588 111112 108628 111152
rect 108670 111112 108710 111152
rect 108752 111112 108792 111152
rect 123544 111112 123584 111152
rect 123626 111112 123666 111152
rect 123708 111112 123748 111152
rect 123790 111112 123830 111152
rect 123872 111112 123912 111152
rect 138664 111112 138704 111152
rect 138746 111112 138786 111152
rect 138828 111112 138868 111152
rect 138910 111112 138950 111152
rect 138992 111112 139032 111152
rect 79424 110356 79464 110396
rect 79506 110356 79546 110396
rect 79588 110356 79628 110396
rect 79670 110356 79710 110396
rect 79752 110356 79792 110396
rect 94544 110356 94584 110396
rect 94626 110356 94666 110396
rect 94708 110356 94748 110396
rect 94790 110356 94830 110396
rect 94872 110356 94912 110396
rect 109664 110356 109704 110396
rect 109746 110356 109786 110396
rect 109828 110356 109868 110396
rect 109910 110356 109950 110396
rect 109992 110356 110032 110396
rect 124784 110356 124824 110396
rect 124866 110356 124906 110396
rect 124948 110356 124988 110396
rect 125030 110356 125070 110396
rect 125112 110356 125152 110396
rect 139904 110356 139944 110396
rect 139986 110356 140026 110396
rect 140068 110356 140108 110396
rect 140150 110356 140190 110396
rect 140232 110356 140272 110396
rect 78184 109600 78224 109640
rect 78266 109600 78306 109640
rect 78348 109600 78388 109640
rect 78430 109600 78470 109640
rect 78512 109600 78552 109640
rect 93304 109600 93344 109640
rect 93386 109600 93426 109640
rect 93468 109600 93508 109640
rect 93550 109600 93590 109640
rect 93632 109600 93672 109640
rect 108424 109600 108464 109640
rect 108506 109600 108546 109640
rect 108588 109600 108628 109640
rect 108670 109600 108710 109640
rect 108752 109600 108792 109640
rect 123544 109600 123584 109640
rect 123626 109600 123666 109640
rect 123708 109600 123748 109640
rect 123790 109600 123830 109640
rect 123872 109600 123912 109640
rect 138664 109600 138704 109640
rect 138746 109600 138786 109640
rect 138828 109600 138868 109640
rect 138910 109600 138950 109640
rect 138992 109600 139032 109640
rect 79424 108844 79464 108884
rect 79506 108844 79546 108884
rect 79588 108844 79628 108884
rect 79670 108844 79710 108884
rect 79752 108844 79792 108884
rect 94544 108844 94584 108884
rect 94626 108844 94666 108884
rect 94708 108844 94748 108884
rect 94790 108844 94830 108884
rect 94872 108844 94912 108884
rect 109664 108844 109704 108884
rect 109746 108844 109786 108884
rect 109828 108844 109868 108884
rect 109910 108844 109950 108884
rect 109992 108844 110032 108884
rect 124784 108844 124824 108884
rect 124866 108844 124906 108884
rect 124948 108844 124988 108884
rect 125030 108844 125070 108884
rect 125112 108844 125152 108884
rect 139904 108844 139944 108884
rect 139986 108844 140026 108884
rect 140068 108844 140108 108884
rect 140150 108844 140190 108884
rect 140232 108844 140272 108884
rect 78184 108088 78224 108128
rect 78266 108088 78306 108128
rect 78348 108088 78388 108128
rect 78430 108088 78470 108128
rect 78512 108088 78552 108128
rect 93304 108088 93344 108128
rect 93386 108088 93426 108128
rect 93468 108088 93508 108128
rect 93550 108088 93590 108128
rect 93632 108088 93672 108128
rect 108424 108088 108464 108128
rect 108506 108088 108546 108128
rect 108588 108088 108628 108128
rect 108670 108088 108710 108128
rect 108752 108088 108792 108128
rect 123544 108088 123584 108128
rect 123626 108088 123666 108128
rect 123708 108088 123748 108128
rect 123790 108088 123830 108128
rect 123872 108088 123912 108128
rect 138664 108088 138704 108128
rect 138746 108088 138786 108128
rect 138828 108088 138868 108128
rect 138910 108088 138950 108128
rect 138992 108088 139032 108128
rect 79424 107332 79464 107372
rect 79506 107332 79546 107372
rect 79588 107332 79628 107372
rect 79670 107332 79710 107372
rect 79752 107332 79792 107372
rect 94544 107332 94584 107372
rect 94626 107332 94666 107372
rect 94708 107332 94748 107372
rect 94790 107332 94830 107372
rect 94872 107332 94912 107372
rect 109664 107332 109704 107372
rect 109746 107332 109786 107372
rect 109828 107332 109868 107372
rect 109910 107332 109950 107372
rect 109992 107332 110032 107372
rect 124784 107332 124824 107372
rect 124866 107332 124906 107372
rect 124948 107332 124988 107372
rect 125030 107332 125070 107372
rect 125112 107332 125152 107372
rect 139904 107332 139944 107372
rect 139986 107332 140026 107372
rect 140068 107332 140108 107372
rect 140150 107332 140190 107372
rect 140232 107332 140272 107372
rect 78184 106576 78224 106616
rect 78266 106576 78306 106616
rect 78348 106576 78388 106616
rect 78430 106576 78470 106616
rect 78512 106576 78552 106616
rect 93304 106576 93344 106616
rect 93386 106576 93426 106616
rect 93468 106576 93508 106616
rect 93550 106576 93590 106616
rect 93632 106576 93672 106616
rect 108424 106576 108464 106616
rect 108506 106576 108546 106616
rect 108588 106576 108628 106616
rect 108670 106576 108710 106616
rect 108752 106576 108792 106616
rect 123544 106576 123584 106616
rect 123626 106576 123666 106616
rect 123708 106576 123748 106616
rect 123790 106576 123830 106616
rect 123872 106576 123912 106616
rect 138664 106576 138704 106616
rect 138746 106576 138786 106616
rect 138828 106576 138868 106616
rect 138910 106576 138950 106616
rect 138992 106576 139032 106616
rect 79424 105820 79464 105860
rect 79506 105820 79546 105860
rect 79588 105820 79628 105860
rect 79670 105820 79710 105860
rect 79752 105820 79792 105860
rect 94544 105820 94584 105860
rect 94626 105820 94666 105860
rect 94708 105820 94748 105860
rect 94790 105820 94830 105860
rect 94872 105820 94912 105860
rect 109664 105820 109704 105860
rect 109746 105820 109786 105860
rect 109828 105820 109868 105860
rect 109910 105820 109950 105860
rect 109992 105820 110032 105860
rect 124784 105820 124824 105860
rect 124866 105820 124906 105860
rect 124948 105820 124988 105860
rect 125030 105820 125070 105860
rect 125112 105820 125152 105860
rect 139904 105820 139944 105860
rect 139986 105820 140026 105860
rect 140068 105820 140108 105860
rect 140150 105820 140190 105860
rect 140232 105820 140272 105860
rect 78184 105064 78224 105104
rect 78266 105064 78306 105104
rect 78348 105064 78388 105104
rect 78430 105064 78470 105104
rect 78512 105064 78552 105104
rect 93304 105064 93344 105104
rect 93386 105064 93426 105104
rect 93468 105064 93508 105104
rect 93550 105064 93590 105104
rect 93632 105064 93672 105104
rect 108424 105064 108464 105104
rect 108506 105064 108546 105104
rect 108588 105064 108628 105104
rect 108670 105064 108710 105104
rect 108752 105064 108792 105104
rect 123544 105064 123584 105104
rect 123626 105064 123666 105104
rect 123708 105064 123748 105104
rect 123790 105064 123830 105104
rect 123872 105064 123912 105104
rect 138664 105064 138704 105104
rect 138746 105064 138786 105104
rect 138828 105064 138868 105104
rect 138910 105064 138950 105104
rect 138992 105064 139032 105104
rect 79424 104308 79464 104348
rect 79506 104308 79546 104348
rect 79588 104308 79628 104348
rect 79670 104308 79710 104348
rect 79752 104308 79792 104348
rect 94544 104308 94584 104348
rect 94626 104308 94666 104348
rect 94708 104308 94748 104348
rect 94790 104308 94830 104348
rect 94872 104308 94912 104348
rect 109664 104308 109704 104348
rect 109746 104308 109786 104348
rect 109828 104308 109868 104348
rect 109910 104308 109950 104348
rect 109992 104308 110032 104348
rect 124784 104308 124824 104348
rect 124866 104308 124906 104348
rect 124948 104308 124988 104348
rect 125030 104308 125070 104348
rect 125112 104308 125152 104348
rect 139904 104308 139944 104348
rect 139986 104308 140026 104348
rect 140068 104308 140108 104348
rect 140150 104308 140190 104348
rect 140232 104308 140272 104348
rect 78184 103552 78224 103592
rect 78266 103552 78306 103592
rect 78348 103552 78388 103592
rect 78430 103552 78470 103592
rect 78512 103552 78552 103592
rect 93304 103552 93344 103592
rect 93386 103552 93426 103592
rect 93468 103552 93508 103592
rect 93550 103552 93590 103592
rect 93632 103552 93672 103592
rect 108424 103552 108464 103592
rect 108506 103552 108546 103592
rect 108588 103552 108628 103592
rect 108670 103552 108710 103592
rect 108752 103552 108792 103592
rect 123544 103552 123584 103592
rect 123626 103552 123666 103592
rect 123708 103552 123748 103592
rect 123790 103552 123830 103592
rect 123872 103552 123912 103592
rect 138664 103552 138704 103592
rect 138746 103552 138786 103592
rect 138828 103552 138868 103592
rect 138910 103552 138950 103592
rect 138992 103552 139032 103592
rect 79424 102796 79464 102836
rect 79506 102796 79546 102836
rect 79588 102796 79628 102836
rect 79670 102796 79710 102836
rect 79752 102796 79792 102836
rect 94544 102796 94584 102836
rect 94626 102796 94666 102836
rect 94708 102796 94748 102836
rect 94790 102796 94830 102836
rect 94872 102796 94912 102836
rect 109664 102796 109704 102836
rect 109746 102796 109786 102836
rect 109828 102796 109868 102836
rect 109910 102796 109950 102836
rect 109992 102796 110032 102836
rect 124784 102796 124824 102836
rect 124866 102796 124906 102836
rect 124948 102796 124988 102836
rect 125030 102796 125070 102836
rect 125112 102796 125152 102836
rect 139904 102796 139944 102836
rect 139986 102796 140026 102836
rect 140068 102796 140108 102836
rect 140150 102796 140190 102836
rect 140232 102796 140272 102836
rect 78184 102040 78224 102080
rect 78266 102040 78306 102080
rect 78348 102040 78388 102080
rect 78430 102040 78470 102080
rect 78512 102040 78552 102080
rect 93304 102040 93344 102080
rect 93386 102040 93426 102080
rect 93468 102040 93508 102080
rect 93550 102040 93590 102080
rect 93632 102040 93672 102080
rect 108424 102040 108464 102080
rect 108506 102040 108546 102080
rect 108588 102040 108628 102080
rect 108670 102040 108710 102080
rect 108752 102040 108792 102080
rect 123544 102040 123584 102080
rect 123626 102040 123666 102080
rect 123708 102040 123748 102080
rect 123790 102040 123830 102080
rect 123872 102040 123912 102080
rect 138664 102040 138704 102080
rect 138746 102040 138786 102080
rect 138828 102040 138868 102080
rect 138910 102040 138950 102080
rect 138992 102040 139032 102080
rect 79424 101284 79464 101324
rect 79506 101284 79546 101324
rect 79588 101284 79628 101324
rect 79670 101284 79710 101324
rect 79752 101284 79792 101324
rect 94544 101284 94584 101324
rect 94626 101284 94666 101324
rect 94708 101284 94748 101324
rect 94790 101284 94830 101324
rect 94872 101284 94912 101324
rect 109664 101284 109704 101324
rect 109746 101284 109786 101324
rect 109828 101284 109868 101324
rect 109910 101284 109950 101324
rect 109992 101284 110032 101324
rect 124784 101284 124824 101324
rect 124866 101284 124906 101324
rect 124948 101284 124988 101324
rect 125030 101284 125070 101324
rect 125112 101284 125152 101324
rect 139904 101284 139944 101324
rect 139986 101284 140026 101324
rect 140068 101284 140108 101324
rect 140150 101284 140190 101324
rect 140232 101284 140272 101324
rect 78184 100528 78224 100568
rect 78266 100528 78306 100568
rect 78348 100528 78388 100568
rect 78430 100528 78470 100568
rect 78512 100528 78552 100568
rect 93304 100528 93344 100568
rect 93386 100528 93426 100568
rect 93468 100528 93508 100568
rect 93550 100528 93590 100568
rect 93632 100528 93672 100568
rect 108424 100528 108464 100568
rect 108506 100528 108546 100568
rect 108588 100528 108628 100568
rect 108670 100528 108710 100568
rect 108752 100528 108792 100568
rect 123544 100528 123584 100568
rect 123626 100528 123666 100568
rect 123708 100528 123748 100568
rect 123790 100528 123830 100568
rect 123872 100528 123912 100568
rect 138664 100528 138704 100568
rect 138746 100528 138786 100568
rect 138828 100528 138868 100568
rect 138910 100528 138950 100568
rect 138992 100528 139032 100568
rect 79424 99772 79464 99812
rect 79506 99772 79546 99812
rect 79588 99772 79628 99812
rect 79670 99772 79710 99812
rect 79752 99772 79792 99812
rect 94544 99772 94584 99812
rect 94626 99772 94666 99812
rect 94708 99772 94748 99812
rect 94790 99772 94830 99812
rect 94872 99772 94912 99812
rect 109664 99772 109704 99812
rect 109746 99772 109786 99812
rect 109828 99772 109868 99812
rect 109910 99772 109950 99812
rect 109992 99772 110032 99812
rect 124784 99772 124824 99812
rect 124866 99772 124906 99812
rect 124948 99772 124988 99812
rect 125030 99772 125070 99812
rect 125112 99772 125152 99812
rect 139904 99772 139944 99812
rect 139986 99772 140026 99812
rect 140068 99772 140108 99812
rect 140150 99772 140190 99812
rect 140232 99772 140272 99812
rect 78184 99016 78224 99056
rect 78266 99016 78306 99056
rect 78348 99016 78388 99056
rect 78430 99016 78470 99056
rect 78512 99016 78552 99056
rect 93304 99016 93344 99056
rect 93386 99016 93426 99056
rect 93468 99016 93508 99056
rect 93550 99016 93590 99056
rect 93632 99016 93672 99056
rect 108424 99016 108464 99056
rect 108506 99016 108546 99056
rect 108588 99016 108628 99056
rect 108670 99016 108710 99056
rect 108752 99016 108792 99056
rect 123544 99016 123584 99056
rect 123626 99016 123666 99056
rect 123708 99016 123748 99056
rect 123790 99016 123830 99056
rect 123872 99016 123912 99056
rect 138664 99016 138704 99056
rect 138746 99016 138786 99056
rect 138828 99016 138868 99056
rect 138910 99016 138950 99056
rect 138992 99016 139032 99056
rect 79424 98260 79464 98300
rect 79506 98260 79546 98300
rect 79588 98260 79628 98300
rect 79670 98260 79710 98300
rect 79752 98260 79792 98300
rect 94544 98260 94584 98300
rect 94626 98260 94666 98300
rect 94708 98260 94748 98300
rect 94790 98260 94830 98300
rect 94872 98260 94912 98300
rect 109664 98260 109704 98300
rect 109746 98260 109786 98300
rect 109828 98260 109868 98300
rect 109910 98260 109950 98300
rect 109992 98260 110032 98300
rect 124784 98260 124824 98300
rect 124866 98260 124906 98300
rect 124948 98260 124988 98300
rect 125030 98260 125070 98300
rect 125112 98260 125152 98300
rect 139904 98260 139944 98300
rect 139986 98260 140026 98300
rect 140068 98260 140108 98300
rect 140150 98260 140190 98300
rect 140232 98260 140272 98300
rect 78184 97504 78224 97544
rect 78266 97504 78306 97544
rect 78348 97504 78388 97544
rect 78430 97504 78470 97544
rect 78512 97504 78552 97544
rect 93304 97504 93344 97544
rect 93386 97504 93426 97544
rect 93468 97504 93508 97544
rect 93550 97504 93590 97544
rect 93632 97504 93672 97544
rect 108424 97504 108464 97544
rect 108506 97504 108546 97544
rect 108588 97504 108628 97544
rect 108670 97504 108710 97544
rect 108752 97504 108792 97544
rect 123544 97504 123584 97544
rect 123626 97504 123666 97544
rect 123708 97504 123748 97544
rect 123790 97504 123830 97544
rect 123872 97504 123912 97544
rect 138664 97504 138704 97544
rect 138746 97504 138786 97544
rect 138828 97504 138868 97544
rect 138910 97504 138950 97544
rect 138992 97504 139032 97544
rect 79424 96748 79464 96788
rect 79506 96748 79546 96788
rect 79588 96748 79628 96788
rect 79670 96748 79710 96788
rect 79752 96748 79792 96788
rect 94544 96748 94584 96788
rect 94626 96748 94666 96788
rect 94708 96748 94748 96788
rect 94790 96748 94830 96788
rect 94872 96748 94912 96788
rect 109664 96748 109704 96788
rect 109746 96748 109786 96788
rect 109828 96748 109868 96788
rect 109910 96748 109950 96788
rect 109992 96748 110032 96788
rect 124784 96748 124824 96788
rect 124866 96748 124906 96788
rect 124948 96748 124988 96788
rect 125030 96748 125070 96788
rect 125112 96748 125152 96788
rect 139904 96748 139944 96788
rect 139986 96748 140026 96788
rect 140068 96748 140108 96788
rect 140150 96748 140190 96788
rect 140232 96748 140272 96788
rect 78184 95992 78224 96032
rect 78266 95992 78306 96032
rect 78348 95992 78388 96032
rect 78430 95992 78470 96032
rect 78512 95992 78552 96032
rect 93304 95992 93344 96032
rect 93386 95992 93426 96032
rect 93468 95992 93508 96032
rect 93550 95992 93590 96032
rect 93632 95992 93672 96032
rect 108424 95992 108464 96032
rect 108506 95992 108546 96032
rect 108588 95992 108628 96032
rect 108670 95992 108710 96032
rect 108752 95992 108792 96032
rect 123544 95992 123584 96032
rect 123626 95992 123666 96032
rect 123708 95992 123748 96032
rect 123790 95992 123830 96032
rect 123872 95992 123912 96032
rect 138664 95992 138704 96032
rect 138746 95992 138786 96032
rect 138828 95992 138868 96032
rect 138910 95992 138950 96032
rect 138992 95992 139032 96032
rect 79424 95236 79464 95276
rect 79506 95236 79546 95276
rect 79588 95236 79628 95276
rect 79670 95236 79710 95276
rect 79752 95236 79792 95276
rect 94544 95236 94584 95276
rect 94626 95236 94666 95276
rect 94708 95236 94748 95276
rect 94790 95236 94830 95276
rect 94872 95236 94912 95276
rect 109664 95236 109704 95276
rect 109746 95236 109786 95276
rect 109828 95236 109868 95276
rect 109910 95236 109950 95276
rect 109992 95236 110032 95276
rect 124784 95236 124824 95276
rect 124866 95236 124906 95276
rect 124948 95236 124988 95276
rect 125030 95236 125070 95276
rect 125112 95236 125152 95276
rect 139904 95236 139944 95276
rect 139986 95236 140026 95276
rect 140068 95236 140108 95276
rect 140150 95236 140190 95276
rect 140232 95236 140272 95276
rect 78184 94480 78224 94520
rect 78266 94480 78306 94520
rect 78348 94480 78388 94520
rect 78430 94480 78470 94520
rect 78512 94480 78552 94520
rect 93304 94480 93344 94520
rect 93386 94480 93426 94520
rect 93468 94480 93508 94520
rect 93550 94480 93590 94520
rect 93632 94480 93672 94520
rect 108424 94480 108464 94520
rect 108506 94480 108546 94520
rect 108588 94480 108628 94520
rect 108670 94480 108710 94520
rect 108752 94480 108792 94520
rect 123544 94480 123584 94520
rect 123626 94480 123666 94520
rect 123708 94480 123748 94520
rect 123790 94480 123830 94520
rect 123872 94480 123912 94520
rect 138664 94480 138704 94520
rect 138746 94480 138786 94520
rect 138828 94480 138868 94520
rect 138910 94480 138950 94520
rect 138992 94480 139032 94520
rect 79424 93724 79464 93764
rect 79506 93724 79546 93764
rect 79588 93724 79628 93764
rect 79670 93724 79710 93764
rect 79752 93724 79792 93764
rect 94544 93724 94584 93764
rect 94626 93724 94666 93764
rect 94708 93724 94748 93764
rect 94790 93724 94830 93764
rect 94872 93724 94912 93764
rect 109664 93724 109704 93764
rect 109746 93724 109786 93764
rect 109828 93724 109868 93764
rect 109910 93724 109950 93764
rect 109992 93724 110032 93764
rect 124784 93724 124824 93764
rect 124866 93724 124906 93764
rect 124948 93724 124988 93764
rect 125030 93724 125070 93764
rect 125112 93724 125152 93764
rect 139904 93724 139944 93764
rect 139986 93724 140026 93764
rect 140068 93724 140108 93764
rect 140150 93724 140190 93764
rect 140232 93724 140272 93764
rect 78184 92968 78224 93008
rect 78266 92968 78306 93008
rect 78348 92968 78388 93008
rect 78430 92968 78470 93008
rect 78512 92968 78552 93008
rect 93304 92968 93344 93008
rect 93386 92968 93426 93008
rect 93468 92968 93508 93008
rect 93550 92968 93590 93008
rect 93632 92968 93672 93008
rect 108424 92968 108464 93008
rect 108506 92968 108546 93008
rect 108588 92968 108628 93008
rect 108670 92968 108710 93008
rect 108752 92968 108792 93008
rect 123544 92968 123584 93008
rect 123626 92968 123666 93008
rect 123708 92968 123748 93008
rect 123790 92968 123830 93008
rect 123872 92968 123912 93008
rect 138664 92968 138704 93008
rect 138746 92968 138786 93008
rect 138828 92968 138868 93008
rect 138910 92968 138950 93008
rect 138992 92968 139032 93008
rect 79424 92212 79464 92252
rect 79506 92212 79546 92252
rect 79588 92212 79628 92252
rect 79670 92212 79710 92252
rect 79752 92212 79792 92252
rect 94544 92212 94584 92252
rect 94626 92212 94666 92252
rect 94708 92212 94748 92252
rect 94790 92212 94830 92252
rect 94872 92212 94912 92252
rect 109664 92212 109704 92252
rect 109746 92212 109786 92252
rect 109828 92212 109868 92252
rect 109910 92212 109950 92252
rect 109992 92212 110032 92252
rect 124784 92212 124824 92252
rect 124866 92212 124906 92252
rect 124948 92212 124988 92252
rect 125030 92212 125070 92252
rect 125112 92212 125152 92252
rect 139904 92212 139944 92252
rect 139986 92212 140026 92252
rect 140068 92212 140108 92252
rect 140150 92212 140190 92252
rect 140232 92212 140272 92252
rect 78184 91456 78224 91496
rect 78266 91456 78306 91496
rect 78348 91456 78388 91496
rect 78430 91456 78470 91496
rect 78512 91456 78552 91496
rect 93304 91456 93344 91496
rect 93386 91456 93426 91496
rect 93468 91456 93508 91496
rect 93550 91456 93590 91496
rect 93632 91456 93672 91496
rect 108424 91456 108464 91496
rect 108506 91456 108546 91496
rect 108588 91456 108628 91496
rect 108670 91456 108710 91496
rect 108752 91456 108792 91496
rect 123544 91456 123584 91496
rect 123626 91456 123666 91496
rect 123708 91456 123748 91496
rect 123790 91456 123830 91496
rect 123872 91456 123912 91496
rect 138664 91456 138704 91496
rect 138746 91456 138786 91496
rect 138828 91456 138868 91496
rect 138910 91456 138950 91496
rect 138992 91456 139032 91496
rect 79424 90700 79464 90740
rect 79506 90700 79546 90740
rect 79588 90700 79628 90740
rect 79670 90700 79710 90740
rect 79752 90700 79792 90740
rect 94544 90700 94584 90740
rect 94626 90700 94666 90740
rect 94708 90700 94748 90740
rect 94790 90700 94830 90740
rect 94872 90700 94912 90740
rect 109664 90700 109704 90740
rect 109746 90700 109786 90740
rect 109828 90700 109868 90740
rect 109910 90700 109950 90740
rect 109992 90700 110032 90740
rect 124784 90700 124824 90740
rect 124866 90700 124906 90740
rect 124948 90700 124988 90740
rect 125030 90700 125070 90740
rect 125112 90700 125152 90740
rect 139904 90700 139944 90740
rect 139986 90700 140026 90740
rect 140068 90700 140108 90740
rect 140150 90700 140190 90740
rect 140232 90700 140272 90740
rect 78184 89944 78224 89984
rect 78266 89944 78306 89984
rect 78348 89944 78388 89984
rect 78430 89944 78470 89984
rect 78512 89944 78552 89984
rect 93304 89944 93344 89984
rect 93386 89944 93426 89984
rect 93468 89944 93508 89984
rect 93550 89944 93590 89984
rect 93632 89944 93672 89984
rect 108424 89944 108464 89984
rect 108506 89944 108546 89984
rect 108588 89944 108628 89984
rect 108670 89944 108710 89984
rect 108752 89944 108792 89984
rect 123544 89944 123584 89984
rect 123626 89944 123666 89984
rect 123708 89944 123748 89984
rect 123790 89944 123830 89984
rect 123872 89944 123912 89984
rect 138664 89944 138704 89984
rect 138746 89944 138786 89984
rect 138828 89944 138868 89984
rect 138910 89944 138950 89984
rect 138992 89944 139032 89984
rect 79424 89188 79464 89228
rect 79506 89188 79546 89228
rect 79588 89188 79628 89228
rect 79670 89188 79710 89228
rect 79752 89188 79792 89228
rect 94544 89188 94584 89228
rect 94626 89188 94666 89228
rect 94708 89188 94748 89228
rect 94790 89188 94830 89228
rect 94872 89188 94912 89228
rect 109664 89188 109704 89228
rect 109746 89188 109786 89228
rect 109828 89188 109868 89228
rect 109910 89188 109950 89228
rect 109992 89188 110032 89228
rect 124784 89188 124824 89228
rect 124866 89188 124906 89228
rect 124948 89188 124988 89228
rect 125030 89188 125070 89228
rect 125112 89188 125152 89228
rect 139904 89188 139944 89228
rect 139986 89188 140026 89228
rect 140068 89188 140108 89228
rect 140150 89188 140190 89228
rect 140232 89188 140272 89228
rect 90700 89104 90740 89144
rect 92140 89104 92180 89144
rect 78184 88432 78224 88472
rect 78266 88432 78306 88472
rect 78348 88432 78388 88472
rect 78430 88432 78470 88472
rect 78512 88432 78552 88472
rect 93304 88432 93344 88472
rect 93386 88432 93426 88472
rect 93468 88432 93508 88472
rect 93550 88432 93590 88472
rect 93632 88432 93672 88472
rect 108424 88432 108464 88472
rect 108506 88432 108546 88472
rect 108588 88432 108628 88472
rect 108670 88432 108710 88472
rect 108752 88432 108792 88472
rect 123544 88432 123584 88472
rect 123626 88432 123666 88472
rect 123708 88432 123748 88472
rect 123790 88432 123830 88472
rect 123872 88432 123912 88472
rect 138664 88432 138704 88472
rect 138746 88432 138786 88472
rect 138828 88432 138868 88472
rect 138910 88432 138950 88472
rect 138992 88432 139032 88472
rect 79424 87676 79464 87716
rect 79506 87676 79546 87716
rect 79588 87676 79628 87716
rect 79670 87676 79710 87716
rect 79752 87676 79792 87716
rect 94544 87676 94584 87716
rect 94626 87676 94666 87716
rect 94708 87676 94748 87716
rect 94790 87676 94830 87716
rect 94872 87676 94912 87716
rect 109664 87676 109704 87716
rect 109746 87676 109786 87716
rect 109828 87676 109868 87716
rect 109910 87676 109950 87716
rect 109992 87676 110032 87716
rect 124784 87676 124824 87716
rect 124866 87676 124906 87716
rect 124948 87676 124988 87716
rect 125030 87676 125070 87716
rect 125112 87676 125152 87716
rect 139904 87676 139944 87716
rect 139986 87676 140026 87716
rect 140068 87676 140108 87716
rect 140150 87676 140190 87716
rect 140232 87676 140272 87716
rect 78184 86920 78224 86960
rect 78266 86920 78306 86960
rect 78348 86920 78388 86960
rect 78430 86920 78470 86960
rect 78512 86920 78552 86960
rect 93304 86920 93344 86960
rect 93386 86920 93426 86960
rect 93468 86920 93508 86960
rect 93550 86920 93590 86960
rect 93632 86920 93672 86960
rect 108424 86920 108464 86960
rect 108506 86920 108546 86960
rect 108588 86920 108628 86960
rect 108670 86920 108710 86960
rect 108752 86920 108792 86960
rect 123544 86920 123584 86960
rect 123626 86920 123666 86960
rect 123708 86920 123748 86960
rect 123790 86920 123830 86960
rect 123872 86920 123912 86960
rect 138664 86920 138704 86960
rect 138746 86920 138786 86960
rect 138828 86920 138868 86960
rect 138910 86920 138950 86960
rect 138992 86920 139032 86960
rect 79424 86164 79464 86204
rect 79506 86164 79546 86204
rect 79588 86164 79628 86204
rect 79670 86164 79710 86204
rect 79752 86164 79792 86204
rect 94544 86164 94584 86204
rect 94626 86164 94666 86204
rect 94708 86164 94748 86204
rect 94790 86164 94830 86204
rect 94872 86164 94912 86204
rect 109664 86164 109704 86204
rect 109746 86164 109786 86204
rect 109828 86164 109868 86204
rect 109910 86164 109950 86204
rect 109992 86164 110032 86204
rect 124784 86164 124824 86204
rect 124866 86164 124906 86204
rect 124948 86164 124988 86204
rect 125030 86164 125070 86204
rect 125112 86164 125152 86204
rect 139904 86164 139944 86204
rect 139986 86164 140026 86204
rect 140068 86164 140108 86204
rect 140150 86164 140190 86204
rect 140232 86164 140272 86204
rect 78184 85408 78224 85448
rect 78266 85408 78306 85448
rect 78348 85408 78388 85448
rect 78430 85408 78470 85448
rect 78512 85408 78552 85448
rect 93304 85408 93344 85448
rect 93386 85408 93426 85448
rect 93468 85408 93508 85448
rect 93550 85408 93590 85448
rect 93632 85408 93672 85448
rect 108424 85408 108464 85448
rect 108506 85408 108546 85448
rect 108588 85408 108628 85448
rect 108670 85408 108710 85448
rect 108752 85408 108792 85448
rect 123544 85408 123584 85448
rect 123626 85408 123666 85448
rect 123708 85408 123748 85448
rect 123790 85408 123830 85448
rect 123872 85408 123912 85448
rect 138664 85408 138704 85448
rect 138746 85408 138786 85448
rect 138828 85408 138868 85448
rect 138910 85408 138950 85448
rect 138992 85408 139032 85448
rect 79424 84652 79464 84692
rect 79506 84652 79546 84692
rect 79588 84652 79628 84692
rect 79670 84652 79710 84692
rect 79752 84652 79792 84692
rect 94544 84652 94584 84692
rect 94626 84652 94666 84692
rect 94708 84652 94748 84692
rect 94790 84652 94830 84692
rect 94872 84652 94912 84692
rect 109664 84652 109704 84692
rect 109746 84652 109786 84692
rect 109828 84652 109868 84692
rect 109910 84652 109950 84692
rect 109992 84652 110032 84692
rect 124784 84652 124824 84692
rect 124866 84652 124906 84692
rect 124948 84652 124988 84692
rect 125030 84652 125070 84692
rect 125112 84652 125152 84692
rect 139904 84652 139944 84692
rect 139986 84652 140026 84692
rect 140068 84652 140108 84692
rect 140150 84652 140190 84692
rect 140232 84652 140272 84692
rect 78184 83896 78224 83936
rect 78266 83896 78306 83936
rect 78348 83896 78388 83936
rect 78430 83896 78470 83936
rect 78512 83896 78552 83936
rect 93304 83896 93344 83936
rect 93386 83896 93426 83936
rect 93468 83896 93508 83936
rect 93550 83896 93590 83936
rect 93632 83896 93672 83936
rect 108424 83896 108464 83936
rect 108506 83896 108546 83936
rect 108588 83896 108628 83936
rect 108670 83896 108710 83936
rect 108752 83896 108792 83936
rect 123544 83896 123584 83936
rect 123626 83896 123666 83936
rect 123708 83896 123748 83936
rect 123790 83896 123830 83936
rect 123872 83896 123912 83936
rect 138664 83896 138704 83936
rect 138746 83896 138786 83936
rect 138828 83896 138868 83936
rect 138910 83896 138950 83936
rect 138992 83896 139032 83936
rect 79424 83140 79464 83180
rect 79506 83140 79546 83180
rect 79588 83140 79628 83180
rect 79670 83140 79710 83180
rect 79752 83140 79792 83180
rect 94544 83140 94584 83180
rect 94626 83140 94666 83180
rect 94708 83140 94748 83180
rect 94790 83140 94830 83180
rect 94872 83140 94912 83180
rect 109664 83140 109704 83180
rect 109746 83140 109786 83180
rect 109828 83140 109868 83180
rect 109910 83140 109950 83180
rect 109992 83140 110032 83180
rect 124784 83140 124824 83180
rect 124866 83140 124906 83180
rect 124948 83140 124988 83180
rect 125030 83140 125070 83180
rect 125112 83140 125152 83180
rect 139904 83140 139944 83180
rect 139986 83140 140026 83180
rect 140068 83140 140108 83180
rect 140150 83140 140190 83180
rect 140232 83140 140272 83180
rect 78184 82384 78224 82424
rect 78266 82384 78306 82424
rect 78348 82384 78388 82424
rect 78430 82384 78470 82424
rect 78512 82384 78552 82424
rect 93304 82384 93344 82424
rect 93386 82384 93426 82424
rect 93468 82384 93508 82424
rect 93550 82384 93590 82424
rect 93632 82384 93672 82424
rect 108424 82384 108464 82424
rect 108506 82384 108546 82424
rect 108588 82384 108628 82424
rect 108670 82384 108710 82424
rect 108752 82384 108792 82424
rect 123544 82384 123584 82424
rect 123626 82384 123666 82424
rect 123708 82384 123748 82424
rect 123790 82384 123830 82424
rect 123872 82384 123912 82424
rect 138664 82384 138704 82424
rect 138746 82384 138786 82424
rect 138828 82384 138868 82424
rect 138910 82384 138950 82424
rect 138992 82384 139032 82424
rect 79424 81628 79464 81668
rect 79506 81628 79546 81668
rect 79588 81628 79628 81668
rect 79670 81628 79710 81668
rect 79752 81628 79792 81668
rect 94544 81628 94584 81668
rect 94626 81628 94666 81668
rect 94708 81628 94748 81668
rect 94790 81628 94830 81668
rect 94872 81628 94912 81668
rect 109664 81628 109704 81668
rect 109746 81628 109786 81668
rect 109828 81628 109868 81668
rect 109910 81628 109950 81668
rect 109992 81628 110032 81668
rect 124784 81628 124824 81668
rect 124866 81628 124906 81668
rect 124948 81628 124988 81668
rect 125030 81628 125070 81668
rect 125112 81628 125152 81668
rect 139904 81628 139944 81668
rect 139986 81628 140026 81668
rect 140068 81628 140108 81668
rect 140150 81628 140190 81668
rect 140232 81628 140272 81668
rect 78184 80872 78224 80912
rect 78266 80872 78306 80912
rect 78348 80872 78388 80912
rect 78430 80872 78470 80912
rect 78512 80872 78552 80912
rect 93304 80872 93344 80912
rect 93386 80872 93426 80912
rect 93468 80872 93508 80912
rect 93550 80872 93590 80912
rect 93632 80872 93672 80912
rect 108424 80872 108464 80912
rect 108506 80872 108546 80912
rect 108588 80872 108628 80912
rect 108670 80872 108710 80912
rect 108752 80872 108792 80912
rect 123544 80872 123584 80912
rect 123626 80872 123666 80912
rect 123708 80872 123748 80912
rect 123790 80872 123830 80912
rect 123872 80872 123912 80912
rect 138664 80872 138704 80912
rect 138746 80872 138786 80912
rect 138828 80872 138868 80912
rect 138910 80872 138950 80912
rect 138992 80872 139032 80912
rect 79424 80116 79464 80156
rect 79506 80116 79546 80156
rect 79588 80116 79628 80156
rect 79670 80116 79710 80156
rect 79752 80116 79792 80156
rect 94544 80116 94584 80156
rect 94626 80116 94666 80156
rect 94708 80116 94748 80156
rect 94790 80116 94830 80156
rect 94872 80116 94912 80156
rect 109664 80116 109704 80156
rect 109746 80116 109786 80156
rect 109828 80116 109868 80156
rect 109910 80116 109950 80156
rect 109992 80116 110032 80156
rect 124784 80116 124824 80156
rect 124866 80116 124906 80156
rect 124948 80116 124988 80156
rect 125030 80116 125070 80156
rect 125112 80116 125152 80156
rect 139904 80116 139944 80156
rect 139986 80116 140026 80156
rect 140068 80116 140108 80156
rect 140150 80116 140190 80156
rect 140232 80116 140272 80156
rect 78184 79360 78224 79400
rect 78266 79360 78306 79400
rect 78348 79360 78388 79400
rect 78430 79360 78470 79400
rect 78512 79360 78552 79400
rect 93304 79360 93344 79400
rect 93386 79360 93426 79400
rect 93468 79360 93508 79400
rect 93550 79360 93590 79400
rect 93632 79360 93672 79400
rect 108424 79360 108464 79400
rect 108506 79360 108546 79400
rect 108588 79360 108628 79400
rect 108670 79360 108710 79400
rect 108752 79360 108792 79400
rect 123544 79360 123584 79400
rect 123626 79360 123666 79400
rect 123708 79360 123748 79400
rect 123790 79360 123830 79400
rect 123872 79360 123912 79400
rect 138664 79360 138704 79400
rect 138746 79360 138786 79400
rect 138828 79360 138868 79400
rect 138910 79360 138950 79400
rect 138992 79360 139032 79400
rect 79424 78604 79464 78644
rect 79506 78604 79546 78644
rect 79588 78604 79628 78644
rect 79670 78604 79710 78644
rect 79752 78604 79792 78644
rect 94544 78604 94584 78644
rect 94626 78604 94666 78644
rect 94708 78604 94748 78644
rect 94790 78604 94830 78644
rect 94872 78604 94912 78644
rect 109664 78604 109704 78644
rect 109746 78604 109786 78644
rect 109828 78604 109868 78644
rect 109910 78604 109950 78644
rect 109992 78604 110032 78644
rect 124784 78604 124824 78644
rect 124866 78604 124906 78644
rect 124948 78604 124988 78644
rect 125030 78604 125070 78644
rect 125112 78604 125152 78644
rect 139904 78604 139944 78644
rect 139986 78604 140026 78644
rect 140068 78604 140108 78644
rect 140150 78604 140190 78644
rect 140232 78604 140272 78644
rect 78184 77848 78224 77888
rect 78266 77848 78306 77888
rect 78348 77848 78388 77888
rect 78430 77848 78470 77888
rect 78512 77848 78552 77888
rect 93304 77848 93344 77888
rect 93386 77848 93426 77888
rect 93468 77848 93508 77888
rect 93550 77848 93590 77888
rect 93632 77848 93672 77888
rect 108424 77848 108464 77888
rect 108506 77848 108546 77888
rect 108588 77848 108628 77888
rect 108670 77848 108710 77888
rect 108752 77848 108792 77888
rect 123544 77848 123584 77888
rect 123626 77848 123666 77888
rect 123708 77848 123748 77888
rect 123790 77848 123830 77888
rect 123872 77848 123912 77888
rect 138664 77848 138704 77888
rect 138746 77848 138786 77888
rect 138828 77848 138868 77888
rect 138910 77848 138950 77888
rect 138992 77848 139032 77888
rect 79424 77092 79464 77132
rect 79506 77092 79546 77132
rect 79588 77092 79628 77132
rect 79670 77092 79710 77132
rect 79752 77092 79792 77132
rect 94544 77092 94584 77132
rect 94626 77092 94666 77132
rect 94708 77092 94748 77132
rect 94790 77092 94830 77132
rect 94872 77092 94912 77132
rect 109664 77092 109704 77132
rect 109746 77092 109786 77132
rect 109828 77092 109868 77132
rect 109910 77092 109950 77132
rect 109992 77092 110032 77132
rect 124784 77092 124824 77132
rect 124866 77092 124906 77132
rect 124948 77092 124988 77132
rect 125030 77092 125070 77132
rect 125112 77092 125152 77132
rect 139904 77092 139944 77132
rect 139986 77092 140026 77132
rect 140068 77092 140108 77132
rect 140150 77092 140190 77132
rect 140232 77092 140272 77132
rect 78184 76336 78224 76376
rect 78266 76336 78306 76376
rect 78348 76336 78388 76376
rect 78430 76336 78470 76376
rect 78512 76336 78552 76376
rect 93304 76336 93344 76376
rect 93386 76336 93426 76376
rect 93468 76336 93508 76376
rect 93550 76336 93590 76376
rect 93632 76336 93672 76376
rect 108424 76336 108464 76376
rect 108506 76336 108546 76376
rect 108588 76336 108628 76376
rect 108670 76336 108710 76376
rect 108752 76336 108792 76376
rect 123544 76336 123584 76376
rect 123626 76336 123666 76376
rect 123708 76336 123748 76376
rect 123790 76336 123830 76376
rect 123872 76336 123912 76376
rect 138664 76336 138704 76376
rect 138746 76336 138786 76376
rect 138828 76336 138868 76376
rect 138910 76336 138950 76376
rect 138992 76336 139032 76376
rect 79424 75580 79464 75620
rect 79506 75580 79546 75620
rect 79588 75580 79628 75620
rect 79670 75580 79710 75620
rect 79752 75580 79792 75620
rect 94544 75580 94584 75620
rect 94626 75580 94666 75620
rect 94708 75580 94748 75620
rect 94790 75580 94830 75620
rect 94872 75580 94912 75620
rect 109664 75580 109704 75620
rect 109746 75580 109786 75620
rect 109828 75580 109868 75620
rect 109910 75580 109950 75620
rect 109992 75580 110032 75620
rect 124784 75580 124824 75620
rect 124866 75580 124906 75620
rect 124948 75580 124988 75620
rect 125030 75580 125070 75620
rect 125112 75580 125152 75620
rect 139904 75580 139944 75620
rect 139986 75580 140026 75620
rect 140068 75580 140108 75620
rect 140150 75580 140190 75620
rect 140232 75580 140272 75620
rect 90700 71212 90740 71252
rect 92140 71212 92180 71252
<< metal4 >>
rect 79424 148196 79792 148205
rect 79464 148156 79506 148196
rect 79546 148156 79588 148196
rect 79628 148156 79670 148196
rect 79710 148156 79752 148196
rect 79424 148147 79792 148156
rect 94544 148196 94912 148205
rect 94584 148156 94626 148196
rect 94666 148156 94708 148196
rect 94748 148156 94790 148196
rect 94830 148156 94872 148196
rect 94544 148147 94912 148156
rect 109664 148196 110032 148205
rect 109704 148156 109746 148196
rect 109786 148156 109828 148196
rect 109868 148156 109910 148196
rect 109950 148156 109992 148196
rect 109664 148147 110032 148156
rect 124784 148196 125152 148205
rect 124824 148156 124866 148196
rect 124906 148156 124948 148196
rect 124988 148156 125030 148196
rect 125070 148156 125112 148196
rect 124784 148147 125152 148156
rect 139904 148196 140272 148205
rect 139944 148156 139986 148196
rect 140026 148156 140068 148196
rect 140108 148156 140150 148196
rect 140190 148156 140232 148196
rect 139904 148147 140272 148156
rect 78184 147440 78552 147449
rect 78224 147400 78266 147440
rect 78306 147400 78348 147440
rect 78388 147400 78430 147440
rect 78470 147400 78512 147440
rect 78184 147391 78552 147400
rect 93304 147440 93672 147449
rect 93344 147400 93386 147440
rect 93426 147400 93468 147440
rect 93508 147400 93550 147440
rect 93590 147400 93632 147440
rect 93304 147391 93672 147400
rect 108424 147440 108792 147449
rect 108464 147400 108506 147440
rect 108546 147400 108588 147440
rect 108628 147400 108670 147440
rect 108710 147400 108752 147440
rect 108424 147391 108792 147400
rect 123544 147440 123912 147449
rect 123584 147400 123626 147440
rect 123666 147400 123708 147440
rect 123748 147400 123790 147440
rect 123830 147400 123872 147440
rect 123544 147391 123912 147400
rect 138664 147440 139032 147449
rect 138704 147400 138746 147440
rect 138786 147400 138828 147440
rect 138868 147400 138910 147440
rect 138950 147400 138992 147440
rect 138664 147391 139032 147400
rect 79424 146684 79792 146693
rect 79464 146644 79506 146684
rect 79546 146644 79588 146684
rect 79628 146644 79670 146684
rect 79710 146644 79752 146684
rect 79424 146635 79792 146644
rect 94544 146684 94912 146693
rect 94584 146644 94626 146684
rect 94666 146644 94708 146684
rect 94748 146644 94790 146684
rect 94830 146644 94872 146684
rect 94544 146635 94912 146644
rect 109664 146684 110032 146693
rect 109704 146644 109746 146684
rect 109786 146644 109828 146684
rect 109868 146644 109910 146684
rect 109950 146644 109992 146684
rect 109664 146635 110032 146644
rect 124784 146684 125152 146693
rect 124824 146644 124866 146684
rect 124906 146644 124948 146684
rect 124988 146644 125030 146684
rect 125070 146644 125112 146684
rect 124784 146635 125152 146644
rect 139904 146684 140272 146693
rect 139944 146644 139986 146684
rect 140026 146644 140068 146684
rect 140108 146644 140150 146684
rect 140190 146644 140232 146684
rect 139904 146635 140272 146644
rect 78184 145928 78552 145937
rect 78224 145888 78266 145928
rect 78306 145888 78348 145928
rect 78388 145888 78430 145928
rect 78470 145888 78512 145928
rect 78184 145879 78552 145888
rect 93304 145928 93672 145937
rect 93344 145888 93386 145928
rect 93426 145888 93468 145928
rect 93508 145888 93550 145928
rect 93590 145888 93632 145928
rect 93304 145879 93672 145888
rect 108424 145928 108792 145937
rect 108464 145888 108506 145928
rect 108546 145888 108588 145928
rect 108628 145888 108670 145928
rect 108710 145888 108752 145928
rect 108424 145879 108792 145888
rect 123544 145928 123912 145937
rect 123584 145888 123626 145928
rect 123666 145888 123708 145928
rect 123748 145888 123790 145928
rect 123830 145888 123872 145928
rect 123544 145879 123912 145888
rect 138664 145928 139032 145937
rect 138704 145888 138746 145928
rect 138786 145888 138828 145928
rect 138868 145888 138910 145928
rect 138950 145888 138992 145928
rect 138664 145879 139032 145888
rect 79424 145172 79792 145181
rect 79464 145132 79506 145172
rect 79546 145132 79588 145172
rect 79628 145132 79670 145172
rect 79710 145132 79752 145172
rect 79424 145123 79792 145132
rect 94544 145172 94912 145181
rect 94584 145132 94626 145172
rect 94666 145132 94708 145172
rect 94748 145132 94790 145172
rect 94830 145132 94872 145172
rect 94544 145123 94912 145132
rect 109664 145172 110032 145181
rect 109704 145132 109746 145172
rect 109786 145132 109828 145172
rect 109868 145132 109910 145172
rect 109950 145132 109992 145172
rect 109664 145123 110032 145132
rect 124784 145172 125152 145181
rect 124824 145132 124866 145172
rect 124906 145132 124948 145172
rect 124988 145132 125030 145172
rect 125070 145132 125112 145172
rect 124784 145123 125152 145132
rect 139904 145172 140272 145181
rect 139944 145132 139986 145172
rect 140026 145132 140068 145172
rect 140108 145132 140150 145172
rect 140190 145132 140232 145172
rect 139904 145123 140272 145132
rect 78184 144416 78552 144425
rect 78224 144376 78266 144416
rect 78306 144376 78348 144416
rect 78388 144376 78430 144416
rect 78470 144376 78512 144416
rect 78184 144367 78552 144376
rect 93304 144416 93672 144425
rect 93344 144376 93386 144416
rect 93426 144376 93468 144416
rect 93508 144376 93550 144416
rect 93590 144376 93632 144416
rect 93304 144367 93672 144376
rect 108424 144416 108792 144425
rect 108464 144376 108506 144416
rect 108546 144376 108588 144416
rect 108628 144376 108670 144416
rect 108710 144376 108752 144416
rect 108424 144367 108792 144376
rect 123544 144416 123912 144425
rect 123584 144376 123626 144416
rect 123666 144376 123708 144416
rect 123748 144376 123790 144416
rect 123830 144376 123872 144416
rect 123544 144367 123912 144376
rect 138664 144416 139032 144425
rect 138704 144376 138746 144416
rect 138786 144376 138828 144416
rect 138868 144376 138910 144416
rect 138950 144376 138992 144416
rect 138664 144367 139032 144376
rect 79424 143660 79792 143669
rect 79464 143620 79506 143660
rect 79546 143620 79588 143660
rect 79628 143620 79670 143660
rect 79710 143620 79752 143660
rect 79424 143611 79792 143620
rect 94544 143660 94912 143669
rect 94584 143620 94626 143660
rect 94666 143620 94708 143660
rect 94748 143620 94790 143660
rect 94830 143620 94872 143660
rect 94544 143611 94912 143620
rect 109664 143660 110032 143669
rect 109704 143620 109746 143660
rect 109786 143620 109828 143660
rect 109868 143620 109910 143660
rect 109950 143620 109992 143660
rect 109664 143611 110032 143620
rect 124784 143660 125152 143669
rect 124824 143620 124866 143660
rect 124906 143620 124948 143660
rect 124988 143620 125030 143660
rect 125070 143620 125112 143660
rect 124784 143611 125152 143620
rect 139904 143660 140272 143669
rect 139944 143620 139986 143660
rect 140026 143620 140068 143660
rect 140108 143620 140150 143660
rect 140190 143620 140232 143660
rect 139904 143611 140272 143620
rect 78184 142904 78552 142913
rect 78224 142864 78266 142904
rect 78306 142864 78348 142904
rect 78388 142864 78430 142904
rect 78470 142864 78512 142904
rect 78184 142855 78552 142864
rect 93304 142904 93672 142913
rect 93344 142864 93386 142904
rect 93426 142864 93468 142904
rect 93508 142864 93550 142904
rect 93590 142864 93632 142904
rect 93304 142855 93672 142864
rect 108424 142904 108792 142913
rect 108464 142864 108506 142904
rect 108546 142864 108588 142904
rect 108628 142864 108670 142904
rect 108710 142864 108752 142904
rect 108424 142855 108792 142864
rect 123544 142904 123912 142913
rect 123584 142864 123626 142904
rect 123666 142864 123708 142904
rect 123748 142864 123790 142904
rect 123830 142864 123872 142904
rect 123544 142855 123912 142864
rect 138664 142904 139032 142913
rect 138704 142864 138746 142904
rect 138786 142864 138828 142904
rect 138868 142864 138910 142904
rect 138950 142864 138992 142904
rect 138664 142855 139032 142864
rect 79424 142148 79792 142157
rect 79464 142108 79506 142148
rect 79546 142108 79588 142148
rect 79628 142108 79670 142148
rect 79710 142108 79752 142148
rect 79424 142099 79792 142108
rect 94544 142148 94912 142157
rect 94584 142108 94626 142148
rect 94666 142108 94708 142148
rect 94748 142108 94790 142148
rect 94830 142108 94872 142148
rect 94544 142099 94912 142108
rect 109664 142148 110032 142157
rect 109704 142108 109746 142148
rect 109786 142108 109828 142148
rect 109868 142108 109910 142148
rect 109950 142108 109992 142148
rect 109664 142099 110032 142108
rect 124784 142148 125152 142157
rect 124824 142108 124866 142148
rect 124906 142108 124948 142148
rect 124988 142108 125030 142148
rect 125070 142108 125112 142148
rect 124784 142099 125152 142108
rect 139904 142148 140272 142157
rect 139944 142108 139986 142148
rect 140026 142108 140068 142148
rect 140108 142108 140150 142148
rect 140190 142108 140232 142148
rect 139904 142099 140272 142108
rect 78184 141392 78552 141401
rect 78224 141352 78266 141392
rect 78306 141352 78348 141392
rect 78388 141352 78430 141392
rect 78470 141352 78512 141392
rect 78184 141343 78552 141352
rect 93304 141392 93672 141401
rect 93344 141352 93386 141392
rect 93426 141352 93468 141392
rect 93508 141352 93550 141392
rect 93590 141352 93632 141392
rect 93304 141343 93672 141352
rect 108424 141392 108792 141401
rect 108464 141352 108506 141392
rect 108546 141352 108588 141392
rect 108628 141352 108670 141392
rect 108710 141352 108752 141392
rect 108424 141343 108792 141352
rect 123544 141392 123912 141401
rect 123584 141352 123626 141392
rect 123666 141352 123708 141392
rect 123748 141352 123790 141392
rect 123830 141352 123872 141392
rect 123544 141343 123912 141352
rect 138664 141392 139032 141401
rect 138704 141352 138746 141392
rect 138786 141352 138828 141392
rect 138868 141352 138910 141392
rect 138950 141352 138992 141392
rect 138664 141343 139032 141352
rect 79424 140636 79792 140645
rect 79464 140596 79506 140636
rect 79546 140596 79588 140636
rect 79628 140596 79670 140636
rect 79710 140596 79752 140636
rect 79424 140587 79792 140596
rect 94544 140636 94912 140645
rect 94584 140596 94626 140636
rect 94666 140596 94708 140636
rect 94748 140596 94790 140636
rect 94830 140596 94872 140636
rect 94544 140587 94912 140596
rect 109664 140636 110032 140645
rect 109704 140596 109746 140636
rect 109786 140596 109828 140636
rect 109868 140596 109910 140636
rect 109950 140596 109992 140636
rect 109664 140587 110032 140596
rect 124784 140636 125152 140645
rect 124824 140596 124866 140636
rect 124906 140596 124948 140636
rect 124988 140596 125030 140636
rect 125070 140596 125112 140636
rect 124784 140587 125152 140596
rect 139904 140636 140272 140645
rect 139944 140596 139986 140636
rect 140026 140596 140068 140636
rect 140108 140596 140150 140636
rect 140190 140596 140232 140636
rect 139904 140587 140272 140596
rect 78184 139880 78552 139889
rect 78224 139840 78266 139880
rect 78306 139840 78348 139880
rect 78388 139840 78430 139880
rect 78470 139840 78512 139880
rect 78184 139831 78552 139840
rect 93304 139880 93672 139889
rect 93344 139840 93386 139880
rect 93426 139840 93468 139880
rect 93508 139840 93550 139880
rect 93590 139840 93632 139880
rect 93304 139831 93672 139840
rect 108424 139880 108792 139889
rect 108464 139840 108506 139880
rect 108546 139840 108588 139880
rect 108628 139840 108670 139880
rect 108710 139840 108752 139880
rect 108424 139831 108792 139840
rect 123544 139880 123912 139889
rect 123584 139840 123626 139880
rect 123666 139840 123708 139880
rect 123748 139840 123790 139880
rect 123830 139840 123872 139880
rect 123544 139831 123912 139840
rect 138664 139880 139032 139889
rect 138704 139840 138746 139880
rect 138786 139840 138828 139880
rect 138868 139840 138910 139880
rect 138950 139840 138992 139880
rect 138664 139831 139032 139840
rect 79424 139124 79792 139133
rect 79464 139084 79506 139124
rect 79546 139084 79588 139124
rect 79628 139084 79670 139124
rect 79710 139084 79752 139124
rect 79424 139075 79792 139084
rect 94544 139124 94912 139133
rect 94584 139084 94626 139124
rect 94666 139084 94708 139124
rect 94748 139084 94790 139124
rect 94830 139084 94872 139124
rect 94544 139075 94912 139084
rect 109664 139124 110032 139133
rect 109704 139084 109746 139124
rect 109786 139084 109828 139124
rect 109868 139084 109910 139124
rect 109950 139084 109992 139124
rect 109664 139075 110032 139084
rect 124784 139124 125152 139133
rect 124824 139084 124866 139124
rect 124906 139084 124948 139124
rect 124988 139084 125030 139124
rect 125070 139084 125112 139124
rect 124784 139075 125152 139084
rect 139904 139124 140272 139133
rect 139944 139084 139986 139124
rect 140026 139084 140068 139124
rect 140108 139084 140150 139124
rect 140190 139084 140232 139124
rect 139904 139075 140272 139084
rect 78184 138368 78552 138377
rect 78224 138328 78266 138368
rect 78306 138328 78348 138368
rect 78388 138328 78430 138368
rect 78470 138328 78512 138368
rect 78184 138319 78552 138328
rect 93304 138368 93672 138377
rect 93344 138328 93386 138368
rect 93426 138328 93468 138368
rect 93508 138328 93550 138368
rect 93590 138328 93632 138368
rect 93304 138319 93672 138328
rect 108424 138368 108792 138377
rect 108464 138328 108506 138368
rect 108546 138328 108588 138368
rect 108628 138328 108670 138368
rect 108710 138328 108752 138368
rect 108424 138319 108792 138328
rect 123544 138368 123912 138377
rect 123584 138328 123626 138368
rect 123666 138328 123708 138368
rect 123748 138328 123790 138368
rect 123830 138328 123872 138368
rect 123544 138319 123912 138328
rect 138664 138368 139032 138377
rect 138704 138328 138746 138368
rect 138786 138328 138828 138368
rect 138868 138328 138910 138368
rect 138950 138328 138992 138368
rect 138664 138319 139032 138328
rect 79424 137612 79792 137621
rect 79464 137572 79506 137612
rect 79546 137572 79588 137612
rect 79628 137572 79670 137612
rect 79710 137572 79752 137612
rect 79424 137563 79792 137572
rect 94544 137612 94912 137621
rect 94584 137572 94626 137612
rect 94666 137572 94708 137612
rect 94748 137572 94790 137612
rect 94830 137572 94872 137612
rect 94544 137563 94912 137572
rect 109664 137612 110032 137621
rect 109704 137572 109746 137612
rect 109786 137572 109828 137612
rect 109868 137572 109910 137612
rect 109950 137572 109992 137612
rect 109664 137563 110032 137572
rect 124784 137612 125152 137621
rect 124824 137572 124866 137612
rect 124906 137572 124948 137612
rect 124988 137572 125030 137612
rect 125070 137572 125112 137612
rect 124784 137563 125152 137572
rect 139904 137612 140272 137621
rect 139944 137572 139986 137612
rect 140026 137572 140068 137612
rect 140108 137572 140150 137612
rect 140190 137572 140232 137612
rect 139904 137563 140272 137572
rect 78184 136856 78552 136865
rect 78224 136816 78266 136856
rect 78306 136816 78348 136856
rect 78388 136816 78430 136856
rect 78470 136816 78512 136856
rect 78184 136807 78552 136816
rect 93304 136856 93672 136865
rect 93344 136816 93386 136856
rect 93426 136816 93468 136856
rect 93508 136816 93550 136856
rect 93590 136816 93632 136856
rect 93304 136807 93672 136816
rect 108424 136856 108792 136865
rect 108464 136816 108506 136856
rect 108546 136816 108588 136856
rect 108628 136816 108670 136856
rect 108710 136816 108752 136856
rect 108424 136807 108792 136816
rect 123544 136856 123912 136865
rect 123584 136816 123626 136856
rect 123666 136816 123708 136856
rect 123748 136816 123790 136856
rect 123830 136816 123872 136856
rect 123544 136807 123912 136816
rect 138664 136856 139032 136865
rect 138704 136816 138746 136856
rect 138786 136816 138828 136856
rect 138868 136816 138910 136856
rect 138950 136816 138992 136856
rect 138664 136807 139032 136816
rect 79424 136100 79792 136109
rect 79464 136060 79506 136100
rect 79546 136060 79588 136100
rect 79628 136060 79670 136100
rect 79710 136060 79752 136100
rect 79424 136051 79792 136060
rect 94544 136100 94912 136109
rect 94584 136060 94626 136100
rect 94666 136060 94708 136100
rect 94748 136060 94790 136100
rect 94830 136060 94872 136100
rect 94544 136051 94912 136060
rect 109664 136100 110032 136109
rect 109704 136060 109746 136100
rect 109786 136060 109828 136100
rect 109868 136060 109910 136100
rect 109950 136060 109992 136100
rect 109664 136051 110032 136060
rect 124784 136100 125152 136109
rect 124824 136060 124866 136100
rect 124906 136060 124948 136100
rect 124988 136060 125030 136100
rect 125070 136060 125112 136100
rect 124784 136051 125152 136060
rect 139904 136100 140272 136109
rect 139944 136060 139986 136100
rect 140026 136060 140068 136100
rect 140108 136060 140150 136100
rect 140190 136060 140232 136100
rect 139904 136051 140272 136060
rect 78184 135344 78552 135353
rect 78224 135304 78266 135344
rect 78306 135304 78348 135344
rect 78388 135304 78430 135344
rect 78470 135304 78512 135344
rect 78184 135295 78552 135304
rect 93304 135344 93672 135353
rect 93344 135304 93386 135344
rect 93426 135304 93468 135344
rect 93508 135304 93550 135344
rect 93590 135304 93632 135344
rect 93304 135295 93672 135304
rect 108424 135344 108792 135353
rect 108464 135304 108506 135344
rect 108546 135304 108588 135344
rect 108628 135304 108670 135344
rect 108710 135304 108752 135344
rect 108424 135295 108792 135304
rect 123544 135344 123912 135353
rect 123584 135304 123626 135344
rect 123666 135304 123708 135344
rect 123748 135304 123790 135344
rect 123830 135304 123872 135344
rect 123544 135295 123912 135304
rect 138664 135344 139032 135353
rect 138704 135304 138746 135344
rect 138786 135304 138828 135344
rect 138868 135304 138910 135344
rect 138950 135304 138992 135344
rect 138664 135295 139032 135304
rect 79424 134588 79792 134597
rect 79464 134548 79506 134588
rect 79546 134548 79588 134588
rect 79628 134548 79670 134588
rect 79710 134548 79752 134588
rect 79424 134539 79792 134548
rect 94544 134588 94912 134597
rect 94584 134548 94626 134588
rect 94666 134548 94708 134588
rect 94748 134548 94790 134588
rect 94830 134548 94872 134588
rect 94544 134539 94912 134548
rect 109664 134588 110032 134597
rect 109704 134548 109746 134588
rect 109786 134548 109828 134588
rect 109868 134548 109910 134588
rect 109950 134548 109992 134588
rect 109664 134539 110032 134548
rect 124784 134588 125152 134597
rect 124824 134548 124866 134588
rect 124906 134548 124948 134588
rect 124988 134548 125030 134588
rect 125070 134548 125112 134588
rect 124784 134539 125152 134548
rect 139904 134588 140272 134597
rect 139944 134548 139986 134588
rect 140026 134548 140068 134588
rect 140108 134548 140150 134588
rect 140190 134548 140232 134588
rect 139904 134539 140272 134548
rect 78184 133832 78552 133841
rect 78224 133792 78266 133832
rect 78306 133792 78348 133832
rect 78388 133792 78430 133832
rect 78470 133792 78512 133832
rect 78184 133783 78552 133792
rect 93304 133832 93672 133841
rect 93344 133792 93386 133832
rect 93426 133792 93468 133832
rect 93508 133792 93550 133832
rect 93590 133792 93632 133832
rect 93304 133783 93672 133792
rect 108424 133832 108792 133841
rect 108464 133792 108506 133832
rect 108546 133792 108588 133832
rect 108628 133792 108670 133832
rect 108710 133792 108752 133832
rect 108424 133783 108792 133792
rect 123544 133832 123912 133841
rect 123584 133792 123626 133832
rect 123666 133792 123708 133832
rect 123748 133792 123790 133832
rect 123830 133792 123872 133832
rect 123544 133783 123912 133792
rect 138664 133832 139032 133841
rect 138704 133792 138746 133832
rect 138786 133792 138828 133832
rect 138868 133792 138910 133832
rect 138950 133792 138992 133832
rect 138664 133783 139032 133792
rect 79424 133076 79792 133085
rect 79464 133036 79506 133076
rect 79546 133036 79588 133076
rect 79628 133036 79670 133076
rect 79710 133036 79752 133076
rect 79424 133027 79792 133036
rect 94544 133076 94912 133085
rect 94584 133036 94626 133076
rect 94666 133036 94708 133076
rect 94748 133036 94790 133076
rect 94830 133036 94872 133076
rect 94544 133027 94912 133036
rect 109664 133076 110032 133085
rect 109704 133036 109746 133076
rect 109786 133036 109828 133076
rect 109868 133036 109910 133076
rect 109950 133036 109992 133076
rect 109664 133027 110032 133036
rect 124784 133076 125152 133085
rect 124824 133036 124866 133076
rect 124906 133036 124948 133076
rect 124988 133036 125030 133076
rect 125070 133036 125112 133076
rect 124784 133027 125152 133036
rect 139904 133076 140272 133085
rect 139944 133036 139986 133076
rect 140026 133036 140068 133076
rect 140108 133036 140150 133076
rect 140190 133036 140232 133076
rect 139904 133027 140272 133036
rect 78184 132320 78552 132329
rect 78224 132280 78266 132320
rect 78306 132280 78348 132320
rect 78388 132280 78430 132320
rect 78470 132280 78512 132320
rect 78184 132271 78552 132280
rect 93304 132320 93672 132329
rect 93344 132280 93386 132320
rect 93426 132280 93468 132320
rect 93508 132280 93550 132320
rect 93590 132280 93632 132320
rect 93304 132271 93672 132280
rect 108424 132320 108792 132329
rect 108464 132280 108506 132320
rect 108546 132280 108588 132320
rect 108628 132280 108670 132320
rect 108710 132280 108752 132320
rect 108424 132271 108792 132280
rect 123544 132320 123912 132329
rect 123584 132280 123626 132320
rect 123666 132280 123708 132320
rect 123748 132280 123790 132320
rect 123830 132280 123872 132320
rect 123544 132271 123912 132280
rect 138664 132320 139032 132329
rect 138704 132280 138746 132320
rect 138786 132280 138828 132320
rect 138868 132280 138910 132320
rect 138950 132280 138992 132320
rect 138664 132271 139032 132280
rect 79424 131564 79792 131573
rect 79464 131524 79506 131564
rect 79546 131524 79588 131564
rect 79628 131524 79670 131564
rect 79710 131524 79752 131564
rect 79424 131515 79792 131524
rect 94544 131564 94912 131573
rect 94584 131524 94626 131564
rect 94666 131524 94708 131564
rect 94748 131524 94790 131564
rect 94830 131524 94872 131564
rect 94544 131515 94912 131524
rect 109664 131564 110032 131573
rect 109704 131524 109746 131564
rect 109786 131524 109828 131564
rect 109868 131524 109910 131564
rect 109950 131524 109992 131564
rect 109664 131515 110032 131524
rect 124784 131564 125152 131573
rect 124824 131524 124866 131564
rect 124906 131524 124948 131564
rect 124988 131524 125030 131564
rect 125070 131524 125112 131564
rect 124784 131515 125152 131524
rect 139904 131564 140272 131573
rect 139944 131524 139986 131564
rect 140026 131524 140068 131564
rect 140108 131524 140150 131564
rect 140190 131524 140232 131564
rect 139904 131515 140272 131524
rect 78184 130808 78552 130817
rect 78224 130768 78266 130808
rect 78306 130768 78348 130808
rect 78388 130768 78430 130808
rect 78470 130768 78512 130808
rect 78184 130759 78552 130768
rect 93304 130808 93672 130817
rect 93344 130768 93386 130808
rect 93426 130768 93468 130808
rect 93508 130768 93550 130808
rect 93590 130768 93632 130808
rect 93304 130759 93672 130768
rect 108424 130808 108792 130817
rect 108464 130768 108506 130808
rect 108546 130768 108588 130808
rect 108628 130768 108670 130808
rect 108710 130768 108752 130808
rect 108424 130759 108792 130768
rect 123544 130808 123912 130817
rect 123584 130768 123626 130808
rect 123666 130768 123708 130808
rect 123748 130768 123790 130808
rect 123830 130768 123872 130808
rect 123544 130759 123912 130768
rect 138664 130808 139032 130817
rect 138704 130768 138746 130808
rect 138786 130768 138828 130808
rect 138868 130768 138910 130808
rect 138950 130768 138992 130808
rect 138664 130759 139032 130768
rect 79424 130052 79792 130061
rect 79464 130012 79506 130052
rect 79546 130012 79588 130052
rect 79628 130012 79670 130052
rect 79710 130012 79752 130052
rect 79424 130003 79792 130012
rect 94544 130052 94912 130061
rect 94584 130012 94626 130052
rect 94666 130012 94708 130052
rect 94748 130012 94790 130052
rect 94830 130012 94872 130052
rect 94544 130003 94912 130012
rect 109664 130052 110032 130061
rect 109704 130012 109746 130052
rect 109786 130012 109828 130052
rect 109868 130012 109910 130052
rect 109950 130012 109992 130052
rect 109664 130003 110032 130012
rect 124784 130052 125152 130061
rect 124824 130012 124866 130052
rect 124906 130012 124948 130052
rect 124988 130012 125030 130052
rect 125070 130012 125112 130052
rect 124784 130003 125152 130012
rect 139904 130052 140272 130061
rect 139944 130012 139986 130052
rect 140026 130012 140068 130052
rect 140108 130012 140150 130052
rect 140190 130012 140232 130052
rect 139904 130003 140272 130012
rect 78184 129296 78552 129305
rect 78224 129256 78266 129296
rect 78306 129256 78348 129296
rect 78388 129256 78430 129296
rect 78470 129256 78512 129296
rect 78184 129247 78552 129256
rect 93304 129296 93672 129305
rect 93344 129256 93386 129296
rect 93426 129256 93468 129296
rect 93508 129256 93550 129296
rect 93590 129256 93632 129296
rect 93304 129247 93672 129256
rect 108424 129296 108792 129305
rect 108464 129256 108506 129296
rect 108546 129256 108588 129296
rect 108628 129256 108670 129296
rect 108710 129256 108752 129296
rect 108424 129247 108792 129256
rect 123544 129296 123912 129305
rect 123584 129256 123626 129296
rect 123666 129256 123708 129296
rect 123748 129256 123790 129296
rect 123830 129256 123872 129296
rect 123544 129247 123912 129256
rect 138664 129296 139032 129305
rect 138704 129256 138746 129296
rect 138786 129256 138828 129296
rect 138868 129256 138910 129296
rect 138950 129256 138992 129296
rect 138664 129247 139032 129256
rect 79424 128540 79792 128549
rect 79464 128500 79506 128540
rect 79546 128500 79588 128540
rect 79628 128500 79670 128540
rect 79710 128500 79752 128540
rect 79424 128491 79792 128500
rect 94544 128540 94912 128549
rect 94584 128500 94626 128540
rect 94666 128500 94708 128540
rect 94748 128500 94790 128540
rect 94830 128500 94872 128540
rect 94544 128491 94912 128500
rect 109664 128540 110032 128549
rect 109704 128500 109746 128540
rect 109786 128500 109828 128540
rect 109868 128500 109910 128540
rect 109950 128500 109992 128540
rect 109664 128491 110032 128500
rect 124784 128540 125152 128549
rect 124824 128500 124866 128540
rect 124906 128500 124948 128540
rect 124988 128500 125030 128540
rect 125070 128500 125112 128540
rect 124784 128491 125152 128500
rect 139904 128540 140272 128549
rect 139944 128500 139986 128540
rect 140026 128500 140068 128540
rect 140108 128500 140150 128540
rect 140190 128500 140232 128540
rect 139904 128491 140272 128500
rect 78184 127784 78552 127793
rect 78224 127744 78266 127784
rect 78306 127744 78348 127784
rect 78388 127744 78430 127784
rect 78470 127744 78512 127784
rect 78184 127735 78552 127744
rect 93304 127784 93672 127793
rect 93344 127744 93386 127784
rect 93426 127744 93468 127784
rect 93508 127744 93550 127784
rect 93590 127744 93632 127784
rect 93304 127735 93672 127744
rect 108424 127784 108792 127793
rect 108464 127744 108506 127784
rect 108546 127744 108588 127784
rect 108628 127744 108670 127784
rect 108710 127744 108752 127784
rect 108424 127735 108792 127744
rect 123544 127784 123912 127793
rect 123584 127744 123626 127784
rect 123666 127744 123708 127784
rect 123748 127744 123790 127784
rect 123830 127744 123872 127784
rect 123544 127735 123912 127744
rect 138664 127784 139032 127793
rect 138704 127744 138746 127784
rect 138786 127744 138828 127784
rect 138868 127744 138910 127784
rect 138950 127744 138992 127784
rect 138664 127735 139032 127744
rect 79424 127028 79792 127037
rect 79464 126988 79506 127028
rect 79546 126988 79588 127028
rect 79628 126988 79670 127028
rect 79710 126988 79752 127028
rect 79424 126979 79792 126988
rect 94544 127028 94912 127037
rect 94584 126988 94626 127028
rect 94666 126988 94708 127028
rect 94748 126988 94790 127028
rect 94830 126988 94872 127028
rect 94544 126979 94912 126988
rect 109664 127028 110032 127037
rect 109704 126988 109746 127028
rect 109786 126988 109828 127028
rect 109868 126988 109910 127028
rect 109950 126988 109992 127028
rect 109664 126979 110032 126988
rect 124784 127028 125152 127037
rect 124824 126988 124866 127028
rect 124906 126988 124948 127028
rect 124988 126988 125030 127028
rect 125070 126988 125112 127028
rect 124784 126979 125152 126988
rect 139904 127028 140272 127037
rect 139944 126988 139986 127028
rect 140026 126988 140068 127028
rect 140108 126988 140150 127028
rect 140190 126988 140232 127028
rect 139904 126979 140272 126988
rect 78184 126272 78552 126281
rect 78224 126232 78266 126272
rect 78306 126232 78348 126272
rect 78388 126232 78430 126272
rect 78470 126232 78512 126272
rect 78184 126223 78552 126232
rect 93304 126272 93672 126281
rect 93344 126232 93386 126272
rect 93426 126232 93468 126272
rect 93508 126232 93550 126272
rect 93590 126232 93632 126272
rect 93304 126223 93672 126232
rect 108424 126272 108792 126281
rect 108464 126232 108506 126272
rect 108546 126232 108588 126272
rect 108628 126232 108670 126272
rect 108710 126232 108752 126272
rect 108424 126223 108792 126232
rect 123544 126272 123912 126281
rect 123584 126232 123626 126272
rect 123666 126232 123708 126272
rect 123748 126232 123790 126272
rect 123830 126232 123872 126272
rect 123544 126223 123912 126232
rect 138664 126272 139032 126281
rect 138704 126232 138746 126272
rect 138786 126232 138828 126272
rect 138868 126232 138910 126272
rect 138950 126232 138992 126272
rect 138664 126223 139032 126232
rect 79424 125516 79792 125525
rect 79464 125476 79506 125516
rect 79546 125476 79588 125516
rect 79628 125476 79670 125516
rect 79710 125476 79752 125516
rect 79424 125467 79792 125476
rect 94544 125516 94912 125525
rect 94584 125476 94626 125516
rect 94666 125476 94708 125516
rect 94748 125476 94790 125516
rect 94830 125476 94872 125516
rect 94544 125467 94912 125476
rect 109664 125516 110032 125525
rect 109704 125476 109746 125516
rect 109786 125476 109828 125516
rect 109868 125476 109910 125516
rect 109950 125476 109992 125516
rect 109664 125467 110032 125476
rect 124784 125516 125152 125525
rect 124824 125476 124866 125516
rect 124906 125476 124948 125516
rect 124988 125476 125030 125516
rect 125070 125476 125112 125516
rect 124784 125467 125152 125476
rect 139904 125516 140272 125525
rect 139944 125476 139986 125516
rect 140026 125476 140068 125516
rect 140108 125476 140150 125516
rect 140190 125476 140232 125516
rect 139904 125467 140272 125476
rect 93772 125264 93812 125273
rect 78184 124760 78552 124769
rect 78224 124720 78266 124760
rect 78306 124720 78348 124760
rect 78388 124720 78430 124760
rect 78470 124720 78512 124760
rect 78184 124711 78552 124720
rect 93304 124760 93672 124769
rect 93344 124720 93386 124760
rect 93426 124720 93468 124760
rect 93508 124720 93550 124760
rect 93590 124720 93632 124760
rect 93304 124711 93672 124720
rect 79424 124004 79792 124013
rect 79464 123964 79506 124004
rect 79546 123964 79588 124004
rect 79628 123964 79670 124004
rect 79710 123964 79752 124004
rect 79424 123955 79792 123964
rect 78184 123248 78552 123257
rect 78224 123208 78266 123248
rect 78306 123208 78348 123248
rect 78388 123208 78430 123248
rect 78470 123208 78512 123248
rect 78184 123199 78552 123208
rect 93304 123248 93672 123257
rect 93344 123208 93386 123248
rect 93426 123208 93468 123248
rect 93508 123208 93550 123248
rect 93590 123208 93632 123248
rect 93304 123199 93672 123208
rect 79424 122492 79792 122501
rect 79464 122452 79506 122492
rect 79546 122452 79588 122492
rect 79628 122452 79670 122492
rect 79710 122452 79752 122492
rect 79424 122443 79792 122452
rect 93772 122408 93812 125224
rect 108424 124760 108792 124769
rect 108464 124720 108506 124760
rect 108546 124720 108588 124760
rect 108628 124720 108670 124760
rect 108710 124720 108752 124760
rect 108424 124711 108792 124720
rect 123544 124760 123912 124769
rect 123584 124720 123626 124760
rect 123666 124720 123708 124760
rect 123748 124720 123790 124760
rect 123830 124720 123872 124760
rect 123544 124711 123912 124720
rect 138664 124760 139032 124769
rect 138704 124720 138746 124760
rect 138786 124720 138828 124760
rect 138868 124720 138910 124760
rect 138950 124720 138992 124760
rect 138664 124711 139032 124720
rect 94544 124004 94912 124013
rect 94584 123964 94626 124004
rect 94666 123964 94708 124004
rect 94748 123964 94790 124004
rect 94830 123964 94872 124004
rect 94544 123955 94912 123964
rect 109664 124004 110032 124013
rect 109704 123964 109746 124004
rect 109786 123964 109828 124004
rect 109868 123964 109910 124004
rect 109950 123964 109992 124004
rect 109664 123955 110032 123964
rect 124784 124004 125152 124013
rect 124824 123964 124866 124004
rect 124906 123964 124948 124004
rect 124988 123964 125030 124004
rect 125070 123964 125112 124004
rect 124784 123955 125152 123964
rect 139904 124004 140272 124013
rect 139944 123964 139986 124004
rect 140026 123964 140068 124004
rect 140108 123964 140150 124004
rect 140190 123964 140232 124004
rect 139904 123955 140272 123964
rect 108424 123248 108792 123257
rect 108464 123208 108506 123248
rect 108546 123208 108588 123248
rect 108628 123208 108670 123248
rect 108710 123208 108752 123248
rect 108424 123199 108792 123208
rect 123544 123248 123912 123257
rect 123584 123208 123626 123248
rect 123666 123208 123708 123248
rect 123748 123208 123790 123248
rect 123830 123208 123872 123248
rect 123544 123199 123912 123208
rect 138664 123248 139032 123257
rect 138704 123208 138746 123248
rect 138786 123208 138828 123248
rect 138868 123208 138910 123248
rect 138950 123208 138992 123248
rect 138664 123199 139032 123208
rect 94544 122492 94912 122501
rect 94584 122452 94626 122492
rect 94666 122452 94708 122492
rect 94748 122452 94790 122492
rect 94830 122452 94872 122492
rect 94544 122443 94912 122452
rect 109664 122492 110032 122501
rect 109704 122452 109746 122492
rect 109786 122452 109828 122492
rect 109868 122452 109910 122492
rect 109950 122452 109992 122492
rect 109664 122443 110032 122452
rect 124784 122492 125152 122501
rect 124824 122452 124866 122492
rect 124906 122452 124948 122492
rect 124988 122452 125030 122492
rect 125070 122452 125112 122492
rect 124784 122443 125152 122452
rect 139904 122492 140272 122501
rect 139944 122452 139986 122492
rect 140026 122452 140068 122492
rect 140108 122452 140150 122492
rect 140190 122452 140232 122492
rect 139904 122443 140272 122452
rect 93772 122359 93812 122368
rect 78184 121736 78552 121745
rect 78224 121696 78266 121736
rect 78306 121696 78348 121736
rect 78388 121696 78430 121736
rect 78470 121696 78512 121736
rect 78184 121687 78552 121696
rect 93304 121736 93672 121745
rect 93344 121696 93386 121736
rect 93426 121696 93468 121736
rect 93508 121696 93550 121736
rect 93590 121696 93632 121736
rect 93304 121687 93672 121696
rect 108424 121736 108792 121745
rect 108464 121696 108506 121736
rect 108546 121696 108588 121736
rect 108628 121696 108670 121736
rect 108710 121696 108752 121736
rect 108424 121687 108792 121696
rect 123544 121736 123912 121745
rect 123584 121696 123626 121736
rect 123666 121696 123708 121736
rect 123748 121696 123790 121736
rect 123830 121696 123872 121736
rect 123544 121687 123912 121696
rect 138664 121736 139032 121745
rect 138704 121696 138746 121736
rect 138786 121696 138828 121736
rect 138868 121696 138910 121736
rect 138950 121696 138992 121736
rect 138664 121687 139032 121696
rect 79424 120980 79792 120989
rect 79464 120940 79506 120980
rect 79546 120940 79588 120980
rect 79628 120940 79670 120980
rect 79710 120940 79752 120980
rect 79424 120931 79792 120940
rect 94544 120980 94912 120989
rect 94584 120940 94626 120980
rect 94666 120940 94708 120980
rect 94748 120940 94790 120980
rect 94830 120940 94872 120980
rect 94544 120931 94912 120940
rect 109664 120980 110032 120989
rect 109704 120940 109746 120980
rect 109786 120940 109828 120980
rect 109868 120940 109910 120980
rect 109950 120940 109992 120980
rect 109664 120931 110032 120940
rect 124784 120980 125152 120989
rect 124824 120940 124866 120980
rect 124906 120940 124948 120980
rect 124988 120940 125030 120980
rect 125070 120940 125112 120980
rect 124784 120931 125152 120940
rect 139904 120980 140272 120989
rect 139944 120940 139986 120980
rect 140026 120940 140068 120980
rect 140108 120940 140150 120980
rect 140190 120940 140232 120980
rect 139904 120931 140272 120940
rect 78184 120224 78552 120233
rect 78224 120184 78266 120224
rect 78306 120184 78348 120224
rect 78388 120184 78430 120224
rect 78470 120184 78512 120224
rect 78184 120175 78552 120184
rect 93304 120224 93672 120233
rect 93344 120184 93386 120224
rect 93426 120184 93468 120224
rect 93508 120184 93550 120224
rect 93590 120184 93632 120224
rect 93304 120175 93672 120184
rect 108424 120224 108792 120233
rect 108464 120184 108506 120224
rect 108546 120184 108588 120224
rect 108628 120184 108670 120224
rect 108710 120184 108752 120224
rect 108424 120175 108792 120184
rect 123544 120224 123912 120233
rect 123584 120184 123626 120224
rect 123666 120184 123708 120224
rect 123748 120184 123790 120224
rect 123830 120184 123872 120224
rect 123544 120175 123912 120184
rect 138664 120224 139032 120233
rect 138704 120184 138746 120224
rect 138786 120184 138828 120224
rect 138868 120184 138910 120224
rect 138950 120184 138992 120224
rect 138664 120175 139032 120184
rect 79424 119468 79792 119477
rect 79464 119428 79506 119468
rect 79546 119428 79588 119468
rect 79628 119428 79670 119468
rect 79710 119428 79752 119468
rect 79424 119419 79792 119428
rect 94544 119468 94912 119477
rect 94584 119428 94626 119468
rect 94666 119428 94708 119468
rect 94748 119428 94790 119468
rect 94830 119428 94872 119468
rect 94544 119419 94912 119428
rect 109664 119468 110032 119477
rect 109704 119428 109746 119468
rect 109786 119428 109828 119468
rect 109868 119428 109910 119468
rect 109950 119428 109992 119468
rect 109664 119419 110032 119428
rect 124784 119468 125152 119477
rect 124824 119428 124866 119468
rect 124906 119428 124948 119468
rect 124988 119428 125030 119468
rect 125070 119428 125112 119468
rect 124784 119419 125152 119428
rect 139904 119468 140272 119477
rect 139944 119428 139986 119468
rect 140026 119428 140068 119468
rect 140108 119428 140150 119468
rect 140190 119428 140232 119468
rect 139904 119419 140272 119428
rect 78184 118712 78552 118721
rect 78224 118672 78266 118712
rect 78306 118672 78348 118712
rect 78388 118672 78430 118712
rect 78470 118672 78512 118712
rect 78184 118663 78552 118672
rect 93304 118712 93672 118721
rect 93344 118672 93386 118712
rect 93426 118672 93468 118712
rect 93508 118672 93550 118712
rect 93590 118672 93632 118712
rect 93304 118663 93672 118672
rect 108424 118712 108792 118721
rect 108464 118672 108506 118712
rect 108546 118672 108588 118712
rect 108628 118672 108670 118712
rect 108710 118672 108752 118712
rect 108424 118663 108792 118672
rect 123544 118712 123912 118721
rect 123584 118672 123626 118712
rect 123666 118672 123708 118712
rect 123748 118672 123790 118712
rect 123830 118672 123872 118712
rect 123544 118663 123912 118672
rect 138664 118712 139032 118721
rect 138704 118672 138746 118712
rect 138786 118672 138828 118712
rect 138868 118672 138910 118712
rect 138950 118672 138992 118712
rect 138664 118663 139032 118672
rect 79424 117956 79792 117965
rect 79464 117916 79506 117956
rect 79546 117916 79588 117956
rect 79628 117916 79670 117956
rect 79710 117916 79752 117956
rect 79424 117907 79792 117916
rect 94544 117956 94912 117965
rect 94584 117916 94626 117956
rect 94666 117916 94708 117956
rect 94748 117916 94790 117956
rect 94830 117916 94872 117956
rect 94544 117907 94912 117916
rect 109664 117956 110032 117965
rect 109704 117916 109746 117956
rect 109786 117916 109828 117956
rect 109868 117916 109910 117956
rect 109950 117916 109992 117956
rect 109664 117907 110032 117916
rect 124784 117956 125152 117965
rect 124824 117916 124866 117956
rect 124906 117916 124948 117956
rect 124988 117916 125030 117956
rect 125070 117916 125112 117956
rect 124784 117907 125152 117916
rect 139904 117956 140272 117965
rect 139944 117916 139986 117956
rect 140026 117916 140068 117956
rect 140108 117916 140150 117956
rect 140190 117916 140232 117956
rect 139904 117907 140272 117916
rect 78184 117200 78552 117209
rect 78224 117160 78266 117200
rect 78306 117160 78348 117200
rect 78388 117160 78430 117200
rect 78470 117160 78512 117200
rect 78184 117151 78552 117160
rect 93304 117200 93672 117209
rect 93344 117160 93386 117200
rect 93426 117160 93468 117200
rect 93508 117160 93550 117200
rect 93590 117160 93632 117200
rect 93304 117151 93672 117160
rect 108424 117200 108792 117209
rect 108464 117160 108506 117200
rect 108546 117160 108588 117200
rect 108628 117160 108670 117200
rect 108710 117160 108752 117200
rect 108424 117151 108792 117160
rect 123544 117200 123912 117209
rect 123584 117160 123626 117200
rect 123666 117160 123708 117200
rect 123748 117160 123790 117200
rect 123830 117160 123872 117200
rect 123544 117151 123912 117160
rect 138664 117200 139032 117209
rect 138704 117160 138746 117200
rect 138786 117160 138828 117200
rect 138868 117160 138910 117200
rect 138950 117160 138992 117200
rect 138664 117151 139032 117160
rect 79424 116444 79792 116453
rect 79464 116404 79506 116444
rect 79546 116404 79588 116444
rect 79628 116404 79670 116444
rect 79710 116404 79752 116444
rect 79424 116395 79792 116404
rect 94544 116444 94912 116453
rect 94584 116404 94626 116444
rect 94666 116404 94708 116444
rect 94748 116404 94790 116444
rect 94830 116404 94872 116444
rect 94544 116395 94912 116404
rect 109664 116444 110032 116453
rect 109704 116404 109746 116444
rect 109786 116404 109828 116444
rect 109868 116404 109910 116444
rect 109950 116404 109992 116444
rect 109664 116395 110032 116404
rect 124784 116444 125152 116453
rect 124824 116404 124866 116444
rect 124906 116404 124948 116444
rect 124988 116404 125030 116444
rect 125070 116404 125112 116444
rect 124784 116395 125152 116404
rect 139904 116444 140272 116453
rect 139944 116404 139986 116444
rect 140026 116404 140068 116444
rect 140108 116404 140150 116444
rect 140190 116404 140232 116444
rect 139904 116395 140272 116404
rect 78184 115688 78552 115697
rect 78224 115648 78266 115688
rect 78306 115648 78348 115688
rect 78388 115648 78430 115688
rect 78470 115648 78512 115688
rect 78184 115639 78552 115648
rect 93304 115688 93672 115697
rect 93344 115648 93386 115688
rect 93426 115648 93468 115688
rect 93508 115648 93550 115688
rect 93590 115648 93632 115688
rect 93304 115639 93672 115648
rect 108424 115688 108792 115697
rect 108464 115648 108506 115688
rect 108546 115648 108588 115688
rect 108628 115648 108670 115688
rect 108710 115648 108752 115688
rect 108424 115639 108792 115648
rect 123544 115688 123912 115697
rect 123584 115648 123626 115688
rect 123666 115648 123708 115688
rect 123748 115648 123790 115688
rect 123830 115648 123872 115688
rect 123544 115639 123912 115648
rect 138664 115688 139032 115697
rect 138704 115648 138746 115688
rect 138786 115648 138828 115688
rect 138868 115648 138910 115688
rect 138950 115648 138992 115688
rect 138664 115639 139032 115648
rect 79424 114932 79792 114941
rect 79464 114892 79506 114932
rect 79546 114892 79588 114932
rect 79628 114892 79670 114932
rect 79710 114892 79752 114932
rect 79424 114883 79792 114892
rect 94544 114932 94912 114941
rect 94584 114892 94626 114932
rect 94666 114892 94708 114932
rect 94748 114892 94790 114932
rect 94830 114892 94872 114932
rect 94544 114883 94912 114892
rect 109664 114932 110032 114941
rect 109704 114892 109746 114932
rect 109786 114892 109828 114932
rect 109868 114892 109910 114932
rect 109950 114892 109992 114932
rect 109664 114883 110032 114892
rect 124784 114932 125152 114941
rect 124824 114892 124866 114932
rect 124906 114892 124948 114932
rect 124988 114892 125030 114932
rect 125070 114892 125112 114932
rect 124784 114883 125152 114892
rect 139904 114932 140272 114941
rect 139944 114892 139986 114932
rect 140026 114892 140068 114932
rect 140108 114892 140150 114932
rect 140190 114892 140232 114932
rect 139904 114883 140272 114892
rect 78184 114176 78552 114185
rect 78224 114136 78266 114176
rect 78306 114136 78348 114176
rect 78388 114136 78430 114176
rect 78470 114136 78512 114176
rect 78184 114127 78552 114136
rect 93304 114176 93672 114185
rect 93344 114136 93386 114176
rect 93426 114136 93468 114176
rect 93508 114136 93550 114176
rect 93590 114136 93632 114176
rect 93304 114127 93672 114136
rect 108424 114176 108792 114185
rect 108464 114136 108506 114176
rect 108546 114136 108588 114176
rect 108628 114136 108670 114176
rect 108710 114136 108752 114176
rect 108424 114127 108792 114136
rect 123544 114176 123912 114185
rect 123584 114136 123626 114176
rect 123666 114136 123708 114176
rect 123748 114136 123790 114176
rect 123830 114136 123872 114176
rect 123544 114127 123912 114136
rect 138664 114176 139032 114185
rect 138704 114136 138746 114176
rect 138786 114136 138828 114176
rect 138868 114136 138910 114176
rect 138950 114136 138992 114176
rect 138664 114127 139032 114136
rect 79424 113420 79792 113429
rect 79464 113380 79506 113420
rect 79546 113380 79588 113420
rect 79628 113380 79670 113420
rect 79710 113380 79752 113420
rect 79424 113371 79792 113380
rect 94544 113420 94912 113429
rect 94584 113380 94626 113420
rect 94666 113380 94708 113420
rect 94748 113380 94790 113420
rect 94830 113380 94872 113420
rect 94544 113371 94912 113380
rect 109664 113420 110032 113429
rect 109704 113380 109746 113420
rect 109786 113380 109828 113420
rect 109868 113380 109910 113420
rect 109950 113380 109992 113420
rect 109664 113371 110032 113380
rect 124784 113420 125152 113429
rect 124824 113380 124866 113420
rect 124906 113380 124948 113420
rect 124988 113380 125030 113420
rect 125070 113380 125112 113420
rect 124784 113371 125152 113380
rect 139904 113420 140272 113429
rect 139944 113380 139986 113420
rect 140026 113380 140068 113420
rect 140108 113380 140150 113420
rect 140190 113380 140232 113420
rect 139904 113371 140272 113380
rect 78184 112664 78552 112673
rect 78224 112624 78266 112664
rect 78306 112624 78348 112664
rect 78388 112624 78430 112664
rect 78470 112624 78512 112664
rect 78184 112615 78552 112624
rect 93304 112664 93672 112673
rect 93344 112624 93386 112664
rect 93426 112624 93468 112664
rect 93508 112624 93550 112664
rect 93590 112624 93632 112664
rect 93304 112615 93672 112624
rect 108424 112664 108792 112673
rect 108464 112624 108506 112664
rect 108546 112624 108588 112664
rect 108628 112624 108670 112664
rect 108710 112624 108752 112664
rect 108424 112615 108792 112624
rect 123544 112664 123912 112673
rect 123584 112624 123626 112664
rect 123666 112624 123708 112664
rect 123748 112624 123790 112664
rect 123830 112624 123872 112664
rect 123544 112615 123912 112624
rect 138664 112664 139032 112673
rect 138704 112624 138746 112664
rect 138786 112624 138828 112664
rect 138868 112624 138910 112664
rect 138950 112624 138992 112664
rect 138664 112615 139032 112624
rect 79424 111908 79792 111917
rect 79464 111868 79506 111908
rect 79546 111868 79588 111908
rect 79628 111868 79670 111908
rect 79710 111868 79752 111908
rect 79424 111859 79792 111868
rect 94544 111908 94912 111917
rect 94584 111868 94626 111908
rect 94666 111868 94708 111908
rect 94748 111868 94790 111908
rect 94830 111868 94872 111908
rect 94544 111859 94912 111868
rect 109664 111908 110032 111917
rect 109704 111868 109746 111908
rect 109786 111868 109828 111908
rect 109868 111868 109910 111908
rect 109950 111868 109992 111908
rect 109664 111859 110032 111868
rect 124784 111908 125152 111917
rect 124824 111868 124866 111908
rect 124906 111868 124948 111908
rect 124988 111868 125030 111908
rect 125070 111868 125112 111908
rect 124784 111859 125152 111868
rect 139904 111908 140272 111917
rect 139944 111868 139986 111908
rect 140026 111868 140068 111908
rect 140108 111868 140150 111908
rect 140190 111868 140232 111908
rect 139904 111859 140272 111868
rect 78184 111152 78552 111161
rect 78224 111112 78266 111152
rect 78306 111112 78348 111152
rect 78388 111112 78430 111152
rect 78470 111112 78512 111152
rect 78184 111103 78552 111112
rect 93304 111152 93672 111161
rect 93344 111112 93386 111152
rect 93426 111112 93468 111152
rect 93508 111112 93550 111152
rect 93590 111112 93632 111152
rect 93304 111103 93672 111112
rect 108424 111152 108792 111161
rect 108464 111112 108506 111152
rect 108546 111112 108588 111152
rect 108628 111112 108670 111152
rect 108710 111112 108752 111152
rect 108424 111103 108792 111112
rect 123544 111152 123912 111161
rect 123584 111112 123626 111152
rect 123666 111112 123708 111152
rect 123748 111112 123790 111152
rect 123830 111112 123872 111152
rect 123544 111103 123912 111112
rect 138664 111152 139032 111161
rect 138704 111112 138746 111152
rect 138786 111112 138828 111152
rect 138868 111112 138910 111152
rect 138950 111112 138992 111152
rect 138664 111103 139032 111112
rect 79424 110396 79792 110405
rect 79464 110356 79506 110396
rect 79546 110356 79588 110396
rect 79628 110356 79670 110396
rect 79710 110356 79752 110396
rect 79424 110347 79792 110356
rect 94544 110396 94912 110405
rect 94584 110356 94626 110396
rect 94666 110356 94708 110396
rect 94748 110356 94790 110396
rect 94830 110356 94872 110396
rect 94544 110347 94912 110356
rect 109664 110396 110032 110405
rect 109704 110356 109746 110396
rect 109786 110356 109828 110396
rect 109868 110356 109910 110396
rect 109950 110356 109992 110396
rect 109664 110347 110032 110356
rect 124784 110396 125152 110405
rect 124824 110356 124866 110396
rect 124906 110356 124948 110396
rect 124988 110356 125030 110396
rect 125070 110356 125112 110396
rect 124784 110347 125152 110356
rect 139904 110396 140272 110405
rect 139944 110356 139986 110396
rect 140026 110356 140068 110396
rect 140108 110356 140150 110396
rect 140190 110356 140232 110396
rect 139904 110347 140272 110356
rect 78184 109640 78552 109649
rect 78224 109600 78266 109640
rect 78306 109600 78348 109640
rect 78388 109600 78430 109640
rect 78470 109600 78512 109640
rect 78184 109591 78552 109600
rect 93304 109640 93672 109649
rect 93344 109600 93386 109640
rect 93426 109600 93468 109640
rect 93508 109600 93550 109640
rect 93590 109600 93632 109640
rect 93304 109591 93672 109600
rect 108424 109640 108792 109649
rect 108464 109600 108506 109640
rect 108546 109600 108588 109640
rect 108628 109600 108670 109640
rect 108710 109600 108752 109640
rect 108424 109591 108792 109600
rect 123544 109640 123912 109649
rect 123584 109600 123626 109640
rect 123666 109600 123708 109640
rect 123748 109600 123790 109640
rect 123830 109600 123872 109640
rect 123544 109591 123912 109600
rect 138664 109640 139032 109649
rect 138704 109600 138746 109640
rect 138786 109600 138828 109640
rect 138868 109600 138910 109640
rect 138950 109600 138992 109640
rect 138664 109591 139032 109600
rect 79424 108884 79792 108893
rect 79464 108844 79506 108884
rect 79546 108844 79588 108884
rect 79628 108844 79670 108884
rect 79710 108844 79752 108884
rect 79424 108835 79792 108844
rect 94544 108884 94912 108893
rect 94584 108844 94626 108884
rect 94666 108844 94708 108884
rect 94748 108844 94790 108884
rect 94830 108844 94872 108884
rect 94544 108835 94912 108844
rect 109664 108884 110032 108893
rect 109704 108844 109746 108884
rect 109786 108844 109828 108884
rect 109868 108844 109910 108884
rect 109950 108844 109992 108884
rect 109664 108835 110032 108844
rect 124784 108884 125152 108893
rect 124824 108844 124866 108884
rect 124906 108844 124948 108884
rect 124988 108844 125030 108884
rect 125070 108844 125112 108884
rect 124784 108835 125152 108844
rect 139904 108884 140272 108893
rect 139944 108844 139986 108884
rect 140026 108844 140068 108884
rect 140108 108844 140150 108884
rect 140190 108844 140232 108884
rect 139904 108835 140272 108844
rect 78184 108128 78552 108137
rect 78224 108088 78266 108128
rect 78306 108088 78348 108128
rect 78388 108088 78430 108128
rect 78470 108088 78512 108128
rect 78184 108079 78552 108088
rect 93304 108128 93672 108137
rect 93344 108088 93386 108128
rect 93426 108088 93468 108128
rect 93508 108088 93550 108128
rect 93590 108088 93632 108128
rect 93304 108079 93672 108088
rect 108424 108128 108792 108137
rect 108464 108088 108506 108128
rect 108546 108088 108588 108128
rect 108628 108088 108670 108128
rect 108710 108088 108752 108128
rect 108424 108079 108792 108088
rect 123544 108128 123912 108137
rect 123584 108088 123626 108128
rect 123666 108088 123708 108128
rect 123748 108088 123790 108128
rect 123830 108088 123872 108128
rect 123544 108079 123912 108088
rect 138664 108128 139032 108137
rect 138704 108088 138746 108128
rect 138786 108088 138828 108128
rect 138868 108088 138910 108128
rect 138950 108088 138992 108128
rect 138664 108079 139032 108088
rect 79424 107372 79792 107381
rect 79464 107332 79506 107372
rect 79546 107332 79588 107372
rect 79628 107332 79670 107372
rect 79710 107332 79752 107372
rect 79424 107323 79792 107332
rect 94544 107372 94912 107381
rect 94584 107332 94626 107372
rect 94666 107332 94708 107372
rect 94748 107332 94790 107372
rect 94830 107332 94872 107372
rect 94544 107323 94912 107332
rect 109664 107372 110032 107381
rect 109704 107332 109746 107372
rect 109786 107332 109828 107372
rect 109868 107332 109910 107372
rect 109950 107332 109992 107372
rect 109664 107323 110032 107332
rect 124784 107372 125152 107381
rect 124824 107332 124866 107372
rect 124906 107332 124948 107372
rect 124988 107332 125030 107372
rect 125070 107332 125112 107372
rect 124784 107323 125152 107332
rect 139904 107372 140272 107381
rect 139944 107332 139986 107372
rect 140026 107332 140068 107372
rect 140108 107332 140150 107372
rect 140190 107332 140232 107372
rect 139904 107323 140272 107332
rect 78184 106616 78552 106625
rect 78224 106576 78266 106616
rect 78306 106576 78348 106616
rect 78388 106576 78430 106616
rect 78470 106576 78512 106616
rect 78184 106567 78552 106576
rect 93304 106616 93672 106625
rect 93344 106576 93386 106616
rect 93426 106576 93468 106616
rect 93508 106576 93550 106616
rect 93590 106576 93632 106616
rect 93304 106567 93672 106576
rect 108424 106616 108792 106625
rect 108464 106576 108506 106616
rect 108546 106576 108588 106616
rect 108628 106576 108670 106616
rect 108710 106576 108752 106616
rect 108424 106567 108792 106576
rect 123544 106616 123912 106625
rect 123584 106576 123626 106616
rect 123666 106576 123708 106616
rect 123748 106576 123790 106616
rect 123830 106576 123872 106616
rect 123544 106567 123912 106576
rect 138664 106616 139032 106625
rect 138704 106576 138746 106616
rect 138786 106576 138828 106616
rect 138868 106576 138910 106616
rect 138950 106576 138992 106616
rect 138664 106567 139032 106576
rect 79424 105860 79792 105869
rect 79464 105820 79506 105860
rect 79546 105820 79588 105860
rect 79628 105820 79670 105860
rect 79710 105820 79752 105860
rect 79424 105811 79792 105820
rect 94544 105860 94912 105869
rect 94584 105820 94626 105860
rect 94666 105820 94708 105860
rect 94748 105820 94790 105860
rect 94830 105820 94872 105860
rect 94544 105811 94912 105820
rect 109664 105860 110032 105869
rect 109704 105820 109746 105860
rect 109786 105820 109828 105860
rect 109868 105820 109910 105860
rect 109950 105820 109992 105860
rect 109664 105811 110032 105820
rect 124784 105860 125152 105869
rect 124824 105820 124866 105860
rect 124906 105820 124948 105860
rect 124988 105820 125030 105860
rect 125070 105820 125112 105860
rect 124784 105811 125152 105820
rect 139904 105860 140272 105869
rect 139944 105820 139986 105860
rect 140026 105820 140068 105860
rect 140108 105820 140150 105860
rect 140190 105820 140232 105860
rect 139904 105811 140272 105820
rect 78184 105104 78552 105113
rect 78224 105064 78266 105104
rect 78306 105064 78348 105104
rect 78388 105064 78430 105104
rect 78470 105064 78512 105104
rect 78184 105055 78552 105064
rect 93304 105104 93672 105113
rect 93344 105064 93386 105104
rect 93426 105064 93468 105104
rect 93508 105064 93550 105104
rect 93590 105064 93632 105104
rect 93304 105055 93672 105064
rect 108424 105104 108792 105113
rect 108464 105064 108506 105104
rect 108546 105064 108588 105104
rect 108628 105064 108670 105104
rect 108710 105064 108752 105104
rect 108424 105055 108792 105064
rect 123544 105104 123912 105113
rect 123584 105064 123626 105104
rect 123666 105064 123708 105104
rect 123748 105064 123790 105104
rect 123830 105064 123872 105104
rect 123544 105055 123912 105064
rect 138664 105104 139032 105113
rect 138704 105064 138746 105104
rect 138786 105064 138828 105104
rect 138868 105064 138910 105104
rect 138950 105064 138992 105104
rect 138664 105055 139032 105064
rect 79424 104348 79792 104357
rect 79464 104308 79506 104348
rect 79546 104308 79588 104348
rect 79628 104308 79670 104348
rect 79710 104308 79752 104348
rect 79424 104299 79792 104308
rect 94544 104348 94912 104357
rect 94584 104308 94626 104348
rect 94666 104308 94708 104348
rect 94748 104308 94790 104348
rect 94830 104308 94872 104348
rect 94544 104299 94912 104308
rect 109664 104348 110032 104357
rect 109704 104308 109746 104348
rect 109786 104308 109828 104348
rect 109868 104308 109910 104348
rect 109950 104308 109992 104348
rect 109664 104299 110032 104308
rect 124784 104348 125152 104357
rect 124824 104308 124866 104348
rect 124906 104308 124948 104348
rect 124988 104308 125030 104348
rect 125070 104308 125112 104348
rect 124784 104299 125152 104308
rect 139904 104348 140272 104357
rect 139944 104308 139986 104348
rect 140026 104308 140068 104348
rect 140108 104308 140150 104348
rect 140190 104308 140232 104348
rect 139904 104299 140272 104308
rect 78184 103592 78552 103601
rect 78224 103552 78266 103592
rect 78306 103552 78348 103592
rect 78388 103552 78430 103592
rect 78470 103552 78512 103592
rect 78184 103543 78552 103552
rect 93304 103592 93672 103601
rect 93344 103552 93386 103592
rect 93426 103552 93468 103592
rect 93508 103552 93550 103592
rect 93590 103552 93632 103592
rect 93304 103543 93672 103552
rect 108424 103592 108792 103601
rect 108464 103552 108506 103592
rect 108546 103552 108588 103592
rect 108628 103552 108670 103592
rect 108710 103552 108752 103592
rect 108424 103543 108792 103552
rect 123544 103592 123912 103601
rect 123584 103552 123626 103592
rect 123666 103552 123708 103592
rect 123748 103552 123790 103592
rect 123830 103552 123872 103592
rect 123544 103543 123912 103552
rect 138664 103592 139032 103601
rect 138704 103552 138746 103592
rect 138786 103552 138828 103592
rect 138868 103552 138910 103592
rect 138950 103552 138992 103592
rect 138664 103543 139032 103552
rect 79424 102836 79792 102845
rect 79464 102796 79506 102836
rect 79546 102796 79588 102836
rect 79628 102796 79670 102836
rect 79710 102796 79752 102836
rect 79424 102787 79792 102796
rect 94544 102836 94912 102845
rect 94584 102796 94626 102836
rect 94666 102796 94708 102836
rect 94748 102796 94790 102836
rect 94830 102796 94872 102836
rect 94544 102787 94912 102796
rect 109664 102836 110032 102845
rect 109704 102796 109746 102836
rect 109786 102796 109828 102836
rect 109868 102796 109910 102836
rect 109950 102796 109992 102836
rect 109664 102787 110032 102796
rect 124784 102836 125152 102845
rect 124824 102796 124866 102836
rect 124906 102796 124948 102836
rect 124988 102796 125030 102836
rect 125070 102796 125112 102836
rect 124784 102787 125152 102796
rect 139904 102836 140272 102845
rect 139944 102796 139986 102836
rect 140026 102796 140068 102836
rect 140108 102796 140150 102836
rect 140190 102796 140232 102836
rect 139904 102787 140272 102796
rect 78184 102080 78552 102089
rect 78224 102040 78266 102080
rect 78306 102040 78348 102080
rect 78388 102040 78430 102080
rect 78470 102040 78512 102080
rect 78184 102031 78552 102040
rect 93304 102080 93672 102089
rect 93344 102040 93386 102080
rect 93426 102040 93468 102080
rect 93508 102040 93550 102080
rect 93590 102040 93632 102080
rect 93304 102031 93672 102040
rect 108424 102080 108792 102089
rect 108464 102040 108506 102080
rect 108546 102040 108588 102080
rect 108628 102040 108670 102080
rect 108710 102040 108752 102080
rect 108424 102031 108792 102040
rect 123544 102080 123912 102089
rect 123584 102040 123626 102080
rect 123666 102040 123708 102080
rect 123748 102040 123790 102080
rect 123830 102040 123872 102080
rect 123544 102031 123912 102040
rect 138664 102080 139032 102089
rect 138704 102040 138746 102080
rect 138786 102040 138828 102080
rect 138868 102040 138910 102080
rect 138950 102040 138992 102080
rect 138664 102031 139032 102040
rect 79424 101324 79792 101333
rect 79464 101284 79506 101324
rect 79546 101284 79588 101324
rect 79628 101284 79670 101324
rect 79710 101284 79752 101324
rect 79424 101275 79792 101284
rect 94544 101324 94912 101333
rect 94584 101284 94626 101324
rect 94666 101284 94708 101324
rect 94748 101284 94790 101324
rect 94830 101284 94872 101324
rect 94544 101275 94912 101284
rect 109664 101324 110032 101333
rect 109704 101284 109746 101324
rect 109786 101284 109828 101324
rect 109868 101284 109910 101324
rect 109950 101284 109992 101324
rect 109664 101275 110032 101284
rect 124784 101324 125152 101333
rect 124824 101284 124866 101324
rect 124906 101284 124948 101324
rect 124988 101284 125030 101324
rect 125070 101284 125112 101324
rect 124784 101275 125152 101284
rect 139904 101324 140272 101333
rect 139944 101284 139986 101324
rect 140026 101284 140068 101324
rect 140108 101284 140150 101324
rect 140190 101284 140232 101324
rect 139904 101275 140272 101284
rect 78184 100568 78552 100577
rect 78224 100528 78266 100568
rect 78306 100528 78348 100568
rect 78388 100528 78430 100568
rect 78470 100528 78512 100568
rect 78184 100519 78552 100528
rect 93304 100568 93672 100577
rect 93344 100528 93386 100568
rect 93426 100528 93468 100568
rect 93508 100528 93550 100568
rect 93590 100528 93632 100568
rect 93304 100519 93672 100528
rect 108424 100568 108792 100577
rect 108464 100528 108506 100568
rect 108546 100528 108588 100568
rect 108628 100528 108670 100568
rect 108710 100528 108752 100568
rect 108424 100519 108792 100528
rect 123544 100568 123912 100577
rect 123584 100528 123626 100568
rect 123666 100528 123708 100568
rect 123748 100528 123790 100568
rect 123830 100528 123872 100568
rect 123544 100519 123912 100528
rect 138664 100568 139032 100577
rect 138704 100528 138746 100568
rect 138786 100528 138828 100568
rect 138868 100528 138910 100568
rect 138950 100528 138992 100568
rect 138664 100519 139032 100528
rect 79424 99812 79792 99821
rect 79464 99772 79506 99812
rect 79546 99772 79588 99812
rect 79628 99772 79670 99812
rect 79710 99772 79752 99812
rect 79424 99763 79792 99772
rect 94544 99812 94912 99821
rect 94584 99772 94626 99812
rect 94666 99772 94708 99812
rect 94748 99772 94790 99812
rect 94830 99772 94872 99812
rect 94544 99763 94912 99772
rect 109664 99812 110032 99821
rect 109704 99772 109746 99812
rect 109786 99772 109828 99812
rect 109868 99772 109910 99812
rect 109950 99772 109992 99812
rect 109664 99763 110032 99772
rect 124784 99812 125152 99821
rect 124824 99772 124866 99812
rect 124906 99772 124948 99812
rect 124988 99772 125030 99812
rect 125070 99772 125112 99812
rect 124784 99763 125152 99772
rect 139904 99812 140272 99821
rect 139944 99772 139986 99812
rect 140026 99772 140068 99812
rect 140108 99772 140150 99812
rect 140190 99772 140232 99812
rect 139904 99763 140272 99772
rect 78184 99056 78552 99065
rect 78224 99016 78266 99056
rect 78306 99016 78348 99056
rect 78388 99016 78430 99056
rect 78470 99016 78512 99056
rect 78184 99007 78552 99016
rect 93304 99056 93672 99065
rect 93344 99016 93386 99056
rect 93426 99016 93468 99056
rect 93508 99016 93550 99056
rect 93590 99016 93632 99056
rect 93304 99007 93672 99016
rect 108424 99056 108792 99065
rect 108464 99016 108506 99056
rect 108546 99016 108588 99056
rect 108628 99016 108670 99056
rect 108710 99016 108752 99056
rect 108424 99007 108792 99016
rect 123544 99056 123912 99065
rect 123584 99016 123626 99056
rect 123666 99016 123708 99056
rect 123748 99016 123790 99056
rect 123830 99016 123872 99056
rect 123544 99007 123912 99016
rect 138664 99056 139032 99065
rect 138704 99016 138746 99056
rect 138786 99016 138828 99056
rect 138868 99016 138910 99056
rect 138950 99016 138992 99056
rect 138664 99007 139032 99016
rect 79424 98300 79792 98309
rect 79464 98260 79506 98300
rect 79546 98260 79588 98300
rect 79628 98260 79670 98300
rect 79710 98260 79752 98300
rect 79424 98251 79792 98260
rect 94544 98300 94912 98309
rect 94584 98260 94626 98300
rect 94666 98260 94708 98300
rect 94748 98260 94790 98300
rect 94830 98260 94872 98300
rect 94544 98251 94912 98260
rect 109664 98300 110032 98309
rect 109704 98260 109746 98300
rect 109786 98260 109828 98300
rect 109868 98260 109910 98300
rect 109950 98260 109992 98300
rect 109664 98251 110032 98260
rect 124784 98300 125152 98309
rect 124824 98260 124866 98300
rect 124906 98260 124948 98300
rect 124988 98260 125030 98300
rect 125070 98260 125112 98300
rect 124784 98251 125152 98260
rect 139904 98300 140272 98309
rect 139944 98260 139986 98300
rect 140026 98260 140068 98300
rect 140108 98260 140150 98300
rect 140190 98260 140232 98300
rect 139904 98251 140272 98260
rect 78184 97544 78552 97553
rect 78224 97504 78266 97544
rect 78306 97504 78348 97544
rect 78388 97504 78430 97544
rect 78470 97504 78512 97544
rect 78184 97495 78552 97504
rect 93304 97544 93672 97553
rect 93344 97504 93386 97544
rect 93426 97504 93468 97544
rect 93508 97504 93550 97544
rect 93590 97504 93632 97544
rect 93304 97495 93672 97504
rect 108424 97544 108792 97553
rect 108464 97504 108506 97544
rect 108546 97504 108588 97544
rect 108628 97504 108670 97544
rect 108710 97504 108752 97544
rect 108424 97495 108792 97504
rect 123544 97544 123912 97553
rect 123584 97504 123626 97544
rect 123666 97504 123708 97544
rect 123748 97504 123790 97544
rect 123830 97504 123872 97544
rect 123544 97495 123912 97504
rect 138664 97544 139032 97553
rect 138704 97504 138746 97544
rect 138786 97504 138828 97544
rect 138868 97504 138910 97544
rect 138950 97504 138992 97544
rect 138664 97495 139032 97504
rect 79424 96788 79792 96797
rect 79464 96748 79506 96788
rect 79546 96748 79588 96788
rect 79628 96748 79670 96788
rect 79710 96748 79752 96788
rect 79424 96739 79792 96748
rect 94544 96788 94912 96797
rect 94584 96748 94626 96788
rect 94666 96748 94708 96788
rect 94748 96748 94790 96788
rect 94830 96748 94872 96788
rect 94544 96739 94912 96748
rect 109664 96788 110032 96797
rect 109704 96748 109746 96788
rect 109786 96748 109828 96788
rect 109868 96748 109910 96788
rect 109950 96748 109992 96788
rect 109664 96739 110032 96748
rect 124784 96788 125152 96797
rect 124824 96748 124866 96788
rect 124906 96748 124948 96788
rect 124988 96748 125030 96788
rect 125070 96748 125112 96788
rect 124784 96739 125152 96748
rect 139904 96788 140272 96797
rect 139944 96748 139986 96788
rect 140026 96748 140068 96788
rect 140108 96748 140150 96788
rect 140190 96748 140232 96788
rect 139904 96739 140272 96748
rect 78184 96032 78552 96041
rect 78224 95992 78266 96032
rect 78306 95992 78348 96032
rect 78388 95992 78430 96032
rect 78470 95992 78512 96032
rect 78184 95983 78552 95992
rect 93304 96032 93672 96041
rect 93344 95992 93386 96032
rect 93426 95992 93468 96032
rect 93508 95992 93550 96032
rect 93590 95992 93632 96032
rect 93304 95983 93672 95992
rect 108424 96032 108792 96041
rect 108464 95992 108506 96032
rect 108546 95992 108588 96032
rect 108628 95992 108670 96032
rect 108710 95992 108752 96032
rect 108424 95983 108792 95992
rect 123544 96032 123912 96041
rect 123584 95992 123626 96032
rect 123666 95992 123708 96032
rect 123748 95992 123790 96032
rect 123830 95992 123872 96032
rect 123544 95983 123912 95992
rect 138664 96032 139032 96041
rect 138704 95992 138746 96032
rect 138786 95992 138828 96032
rect 138868 95992 138910 96032
rect 138950 95992 138992 96032
rect 138664 95983 139032 95992
rect 79424 95276 79792 95285
rect 79464 95236 79506 95276
rect 79546 95236 79588 95276
rect 79628 95236 79670 95276
rect 79710 95236 79752 95276
rect 79424 95227 79792 95236
rect 94544 95276 94912 95285
rect 94584 95236 94626 95276
rect 94666 95236 94708 95276
rect 94748 95236 94790 95276
rect 94830 95236 94872 95276
rect 94544 95227 94912 95236
rect 109664 95276 110032 95285
rect 109704 95236 109746 95276
rect 109786 95236 109828 95276
rect 109868 95236 109910 95276
rect 109950 95236 109992 95276
rect 109664 95227 110032 95236
rect 124784 95276 125152 95285
rect 124824 95236 124866 95276
rect 124906 95236 124948 95276
rect 124988 95236 125030 95276
rect 125070 95236 125112 95276
rect 124784 95227 125152 95236
rect 139904 95276 140272 95285
rect 139944 95236 139986 95276
rect 140026 95236 140068 95276
rect 140108 95236 140150 95276
rect 140190 95236 140232 95276
rect 139904 95227 140272 95236
rect 78184 94520 78552 94529
rect 78224 94480 78266 94520
rect 78306 94480 78348 94520
rect 78388 94480 78430 94520
rect 78470 94480 78512 94520
rect 78184 94471 78552 94480
rect 93304 94520 93672 94529
rect 93344 94480 93386 94520
rect 93426 94480 93468 94520
rect 93508 94480 93550 94520
rect 93590 94480 93632 94520
rect 93304 94471 93672 94480
rect 108424 94520 108792 94529
rect 108464 94480 108506 94520
rect 108546 94480 108588 94520
rect 108628 94480 108670 94520
rect 108710 94480 108752 94520
rect 108424 94471 108792 94480
rect 123544 94520 123912 94529
rect 123584 94480 123626 94520
rect 123666 94480 123708 94520
rect 123748 94480 123790 94520
rect 123830 94480 123872 94520
rect 123544 94471 123912 94480
rect 138664 94520 139032 94529
rect 138704 94480 138746 94520
rect 138786 94480 138828 94520
rect 138868 94480 138910 94520
rect 138950 94480 138992 94520
rect 138664 94471 139032 94480
rect 79424 93764 79792 93773
rect 79464 93724 79506 93764
rect 79546 93724 79588 93764
rect 79628 93724 79670 93764
rect 79710 93724 79752 93764
rect 79424 93715 79792 93724
rect 94544 93764 94912 93773
rect 94584 93724 94626 93764
rect 94666 93724 94708 93764
rect 94748 93724 94790 93764
rect 94830 93724 94872 93764
rect 94544 93715 94912 93724
rect 109664 93764 110032 93773
rect 109704 93724 109746 93764
rect 109786 93724 109828 93764
rect 109868 93724 109910 93764
rect 109950 93724 109992 93764
rect 109664 93715 110032 93724
rect 124784 93764 125152 93773
rect 124824 93724 124866 93764
rect 124906 93724 124948 93764
rect 124988 93724 125030 93764
rect 125070 93724 125112 93764
rect 124784 93715 125152 93724
rect 139904 93764 140272 93773
rect 139944 93724 139986 93764
rect 140026 93724 140068 93764
rect 140108 93724 140150 93764
rect 140190 93724 140232 93764
rect 139904 93715 140272 93724
rect 78184 93008 78552 93017
rect 78224 92968 78266 93008
rect 78306 92968 78348 93008
rect 78388 92968 78430 93008
rect 78470 92968 78512 93008
rect 78184 92959 78552 92968
rect 93304 93008 93672 93017
rect 93344 92968 93386 93008
rect 93426 92968 93468 93008
rect 93508 92968 93550 93008
rect 93590 92968 93632 93008
rect 93304 92959 93672 92968
rect 108424 93008 108792 93017
rect 108464 92968 108506 93008
rect 108546 92968 108588 93008
rect 108628 92968 108670 93008
rect 108710 92968 108752 93008
rect 108424 92959 108792 92968
rect 123544 93008 123912 93017
rect 123584 92968 123626 93008
rect 123666 92968 123708 93008
rect 123748 92968 123790 93008
rect 123830 92968 123872 93008
rect 123544 92959 123912 92968
rect 138664 93008 139032 93017
rect 138704 92968 138746 93008
rect 138786 92968 138828 93008
rect 138868 92968 138910 93008
rect 138950 92968 138992 93008
rect 138664 92959 139032 92968
rect 79424 92252 79792 92261
rect 79464 92212 79506 92252
rect 79546 92212 79588 92252
rect 79628 92212 79670 92252
rect 79710 92212 79752 92252
rect 79424 92203 79792 92212
rect 94544 92252 94912 92261
rect 94584 92212 94626 92252
rect 94666 92212 94708 92252
rect 94748 92212 94790 92252
rect 94830 92212 94872 92252
rect 94544 92203 94912 92212
rect 109664 92252 110032 92261
rect 109704 92212 109746 92252
rect 109786 92212 109828 92252
rect 109868 92212 109910 92252
rect 109950 92212 109992 92252
rect 109664 92203 110032 92212
rect 124784 92252 125152 92261
rect 124824 92212 124866 92252
rect 124906 92212 124948 92252
rect 124988 92212 125030 92252
rect 125070 92212 125112 92252
rect 124784 92203 125152 92212
rect 139904 92252 140272 92261
rect 139944 92212 139986 92252
rect 140026 92212 140068 92252
rect 140108 92212 140150 92252
rect 140190 92212 140232 92252
rect 139904 92203 140272 92212
rect 78184 91496 78552 91505
rect 78224 91456 78266 91496
rect 78306 91456 78348 91496
rect 78388 91456 78430 91496
rect 78470 91456 78512 91496
rect 78184 91447 78552 91456
rect 93304 91496 93672 91505
rect 93344 91456 93386 91496
rect 93426 91456 93468 91496
rect 93508 91456 93550 91496
rect 93590 91456 93632 91496
rect 93304 91447 93672 91456
rect 108424 91496 108792 91505
rect 108464 91456 108506 91496
rect 108546 91456 108588 91496
rect 108628 91456 108670 91496
rect 108710 91456 108752 91496
rect 108424 91447 108792 91456
rect 123544 91496 123912 91505
rect 123584 91456 123626 91496
rect 123666 91456 123708 91496
rect 123748 91456 123790 91496
rect 123830 91456 123872 91496
rect 123544 91447 123912 91456
rect 138664 91496 139032 91505
rect 138704 91456 138746 91496
rect 138786 91456 138828 91496
rect 138868 91456 138910 91496
rect 138950 91456 138992 91496
rect 138664 91447 139032 91456
rect 79424 90740 79792 90749
rect 79464 90700 79506 90740
rect 79546 90700 79588 90740
rect 79628 90700 79670 90740
rect 79710 90700 79752 90740
rect 79424 90691 79792 90700
rect 94544 90740 94912 90749
rect 94584 90700 94626 90740
rect 94666 90700 94708 90740
rect 94748 90700 94790 90740
rect 94830 90700 94872 90740
rect 94544 90691 94912 90700
rect 109664 90740 110032 90749
rect 109704 90700 109746 90740
rect 109786 90700 109828 90740
rect 109868 90700 109910 90740
rect 109950 90700 109992 90740
rect 109664 90691 110032 90700
rect 124784 90740 125152 90749
rect 124824 90700 124866 90740
rect 124906 90700 124948 90740
rect 124988 90700 125030 90740
rect 125070 90700 125112 90740
rect 124784 90691 125152 90700
rect 139904 90740 140272 90749
rect 139944 90700 139986 90740
rect 140026 90700 140068 90740
rect 140108 90700 140150 90740
rect 140190 90700 140232 90740
rect 139904 90691 140272 90700
rect 78184 89984 78552 89993
rect 78224 89944 78266 89984
rect 78306 89944 78348 89984
rect 78388 89944 78430 89984
rect 78470 89944 78512 89984
rect 78184 89935 78552 89944
rect 93304 89984 93672 89993
rect 93344 89944 93386 89984
rect 93426 89944 93468 89984
rect 93508 89944 93550 89984
rect 93590 89944 93632 89984
rect 93304 89935 93672 89944
rect 108424 89984 108792 89993
rect 108464 89944 108506 89984
rect 108546 89944 108588 89984
rect 108628 89944 108670 89984
rect 108710 89944 108752 89984
rect 108424 89935 108792 89944
rect 123544 89984 123912 89993
rect 123584 89944 123626 89984
rect 123666 89944 123708 89984
rect 123748 89944 123790 89984
rect 123830 89944 123872 89984
rect 123544 89935 123912 89944
rect 138664 89984 139032 89993
rect 138704 89944 138746 89984
rect 138786 89944 138828 89984
rect 138868 89944 138910 89984
rect 138950 89944 138992 89984
rect 138664 89935 139032 89944
rect 79424 89228 79792 89237
rect 79464 89188 79506 89228
rect 79546 89188 79588 89228
rect 79628 89188 79670 89228
rect 79710 89188 79752 89228
rect 79424 89179 79792 89188
rect 94544 89228 94912 89237
rect 94584 89188 94626 89228
rect 94666 89188 94708 89228
rect 94748 89188 94790 89228
rect 94830 89188 94872 89228
rect 94544 89179 94912 89188
rect 109664 89228 110032 89237
rect 109704 89188 109746 89228
rect 109786 89188 109828 89228
rect 109868 89188 109910 89228
rect 109950 89188 109992 89228
rect 109664 89179 110032 89188
rect 124784 89228 125152 89237
rect 124824 89188 124866 89228
rect 124906 89188 124948 89228
rect 124988 89188 125030 89228
rect 125070 89188 125112 89228
rect 124784 89179 125152 89188
rect 139904 89228 140272 89237
rect 139944 89188 139986 89228
rect 140026 89188 140068 89228
rect 140108 89188 140150 89228
rect 140190 89188 140232 89228
rect 139904 89179 140272 89188
rect 90699 89144 90741 89153
rect 90699 89104 90700 89144
rect 90740 89104 90741 89144
rect 90699 89095 90741 89104
rect 92139 89144 92181 89153
rect 92139 89104 92140 89144
rect 92180 89104 92181 89144
rect 92139 89095 92181 89104
rect 90700 89010 90740 89095
rect 92140 89010 92180 89095
rect 78184 88472 78552 88481
rect 78224 88432 78266 88472
rect 78306 88432 78348 88472
rect 78388 88432 78430 88472
rect 78470 88432 78512 88472
rect 78184 88423 78552 88432
rect 93304 88472 93672 88481
rect 93344 88432 93386 88472
rect 93426 88432 93468 88472
rect 93508 88432 93550 88472
rect 93590 88432 93632 88472
rect 93304 88423 93672 88432
rect 108424 88472 108792 88481
rect 108464 88432 108506 88472
rect 108546 88432 108588 88472
rect 108628 88432 108670 88472
rect 108710 88432 108752 88472
rect 108424 88423 108792 88432
rect 123544 88472 123912 88481
rect 123584 88432 123626 88472
rect 123666 88432 123708 88472
rect 123748 88432 123790 88472
rect 123830 88432 123872 88472
rect 123544 88423 123912 88432
rect 138664 88472 139032 88481
rect 138704 88432 138746 88472
rect 138786 88432 138828 88472
rect 138868 88432 138910 88472
rect 138950 88432 138992 88472
rect 138664 88423 139032 88432
rect 79424 87716 79792 87725
rect 79464 87676 79506 87716
rect 79546 87676 79588 87716
rect 79628 87676 79670 87716
rect 79710 87676 79752 87716
rect 79424 87667 79792 87676
rect 94544 87716 94912 87725
rect 94584 87676 94626 87716
rect 94666 87676 94708 87716
rect 94748 87676 94790 87716
rect 94830 87676 94872 87716
rect 94544 87667 94912 87676
rect 109664 87716 110032 87725
rect 109704 87676 109746 87716
rect 109786 87676 109828 87716
rect 109868 87676 109910 87716
rect 109950 87676 109992 87716
rect 109664 87667 110032 87676
rect 124784 87716 125152 87725
rect 124824 87676 124866 87716
rect 124906 87676 124948 87716
rect 124988 87676 125030 87716
rect 125070 87676 125112 87716
rect 124784 87667 125152 87676
rect 139904 87716 140272 87725
rect 139944 87676 139986 87716
rect 140026 87676 140068 87716
rect 140108 87676 140150 87716
rect 140190 87676 140232 87716
rect 139904 87667 140272 87676
rect 78184 86960 78552 86969
rect 78224 86920 78266 86960
rect 78306 86920 78348 86960
rect 78388 86920 78430 86960
rect 78470 86920 78512 86960
rect 78184 86911 78552 86920
rect 93304 86960 93672 86969
rect 93344 86920 93386 86960
rect 93426 86920 93468 86960
rect 93508 86920 93550 86960
rect 93590 86920 93632 86960
rect 93304 86911 93672 86920
rect 108424 86960 108792 86969
rect 108464 86920 108506 86960
rect 108546 86920 108588 86960
rect 108628 86920 108670 86960
rect 108710 86920 108752 86960
rect 108424 86911 108792 86920
rect 123544 86960 123912 86969
rect 123584 86920 123626 86960
rect 123666 86920 123708 86960
rect 123748 86920 123790 86960
rect 123830 86920 123872 86960
rect 123544 86911 123912 86920
rect 138664 86960 139032 86969
rect 138704 86920 138746 86960
rect 138786 86920 138828 86960
rect 138868 86920 138910 86960
rect 138950 86920 138992 86960
rect 138664 86911 139032 86920
rect 79424 86204 79792 86213
rect 79464 86164 79506 86204
rect 79546 86164 79588 86204
rect 79628 86164 79670 86204
rect 79710 86164 79752 86204
rect 79424 86155 79792 86164
rect 94544 86204 94912 86213
rect 94584 86164 94626 86204
rect 94666 86164 94708 86204
rect 94748 86164 94790 86204
rect 94830 86164 94872 86204
rect 94544 86155 94912 86164
rect 109664 86204 110032 86213
rect 109704 86164 109746 86204
rect 109786 86164 109828 86204
rect 109868 86164 109910 86204
rect 109950 86164 109992 86204
rect 109664 86155 110032 86164
rect 124784 86204 125152 86213
rect 124824 86164 124866 86204
rect 124906 86164 124948 86204
rect 124988 86164 125030 86204
rect 125070 86164 125112 86204
rect 124784 86155 125152 86164
rect 139904 86204 140272 86213
rect 139944 86164 139986 86204
rect 140026 86164 140068 86204
rect 140108 86164 140150 86204
rect 140190 86164 140232 86204
rect 139904 86155 140272 86164
rect 78184 85448 78552 85457
rect 78224 85408 78266 85448
rect 78306 85408 78348 85448
rect 78388 85408 78430 85448
rect 78470 85408 78512 85448
rect 78184 85399 78552 85408
rect 93304 85448 93672 85457
rect 93344 85408 93386 85448
rect 93426 85408 93468 85448
rect 93508 85408 93550 85448
rect 93590 85408 93632 85448
rect 93304 85399 93672 85408
rect 108424 85448 108792 85457
rect 108464 85408 108506 85448
rect 108546 85408 108588 85448
rect 108628 85408 108670 85448
rect 108710 85408 108752 85448
rect 108424 85399 108792 85408
rect 123544 85448 123912 85457
rect 123584 85408 123626 85448
rect 123666 85408 123708 85448
rect 123748 85408 123790 85448
rect 123830 85408 123872 85448
rect 123544 85399 123912 85408
rect 138664 85448 139032 85457
rect 138704 85408 138746 85448
rect 138786 85408 138828 85448
rect 138868 85408 138910 85448
rect 138950 85408 138992 85448
rect 138664 85399 139032 85408
rect 79424 84692 79792 84701
rect 79464 84652 79506 84692
rect 79546 84652 79588 84692
rect 79628 84652 79670 84692
rect 79710 84652 79752 84692
rect 79424 84643 79792 84652
rect 94544 84692 94912 84701
rect 94584 84652 94626 84692
rect 94666 84652 94708 84692
rect 94748 84652 94790 84692
rect 94830 84652 94872 84692
rect 94544 84643 94912 84652
rect 109664 84692 110032 84701
rect 109704 84652 109746 84692
rect 109786 84652 109828 84692
rect 109868 84652 109910 84692
rect 109950 84652 109992 84692
rect 109664 84643 110032 84652
rect 124784 84692 125152 84701
rect 124824 84652 124866 84692
rect 124906 84652 124948 84692
rect 124988 84652 125030 84692
rect 125070 84652 125112 84692
rect 124784 84643 125152 84652
rect 139904 84692 140272 84701
rect 139944 84652 139986 84692
rect 140026 84652 140068 84692
rect 140108 84652 140150 84692
rect 140190 84652 140232 84692
rect 139904 84643 140272 84652
rect 78184 83936 78552 83945
rect 78224 83896 78266 83936
rect 78306 83896 78348 83936
rect 78388 83896 78430 83936
rect 78470 83896 78512 83936
rect 78184 83887 78552 83896
rect 93304 83936 93672 83945
rect 93344 83896 93386 83936
rect 93426 83896 93468 83936
rect 93508 83896 93550 83936
rect 93590 83896 93632 83936
rect 93304 83887 93672 83896
rect 108424 83936 108792 83945
rect 108464 83896 108506 83936
rect 108546 83896 108588 83936
rect 108628 83896 108670 83936
rect 108710 83896 108752 83936
rect 108424 83887 108792 83896
rect 123544 83936 123912 83945
rect 123584 83896 123626 83936
rect 123666 83896 123708 83936
rect 123748 83896 123790 83936
rect 123830 83896 123872 83936
rect 123544 83887 123912 83896
rect 138664 83936 139032 83945
rect 138704 83896 138746 83936
rect 138786 83896 138828 83936
rect 138868 83896 138910 83936
rect 138950 83896 138992 83936
rect 138664 83887 139032 83896
rect 79424 83180 79792 83189
rect 79464 83140 79506 83180
rect 79546 83140 79588 83180
rect 79628 83140 79670 83180
rect 79710 83140 79752 83180
rect 79424 83131 79792 83140
rect 94544 83180 94912 83189
rect 94584 83140 94626 83180
rect 94666 83140 94708 83180
rect 94748 83140 94790 83180
rect 94830 83140 94872 83180
rect 94544 83131 94912 83140
rect 109664 83180 110032 83189
rect 109704 83140 109746 83180
rect 109786 83140 109828 83180
rect 109868 83140 109910 83180
rect 109950 83140 109992 83180
rect 109664 83131 110032 83140
rect 124784 83180 125152 83189
rect 124824 83140 124866 83180
rect 124906 83140 124948 83180
rect 124988 83140 125030 83180
rect 125070 83140 125112 83180
rect 124784 83131 125152 83140
rect 139904 83180 140272 83189
rect 139944 83140 139986 83180
rect 140026 83140 140068 83180
rect 140108 83140 140150 83180
rect 140190 83140 140232 83180
rect 139904 83131 140272 83140
rect 78184 82424 78552 82433
rect 78224 82384 78266 82424
rect 78306 82384 78348 82424
rect 78388 82384 78430 82424
rect 78470 82384 78512 82424
rect 78184 82375 78552 82384
rect 93304 82424 93672 82433
rect 93344 82384 93386 82424
rect 93426 82384 93468 82424
rect 93508 82384 93550 82424
rect 93590 82384 93632 82424
rect 93304 82375 93672 82384
rect 108424 82424 108792 82433
rect 108464 82384 108506 82424
rect 108546 82384 108588 82424
rect 108628 82384 108670 82424
rect 108710 82384 108752 82424
rect 108424 82375 108792 82384
rect 123544 82424 123912 82433
rect 123584 82384 123626 82424
rect 123666 82384 123708 82424
rect 123748 82384 123790 82424
rect 123830 82384 123872 82424
rect 123544 82375 123912 82384
rect 138664 82424 139032 82433
rect 138704 82384 138746 82424
rect 138786 82384 138828 82424
rect 138868 82384 138910 82424
rect 138950 82384 138992 82424
rect 138664 82375 139032 82384
rect 79424 81668 79792 81677
rect 79464 81628 79506 81668
rect 79546 81628 79588 81668
rect 79628 81628 79670 81668
rect 79710 81628 79752 81668
rect 79424 81619 79792 81628
rect 94544 81668 94912 81677
rect 94584 81628 94626 81668
rect 94666 81628 94708 81668
rect 94748 81628 94790 81668
rect 94830 81628 94872 81668
rect 94544 81619 94912 81628
rect 109664 81668 110032 81677
rect 109704 81628 109746 81668
rect 109786 81628 109828 81668
rect 109868 81628 109910 81668
rect 109950 81628 109992 81668
rect 109664 81619 110032 81628
rect 124784 81668 125152 81677
rect 124824 81628 124866 81668
rect 124906 81628 124948 81668
rect 124988 81628 125030 81668
rect 125070 81628 125112 81668
rect 124784 81619 125152 81628
rect 139904 81668 140272 81677
rect 139944 81628 139986 81668
rect 140026 81628 140068 81668
rect 140108 81628 140150 81668
rect 140190 81628 140232 81668
rect 139904 81619 140272 81628
rect 78184 80912 78552 80921
rect 78224 80872 78266 80912
rect 78306 80872 78348 80912
rect 78388 80872 78430 80912
rect 78470 80872 78512 80912
rect 78184 80863 78552 80872
rect 93304 80912 93672 80921
rect 93344 80872 93386 80912
rect 93426 80872 93468 80912
rect 93508 80872 93550 80912
rect 93590 80872 93632 80912
rect 93304 80863 93672 80872
rect 108424 80912 108792 80921
rect 108464 80872 108506 80912
rect 108546 80872 108588 80912
rect 108628 80872 108670 80912
rect 108710 80872 108752 80912
rect 108424 80863 108792 80872
rect 123544 80912 123912 80921
rect 123584 80872 123626 80912
rect 123666 80872 123708 80912
rect 123748 80872 123790 80912
rect 123830 80872 123872 80912
rect 123544 80863 123912 80872
rect 138664 80912 139032 80921
rect 138704 80872 138746 80912
rect 138786 80872 138828 80912
rect 138868 80872 138910 80912
rect 138950 80872 138992 80912
rect 138664 80863 139032 80872
rect 79424 80156 79792 80165
rect 79464 80116 79506 80156
rect 79546 80116 79588 80156
rect 79628 80116 79670 80156
rect 79710 80116 79752 80156
rect 79424 80107 79792 80116
rect 94544 80156 94912 80165
rect 94584 80116 94626 80156
rect 94666 80116 94708 80156
rect 94748 80116 94790 80156
rect 94830 80116 94872 80156
rect 94544 80107 94912 80116
rect 109664 80156 110032 80165
rect 109704 80116 109746 80156
rect 109786 80116 109828 80156
rect 109868 80116 109910 80156
rect 109950 80116 109992 80156
rect 109664 80107 110032 80116
rect 124784 80156 125152 80165
rect 124824 80116 124866 80156
rect 124906 80116 124948 80156
rect 124988 80116 125030 80156
rect 125070 80116 125112 80156
rect 124784 80107 125152 80116
rect 139904 80156 140272 80165
rect 139944 80116 139986 80156
rect 140026 80116 140068 80156
rect 140108 80116 140150 80156
rect 140190 80116 140232 80156
rect 139904 80107 140272 80116
rect 78184 79400 78552 79409
rect 78224 79360 78266 79400
rect 78306 79360 78348 79400
rect 78388 79360 78430 79400
rect 78470 79360 78512 79400
rect 78184 79351 78552 79360
rect 93304 79400 93672 79409
rect 93344 79360 93386 79400
rect 93426 79360 93468 79400
rect 93508 79360 93550 79400
rect 93590 79360 93632 79400
rect 93304 79351 93672 79360
rect 108424 79400 108792 79409
rect 108464 79360 108506 79400
rect 108546 79360 108588 79400
rect 108628 79360 108670 79400
rect 108710 79360 108752 79400
rect 108424 79351 108792 79360
rect 123544 79400 123912 79409
rect 123584 79360 123626 79400
rect 123666 79360 123708 79400
rect 123748 79360 123790 79400
rect 123830 79360 123872 79400
rect 123544 79351 123912 79360
rect 138664 79400 139032 79409
rect 138704 79360 138746 79400
rect 138786 79360 138828 79400
rect 138868 79360 138910 79400
rect 138950 79360 138992 79400
rect 138664 79351 139032 79360
rect 79424 78644 79792 78653
rect 79464 78604 79506 78644
rect 79546 78604 79588 78644
rect 79628 78604 79670 78644
rect 79710 78604 79752 78644
rect 79424 78595 79792 78604
rect 94544 78644 94912 78653
rect 94584 78604 94626 78644
rect 94666 78604 94708 78644
rect 94748 78604 94790 78644
rect 94830 78604 94872 78644
rect 94544 78595 94912 78604
rect 109664 78644 110032 78653
rect 109704 78604 109746 78644
rect 109786 78604 109828 78644
rect 109868 78604 109910 78644
rect 109950 78604 109992 78644
rect 109664 78595 110032 78604
rect 124784 78644 125152 78653
rect 124824 78604 124866 78644
rect 124906 78604 124948 78644
rect 124988 78604 125030 78644
rect 125070 78604 125112 78644
rect 124784 78595 125152 78604
rect 139904 78644 140272 78653
rect 139944 78604 139986 78644
rect 140026 78604 140068 78644
rect 140108 78604 140150 78644
rect 140190 78604 140232 78644
rect 139904 78595 140272 78604
rect 78184 77888 78552 77897
rect 78224 77848 78266 77888
rect 78306 77848 78348 77888
rect 78388 77848 78430 77888
rect 78470 77848 78512 77888
rect 78184 77839 78552 77848
rect 93304 77888 93672 77897
rect 93344 77848 93386 77888
rect 93426 77848 93468 77888
rect 93508 77848 93550 77888
rect 93590 77848 93632 77888
rect 93304 77839 93672 77848
rect 108424 77888 108792 77897
rect 108464 77848 108506 77888
rect 108546 77848 108588 77888
rect 108628 77848 108670 77888
rect 108710 77848 108752 77888
rect 108424 77839 108792 77848
rect 123544 77888 123912 77897
rect 123584 77848 123626 77888
rect 123666 77848 123708 77888
rect 123748 77848 123790 77888
rect 123830 77848 123872 77888
rect 123544 77839 123912 77848
rect 138664 77888 139032 77897
rect 138704 77848 138746 77888
rect 138786 77848 138828 77888
rect 138868 77848 138910 77888
rect 138950 77848 138992 77888
rect 138664 77839 139032 77848
rect 79424 77132 79792 77141
rect 79464 77092 79506 77132
rect 79546 77092 79588 77132
rect 79628 77092 79670 77132
rect 79710 77092 79752 77132
rect 79424 77083 79792 77092
rect 94544 77132 94912 77141
rect 94584 77092 94626 77132
rect 94666 77092 94708 77132
rect 94748 77092 94790 77132
rect 94830 77092 94872 77132
rect 94544 77083 94912 77092
rect 109664 77132 110032 77141
rect 109704 77092 109746 77132
rect 109786 77092 109828 77132
rect 109868 77092 109910 77132
rect 109950 77092 109992 77132
rect 109664 77083 110032 77092
rect 124784 77132 125152 77141
rect 124824 77092 124866 77132
rect 124906 77092 124948 77132
rect 124988 77092 125030 77132
rect 125070 77092 125112 77132
rect 124784 77083 125152 77092
rect 139904 77132 140272 77141
rect 139944 77092 139986 77132
rect 140026 77092 140068 77132
rect 140108 77092 140150 77132
rect 140190 77092 140232 77132
rect 139904 77083 140272 77092
rect 78184 76376 78552 76385
rect 78224 76336 78266 76376
rect 78306 76336 78348 76376
rect 78388 76336 78430 76376
rect 78470 76336 78512 76376
rect 78184 76327 78552 76336
rect 93304 76376 93672 76385
rect 93344 76336 93386 76376
rect 93426 76336 93468 76376
rect 93508 76336 93550 76376
rect 93590 76336 93632 76376
rect 93304 76327 93672 76336
rect 108424 76376 108792 76385
rect 108464 76336 108506 76376
rect 108546 76336 108588 76376
rect 108628 76336 108670 76376
rect 108710 76336 108752 76376
rect 108424 76327 108792 76336
rect 123544 76376 123912 76385
rect 123584 76336 123626 76376
rect 123666 76336 123708 76376
rect 123748 76336 123790 76376
rect 123830 76336 123872 76376
rect 123544 76327 123912 76336
rect 138664 76376 139032 76385
rect 138704 76336 138746 76376
rect 138786 76336 138828 76376
rect 138868 76336 138910 76376
rect 138950 76336 138992 76376
rect 138664 76327 139032 76336
rect 79424 75620 79792 75629
rect 79464 75580 79506 75620
rect 79546 75580 79588 75620
rect 79628 75580 79670 75620
rect 79710 75580 79752 75620
rect 79424 75571 79792 75580
rect 94544 75620 94912 75629
rect 94584 75580 94626 75620
rect 94666 75580 94708 75620
rect 94748 75580 94790 75620
rect 94830 75580 94872 75620
rect 94544 75571 94912 75580
rect 109664 75620 110032 75629
rect 109704 75580 109746 75620
rect 109786 75580 109828 75620
rect 109868 75580 109910 75620
rect 109950 75580 109992 75620
rect 109664 75571 110032 75580
rect 124784 75620 125152 75629
rect 124824 75580 124866 75620
rect 124906 75580 124948 75620
rect 124988 75580 125030 75620
rect 125070 75580 125112 75620
rect 124784 75571 125152 75580
rect 139904 75620 140272 75629
rect 139944 75580 139986 75620
rect 140026 75580 140068 75620
rect 140108 75580 140150 75620
rect 140190 75580 140232 75620
rect 139904 75571 140272 75580
rect 90699 71252 90741 71261
rect 90699 71212 90700 71252
rect 90740 71212 90741 71252
rect 90699 71203 90741 71212
rect 92139 71252 92181 71261
rect 92139 71212 92140 71252
rect 92180 71212 92181 71252
rect 92139 71203 92181 71212
rect 90700 71118 90740 71203
rect 92140 71118 92180 71203
<< via4 >>
rect 79424 148156 79464 148196
rect 79506 148156 79546 148196
rect 79588 148156 79628 148196
rect 79670 148156 79710 148196
rect 79752 148156 79792 148196
rect 94544 148156 94584 148196
rect 94626 148156 94666 148196
rect 94708 148156 94748 148196
rect 94790 148156 94830 148196
rect 94872 148156 94912 148196
rect 109664 148156 109704 148196
rect 109746 148156 109786 148196
rect 109828 148156 109868 148196
rect 109910 148156 109950 148196
rect 109992 148156 110032 148196
rect 124784 148156 124824 148196
rect 124866 148156 124906 148196
rect 124948 148156 124988 148196
rect 125030 148156 125070 148196
rect 125112 148156 125152 148196
rect 139904 148156 139944 148196
rect 139986 148156 140026 148196
rect 140068 148156 140108 148196
rect 140150 148156 140190 148196
rect 140232 148156 140272 148196
rect 78184 147400 78224 147440
rect 78266 147400 78306 147440
rect 78348 147400 78388 147440
rect 78430 147400 78470 147440
rect 78512 147400 78552 147440
rect 93304 147400 93344 147440
rect 93386 147400 93426 147440
rect 93468 147400 93508 147440
rect 93550 147400 93590 147440
rect 93632 147400 93672 147440
rect 108424 147400 108464 147440
rect 108506 147400 108546 147440
rect 108588 147400 108628 147440
rect 108670 147400 108710 147440
rect 108752 147400 108792 147440
rect 123544 147400 123584 147440
rect 123626 147400 123666 147440
rect 123708 147400 123748 147440
rect 123790 147400 123830 147440
rect 123872 147400 123912 147440
rect 138664 147400 138704 147440
rect 138746 147400 138786 147440
rect 138828 147400 138868 147440
rect 138910 147400 138950 147440
rect 138992 147400 139032 147440
rect 79424 146644 79464 146684
rect 79506 146644 79546 146684
rect 79588 146644 79628 146684
rect 79670 146644 79710 146684
rect 79752 146644 79792 146684
rect 94544 146644 94584 146684
rect 94626 146644 94666 146684
rect 94708 146644 94748 146684
rect 94790 146644 94830 146684
rect 94872 146644 94912 146684
rect 109664 146644 109704 146684
rect 109746 146644 109786 146684
rect 109828 146644 109868 146684
rect 109910 146644 109950 146684
rect 109992 146644 110032 146684
rect 124784 146644 124824 146684
rect 124866 146644 124906 146684
rect 124948 146644 124988 146684
rect 125030 146644 125070 146684
rect 125112 146644 125152 146684
rect 139904 146644 139944 146684
rect 139986 146644 140026 146684
rect 140068 146644 140108 146684
rect 140150 146644 140190 146684
rect 140232 146644 140272 146684
rect 78184 145888 78224 145928
rect 78266 145888 78306 145928
rect 78348 145888 78388 145928
rect 78430 145888 78470 145928
rect 78512 145888 78552 145928
rect 93304 145888 93344 145928
rect 93386 145888 93426 145928
rect 93468 145888 93508 145928
rect 93550 145888 93590 145928
rect 93632 145888 93672 145928
rect 108424 145888 108464 145928
rect 108506 145888 108546 145928
rect 108588 145888 108628 145928
rect 108670 145888 108710 145928
rect 108752 145888 108792 145928
rect 123544 145888 123584 145928
rect 123626 145888 123666 145928
rect 123708 145888 123748 145928
rect 123790 145888 123830 145928
rect 123872 145888 123912 145928
rect 138664 145888 138704 145928
rect 138746 145888 138786 145928
rect 138828 145888 138868 145928
rect 138910 145888 138950 145928
rect 138992 145888 139032 145928
rect 79424 145132 79464 145172
rect 79506 145132 79546 145172
rect 79588 145132 79628 145172
rect 79670 145132 79710 145172
rect 79752 145132 79792 145172
rect 94544 145132 94584 145172
rect 94626 145132 94666 145172
rect 94708 145132 94748 145172
rect 94790 145132 94830 145172
rect 94872 145132 94912 145172
rect 109664 145132 109704 145172
rect 109746 145132 109786 145172
rect 109828 145132 109868 145172
rect 109910 145132 109950 145172
rect 109992 145132 110032 145172
rect 124784 145132 124824 145172
rect 124866 145132 124906 145172
rect 124948 145132 124988 145172
rect 125030 145132 125070 145172
rect 125112 145132 125152 145172
rect 139904 145132 139944 145172
rect 139986 145132 140026 145172
rect 140068 145132 140108 145172
rect 140150 145132 140190 145172
rect 140232 145132 140272 145172
rect 78184 144376 78224 144416
rect 78266 144376 78306 144416
rect 78348 144376 78388 144416
rect 78430 144376 78470 144416
rect 78512 144376 78552 144416
rect 93304 144376 93344 144416
rect 93386 144376 93426 144416
rect 93468 144376 93508 144416
rect 93550 144376 93590 144416
rect 93632 144376 93672 144416
rect 108424 144376 108464 144416
rect 108506 144376 108546 144416
rect 108588 144376 108628 144416
rect 108670 144376 108710 144416
rect 108752 144376 108792 144416
rect 123544 144376 123584 144416
rect 123626 144376 123666 144416
rect 123708 144376 123748 144416
rect 123790 144376 123830 144416
rect 123872 144376 123912 144416
rect 138664 144376 138704 144416
rect 138746 144376 138786 144416
rect 138828 144376 138868 144416
rect 138910 144376 138950 144416
rect 138992 144376 139032 144416
rect 79424 143620 79464 143660
rect 79506 143620 79546 143660
rect 79588 143620 79628 143660
rect 79670 143620 79710 143660
rect 79752 143620 79792 143660
rect 94544 143620 94584 143660
rect 94626 143620 94666 143660
rect 94708 143620 94748 143660
rect 94790 143620 94830 143660
rect 94872 143620 94912 143660
rect 109664 143620 109704 143660
rect 109746 143620 109786 143660
rect 109828 143620 109868 143660
rect 109910 143620 109950 143660
rect 109992 143620 110032 143660
rect 124784 143620 124824 143660
rect 124866 143620 124906 143660
rect 124948 143620 124988 143660
rect 125030 143620 125070 143660
rect 125112 143620 125152 143660
rect 139904 143620 139944 143660
rect 139986 143620 140026 143660
rect 140068 143620 140108 143660
rect 140150 143620 140190 143660
rect 140232 143620 140272 143660
rect 78184 142864 78224 142904
rect 78266 142864 78306 142904
rect 78348 142864 78388 142904
rect 78430 142864 78470 142904
rect 78512 142864 78552 142904
rect 93304 142864 93344 142904
rect 93386 142864 93426 142904
rect 93468 142864 93508 142904
rect 93550 142864 93590 142904
rect 93632 142864 93672 142904
rect 108424 142864 108464 142904
rect 108506 142864 108546 142904
rect 108588 142864 108628 142904
rect 108670 142864 108710 142904
rect 108752 142864 108792 142904
rect 123544 142864 123584 142904
rect 123626 142864 123666 142904
rect 123708 142864 123748 142904
rect 123790 142864 123830 142904
rect 123872 142864 123912 142904
rect 138664 142864 138704 142904
rect 138746 142864 138786 142904
rect 138828 142864 138868 142904
rect 138910 142864 138950 142904
rect 138992 142864 139032 142904
rect 79424 142108 79464 142148
rect 79506 142108 79546 142148
rect 79588 142108 79628 142148
rect 79670 142108 79710 142148
rect 79752 142108 79792 142148
rect 94544 142108 94584 142148
rect 94626 142108 94666 142148
rect 94708 142108 94748 142148
rect 94790 142108 94830 142148
rect 94872 142108 94912 142148
rect 109664 142108 109704 142148
rect 109746 142108 109786 142148
rect 109828 142108 109868 142148
rect 109910 142108 109950 142148
rect 109992 142108 110032 142148
rect 124784 142108 124824 142148
rect 124866 142108 124906 142148
rect 124948 142108 124988 142148
rect 125030 142108 125070 142148
rect 125112 142108 125152 142148
rect 139904 142108 139944 142148
rect 139986 142108 140026 142148
rect 140068 142108 140108 142148
rect 140150 142108 140190 142148
rect 140232 142108 140272 142148
rect 78184 141352 78224 141392
rect 78266 141352 78306 141392
rect 78348 141352 78388 141392
rect 78430 141352 78470 141392
rect 78512 141352 78552 141392
rect 93304 141352 93344 141392
rect 93386 141352 93426 141392
rect 93468 141352 93508 141392
rect 93550 141352 93590 141392
rect 93632 141352 93672 141392
rect 108424 141352 108464 141392
rect 108506 141352 108546 141392
rect 108588 141352 108628 141392
rect 108670 141352 108710 141392
rect 108752 141352 108792 141392
rect 123544 141352 123584 141392
rect 123626 141352 123666 141392
rect 123708 141352 123748 141392
rect 123790 141352 123830 141392
rect 123872 141352 123912 141392
rect 138664 141352 138704 141392
rect 138746 141352 138786 141392
rect 138828 141352 138868 141392
rect 138910 141352 138950 141392
rect 138992 141352 139032 141392
rect 79424 140596 79464 140636
rect 79506 140596 79546 140636
rect 79588 140596 79628 140636
rect 79670 140596 79710 140636
rect 79752 140596 79792 140636
rect 94544 140596 94584 140636
rect 94626 140596 94666 140636
rect 94708 140596 94748 140636
rect 94790 140596 94830 140636
rect 94872 140596 94912 140636
rect 109664 140596 109704 140636
rect 109746 140596 109786 140636
rect 109828 140596 109868 140636
rect 109910 140596 109950 140636
rect 109992 140596 110032 140636
rect 124784 140596 124824 140636
rect 124866 140596 124906 140636
rect 124948 140596 124988 140636
rect 125030 140596 125070 140636
rect 125112 140596 125152 140636
rect 139904 140596 139944 140636
rect 139986 140596 140026 140636
rect 140068 140596 140108 140636
rect 140150 140596 140190 140636
rect 140232 140596 140272 140636
rect 78184 139840 78224 139880
rect 78266 139840 78306 139880
rect 78348 139840 78388 139880
rect 78430 139840 78470 139880
rect 78512 139840 78552 139880
rect 93304 139840 93344 139880
rect 93386 139840 93426 139880
rect 93468 139840 93508 139880
rect 93550 139840 93590 139880
rect 93632 139840 93672 139880
rect 108424 139840 108464 139880
rect 108506 139840 108546 139880
rect 108588 139840 108628 139880
rect 108670 139840 108710 139880
rect 108752 139840 108792 139880
rect 123544 139840 123584 139880
rect 123626 139840 123666 139880
rect 123708 139840 123748 139880
rect 123790 139840 123830 139880
rect 123872 139840 123912 139880
rect 138664 139840 138704 139880
rect 138746 139840 138786 139880
rect 138828 139840 138868 139880
rect 138910 139840 138950 139880
rect 138992 139840 139032 139880
rect 79424 139084 79464 139124
rect 79506 139084 79546 139124
rect 79588 139084 79628 139124
rect 79670 139084 79710 139124
rect 79752 139084 79792 139124
rect 94544 139084 94584 139124
rect 94626 139084 94666 139124
rect 94708 139084 94748 139124
rect 94790 139084 94830 139124
rect 94872 139084 94912 139124
rect 109664 139084 109704 139124
rect 109746 139084 109786 139124
rect 109828 139084 109868 139124
rect 109910 139084 109950 139124
rect 109992 139084 110032 139124
rect 124784 139084 124824 139124
rect 124866 139084 124906 139124
rect 124948 139084 124988 139124
rect 125030 139084 125070 139124
rect 125112 139084 125152 139124
rect 139904 139084 139944 139124
rect 139986 139084 140026 139124
rect 140068 139084 140108 139124
rect 140150 139084 140190 139124
rect 140232 139084 140272 139124
rect 78184 138328 78224 138368
rect 78266 138328 78306 138368
rect 78348 138328 78388 138368
rect 78430 138328 78470 138368
rect 78512 138328 78552 138368
rect 93304 138328 93344 138368
rect 93386 138328 93426 138368
rect 93468 138328 93508 138368
rect 93550 138328 93590 138368
rect 93632 138328 93672 138368
rect 108424 138328 108464 138368
rect 108506 138328 108546 138368
rect 108588 138328 108628 138368
rect 108670 138328 108710 138368
rect 108752 138328 108792 138368
rect 123544 138328 123584 138368
rect 123626 138328 123666 138368
rect 123708 138328 123748 138368
rect 123790 138328 123830 138368
rect 123872 138328 123912 138368
rect 138664 138328 138704 138368
rect 138746 138328 138786 138368
rect 138828 138328 138868 138368
rect 138910 138328 138950 138368
rect 138992 138328 139032 138368
rect 79424 137572 79464 137612
rect 79506 137572 79546 137612
rect 79588 137572 79628 137612
rect 79670 137572 79710 137612
rect 79752 137572 79792 137612
rect 94544 137572 94584 137612
rect 94626 137572 94666 137612
rect 94708 137572 94748 137612
rect 94790 137572 94830 137612
rect 94872 137572 94912 137612
rect 109664 137572 109704 137612
rect 109746 137572 109786 137612
rect 109828 137572 109868 137612
rect 109910 137572 109950 137612
rect 109992 137572 110032 137612
rect 124784 137572 124824 137612
rect 124866 137572 124906 137612
rect 124948 137572 124988 137612
rect 125030 137572 125070 137612
rect 125112 137572 125152 137612
rect 139904 137572 139944 137612
rect 139986 137572 140026 137612
rect 140068 137572 140108 137612
rect 140150 137572 140190 137612
rect 140232 137572 140272 137612
rect 78184 136816 78224 136856
rect 78266 136816 78306 136856
rect 78348 136816 78388 136856
rect 78430 136816 78470 136856
rect 78512 136816 78552 136856
rect 93304 136816 93344 136856
rect 93386 136816 93426 136856
rect 93468 136816 93508 136856
rect 93550 136816 93590 136856
rect 93632 136816 93672 136856
rect 108424 136816 108464 136856
rect 108506 136816 108546 136856
rect 108588 136816 108628 136856
rect 108670 136816 108710 136856
rect 108752 136816 108792 136856
rect 123544 136816 123584 136856
rect 123626 136816 123666 136856
rect 123708 136816 123748 136856
rect 123790 136816 123830 136856
rect 123872 136816 123912 136856
rect 138664 136816 138704 136856
rect 138746 136816 138786 136856
rect 138828 136816 138868 136856
rect 138910 136816 138950 136856
rect 138992 136816 139032 136856
rect 79424 136060 79464 136100
rect 79506 136060 79546 136100
rect 79588 136060 79628 136100
rect 79670 136060 79710 136100
rect 79752 136060 79792 136100
rect 94544 136060 94584 136100
rect 94626 136060 94666 136100
rect 94708 136060 94748 136100
rect 94790 136060 94830 136100
rect 94872 136060 94912 136100
rect 109664 136060 109704 136100
rect 109746 136060 109786 136100
rect 109828 136060 109868 136100
rect 109910 136060 109950 136100
rect 109992 136060 110032 136100
rect 124784 136060 124824 136100
rect 124866 136060 124906 136100
rect 124948 136060 124988 136100
rect 125030 136060 125070 136100
rect 125112 136060 125152 136100
rect 139904 136060 139944 136100
rect 139986 136060 140026 136100
rect 140068 136060 140108 136100
rect 140150 136060 140190 136100
rect 140232 136060 140272 136100
rect 78184 135304 78224 135344
rect 78266 135304 78306 135344
rect 78348 135304 78388 135344
rect 78430 135304 78470 135344
rect 78512 135304 78552 135344
rect 93304 135304 93344 135344
rect 93386 135304 93426 135344
rect 93468 135304 93508 135344
rect 93550 135304 93590 135344
rect 93632 135304 93672 135344
rect 108424 135304 108464 135344
rect 108506 135304 108546 135344
rect 108588 135304 108628 135344
rect 108670 135304 108710 135344
rect 108752 135304 108792 135344
rect 123544 135304 123584 135344
rect 123626 135304 123666 135344
rect 123708 135304 123748 135344
rect 123790 135304 123830 135344
rect 123872 135304 123912 135344
rect 138664 135304 138704 135344
rect 138746 135304 138786 135344
rect 138828 135304 138868 135344
rect 138910 135304 138950 135344
rect 138992 135304 139032 135344
rect 79424 134548 79464 134588
rect 79506 134548 79546 134588
rect 79588 134548 79628 134588
rect 79670 134548 79710 134588
rect 79752 134548 79792 134588
rect 94544 134548 94584 134588
rect 94626 134548 94666 134588
rect 94708 134548 94748 134588
rect 94790 134548 94830 134588
rect 94872 134548 94912 134588
rect 109664 134548 109704 134588
rect 109746 134548 109786 134588
rect 109828 134548 109868 134588
rect 109910 134548 109950 134588
rect 109992 134548 110032 134588
rect 124784 134548 124824 134588
rect 124866 134548 124906 134588
rect 124948 134548 124988 134588
rect 125030 134548 125070 134588
rect 125112 134548 125152 134588
rect 139904 134548 139944 134588
rect 139986 134548 140026 134588
rect 140068 134548 140108 134588
rect 140150 134548 140190 134588
rect 140232 134548 140272 134588
rect 78184 133792 78224 133832
rect 78266 133792 78306 133832
rect 78348 133792 78388 133832
rect 78430 133792 78470 133832
rect 78512 133792 78552 133832
rect 93304 133792 93344 133832
rect 93386 133792 93426 133832
rect 93468 133792 93508 133832
rect 93550 133792 93590 133832
rect 93632 133792 93672 133832
rect 108424 133792 108464 133832
rect 108506 133792 108546 133832
rect 108588 133792 108628 133832
rect 108670 133792 108710 133832
rect 108752 133792 108792 133832
rect 123544 133792 123584 133832
rect 123626 133792 123666 133832
rect 123708 133792 123748 133832
rect 123790 133792 123830 133832
rect 123872 133792 123912 133832
rect 138664 133792 138704 133832
rect 138746 133792 138786 133832
rect 138828 133792 138868 133832
rect 138910 133792 138950 133832
rect 138992 133792 139032 133832
rect 79424 133036 79464 133076
rect 79506 133036 79546 133076
rect 79588 133036 79628 133076
rect 79670 133036 79710 133076
rect 79752 133036 79792 133076
rect 94544 133036 94584 133076
rect 94626 133036 94666 133076
rect 94708 133036 94748 133076
rect 94790 133036 94830 133076
rect 94872 133036 94912 133076
rect 109664 133036 109704 133076
rect 109746 133036 109786 133076
rect 109828 133036 109868 133076
rect 109910 133036 109950 133076
rect 109992 133036 110032 133076
rect 124784 133036 124824 133076
rect 124866 133036 124906 133076
rect 124948 133036 124988 133076
rect 125030 133036 125070 133076
rect 125112 133036 125152 133076
rect 139904 133036 139944 133076
rect 139986 133036 140026 133076
rect 140068 133036 140108 133076
rect 140150 133036 140190 133076
rect 140232 133036 140272 133076
rect 78184 132280 78224 132320
rect 78266 132280 78306 132320
rect 78348 132280 78388 132320
rect 78430 132280 78470 132320
rect 78512 132280 78552 132320
rect 93304 132280 93344 132320
rect 93386 132280 93426 132320
rect 93468 132280 93508 132320
rect 93550 132280 93590 132320
rect 93632 132280 93672 132320
rect 108424 132280 108464 132320
rect 108506 132280 108546 132320
rect 108588 132280 108628 132320
rect 108670 132280 108710 132320
rect 108752 132280 108792 132320
rect 123544 132280 123584 132320
rect 123626 132280 123666 132320
rect 123708 132280 123748 132320
rect 123790 132280 123830 132320
rect 123872 132280 123912 132320
rect 138664 132280 138704 132320
rect 138746 132280 138786 132320
rect 138828 132280 138868 132320
rect 138910 132280 138950 132320
rect 138992 132280 139032 132320
rect 79424 131524 79464 131564
rect 79506 131524 79546 131564
rect 79588 131524 79628 131564
rect 79670 131524 79710 131564
rect 79752 131524 79792 131564
rect 94544 131524 94584 131564
rect 94626 131524 94666 131564
rect 94708 131524 94748 131564
rect 94790 131524 94830 131564
rect 94872 131524 94912 131564
rect 109664 131524 109704 131564
rect 109746 131524 109786 131564
rect 109828 131524 109868 131564
rect 109910 131524 109950 131564
rect 109992 131524 110032 131564
rect 124784 131524 124824 131564
rect 124866 131524 124906 131564
rect 124948 131524 124988 131564
rect 125030 131524 125070 131564
rect 125112 131524 125152 131564
rect 139904 131524 139944 131564
rect 139986 131524 140026 131564
rect 140068 131524 140108 131564
rect 140150 131524 140190 131564
rect 140232 131524 140272 131564
rect 78184 130768 78224 130808
rect 78266 130768 78306 130808
rect 78348 130768 78388 130808
rect 78430 130768 78470 130808
rect 78512 130768 78552 130808
rect 93304 130768 93344 130808
rect 93386 130768 93426 130808
rect 93468 130768 93508 130808
rect 93550 130768 93590 130808
rect 93632 130768 93672 130808
rect 108424 130768 108464 130808
rect 108506 130768 108546 130808
rect 108588 130768 108628 130808
rect 108670 130768 108710 130808
rect 108752 130768 108792 130808
rect 123544 130768 123584 130808
rect 123626 130768 123666 130808
rect 123708 130768 123748 130808
rect 123790 130768 123830 130808
rect 123872 130768 123912 130808
rect 138664 130768 138704 130808
rect 138746 130768 138786 130808
rect 138828 130768 138868 130808
rect 138910 130768 138950 130808
rect 138992 130768 139032 130808
rect 79424 130012 79464 130052
rect 79506 130012 79546 130052
rect 79588 130012 79628 130052
rect 79670 130012 79710 130052
rect 79752 130012 79792 130052
rect 94544 130012 94584 130052
rect 94626 130012 94666 130052
rect 94708 130012 94748 130052
rect 94790 130012 94830 130052
rect 94872 130012 94912 130052
rect 109664 130012 109704 130052
rect 109746 130012 109786 130052
rect 109828 130012 109868 130052
rect 109910 130012 109950 130052
rect 109992 130012 110032 130052
rect 124784 130012 124824 130052
rect 124866 130012 124906 130052
rect 124948 130012 124988 130052
rect 125030 130012 125070 130052
rect 125112 130012 125152 130052
rect 139904 130012 139944 130052
rect 139986 130012 140026 130052
rect 140068 130012 140108 130052
rect 140150 130012 140190 130052
rect 140232 130012 140272 130052
rect 78184 129256 78224 129296
rect 78266 129256 78306 129296
rect 78348 129256 78388 129296
rect 78430 129256 78470 129296
rect 78512 129256 78552 129296
rect 93304 129256 93344 129296
rect 93386 129256 93426 129296
rect 93468 129256 93508 129296
rect 93550 129256 93590 129296
rect 93632 129256 93672 129296
rect 108424 129256 108464 129296
rect 108506 129256 108546 129296
rect 108588 129256 108628 129296
rect 108670 129256 108710 129296
rect 108752 129256 108792 129296
rect 123544 129256 123584 129296
rect 123626 129256 123666 129296
rect 123708 129256 123748 129296
rect 123790 129256 123830 129296
rect 123872 129256 123912 129296
rect 138664 129256 138704 129296
rect 138746 129256 138786 129296
rect 138828 129256 138868 129296
rect 138910 129256 138950 129296
rect 138992 129256 139032 129296
rect 79424 128500 79464 128540
rect 79506 128500 79546 128540
rect 79588 128500 79628 128540
rect 79670 128500 79710 128540
rect 79752 128500 79792 128540
rect 94544 128500 94584 128540
rect 94626 128500 94666 128540
rect 94708 128500 94748 128540
rect 94790 128500 94830 128540
rect 94872 128500 94912 128540
rect 109664 128500 109704 128540
rect 109746 128500 109786 128540
rect 109828 128500 109868 128540
rect 109910 128500 109950 128540
rect 109992 128500 110032 128540
rect 124784 128500 124824 128540
rect 124866 128500 124906 128540
rect 124948 128500 124988 128540
rect 125030 128500 125070 128540
rect 125112 128500 125152 128540
rect 139904 128500 139944 128540
rect 139986 128500 140026 128540
rect 140068 128500 140108 128540
rect 140150 128500 140190 128540
rect 140232 128500 140272 128540
rect 78184 127744 78224 127784
rect 78266 127744 78306 127784
rect 78348 127744 78388 127784
rect 78430 127744 78470 127784
rect 78512 127744 78552 127784
rect 93304 127744 93344 127784
rect 93386 127744 93426 127784
rect 93468 127744 93508 127784
rect 93550 127744 93590 127784
rect 93632 127744 93672 127784
rect 108424 127744 108464 127784
rect 108506 127744 108546 127784
rect 108588 127744 108628 127784
rect 108670 127744 108710 127784
rect 108752 127744 108792 127784
rect 123544 127744 123584 127784
rect 123626 127744 123666 127784
rect 123708 127744 123748 127784
rect 123790 127744 123830 127784
rect 123872 127744 123912 127784
rect 138664 127744 138704 127784
rect 138746 127744 138786 127784
rect 138828 127744 138868 127784
rect 138910 127744 138950 127784
rect 138992 127744 139032 127784
rect 79424 126988 79464 127028
rect 79506 126988 79546 127028
rect 79588 126988 79628 127028
rect 79670 126988 79710 127028
rect 79752 126988 79792 127028
rect 94544 126988 94584 127028
rect 94626 126988 94666 127028
rect 94708 126988 94748 127028
rect 94790 126988 94830 127028
rect 94872 126988 94912 127028
rect 109664 126988 109704 127028
rect 109746 126988 109786 127028
rect 109828 126988 109868 127028
rect 109910 126988 109950 127028
rect 109992 126988 110032 127028
rect 124784 126988 124824 127028
rect 124866 126988 124906 127028
rect 124948 126988 124988 127028
rect 125030 126988 125070 127028
rect 125112 126988 125152 127028
rect 139904 126988 139944 127028
rect 139986 126988 140026 127028
rect 140068 126988 140108 127028
rect 140150 126988 140190 127028
rect 140232 126988 140272 127028
rect 78184 126232 78224 126272
rect 78266 126232 78306 126272
rect 78348 126232 78388 126272
rect 78430 126232 78470 126272
rect 78512 126232 78552 126272
rect 93304 126232 93344 126272
rect 93386 126232 93426 126272
rect 93468 126232 93508 126272
rect 93550 126232 93590 126272
rect 93632 126232 93672 126272
rect 108424 126232 108464 126272
rect 108506 126232 108546 126272
rect 108588 126232 108628 126272
rect 108670 126232 108710 126272
rect 108752 126232 108792 126272
rect 123544 126232 123584 126272
rect 123626 126232 123666 126272
rect 123708 126232 123748 126272
rect 123790 126232 123830 126272
rect 123872 126232 123912 126272
rect 138664 126232 138704 126272
rect 138746 126232 138786 126272
rect 138828 126232 138868 126272
rect 138910 126232 138950 126272
rect 138992 126232 139032 126272
rect 79424 125476 79464 125516
rect 79506 125476 79546 125516
rect 79588 125476 79628 125516
rect 79670 125476 79710 125516
rect 79752 125476 79792 125516
rect 94544 125476 94584 125516
rect 94626 125476 94666 125516
rect 94708 125476 94748 125516
rect 94790 125476 94830 125516
rect 94872 125476 94912 125516
rect 109664 125476 109704 125516
rect 109746 125476 109786 125516
rect 109828 125476 109868 125516
rect 109910 125476 109950 125516
rect 109992 125476 110032 125516
rect 124784 125476 124824 125516
rect 124866 125476 124906 125516
rect 124948 125476 124988 125516
rect 125030 125476 125070 125516
rect 125112 125476 125152 125516
rect 139904 125476 139944 125516
rect 139986 125476 140026 125516
rect 140068 125476 140108 125516
rect 140150 125476 140190 125516
rect 140232 125476 140272 125516
rect 78184 124720 78224 124760
rect 78266 124720 78306 124760
rect 78348 124720 78388 124760
rect 78430 124720 78470 124760
rect 78512 124720 78552 124760
rect 93304 124720 93344 124760
rect 93386 124720 93426 124760
rect 93468 124720 93508 124760
rect 93550 124720 93590 124760
rect 93632 124720 93672 124760
rect 79424 123964 79464 124004
rect 79506 123964 79546 124004
rect 79588 123964 79628 124004
rect 79670 123964 79710 124004
rect 79752 123964 79792 124004
rect 78184 123208 78224 123248
rect 78266 123208 78306 123248
rect 78348 123208 78388 123248
rect 78430 123208 78470 123248
rect 78512 123208 78552 123248
rect 93304 123208 93344 123248
rect 93386 123208 93426 123248
rect 93468 123208 93508 123248
rect 93550 123208 93590 123248
rect 93632 123208 93672 123248
rect 79424 122452 79464 122492
rect 79506 122452 79546 122492
rect 79588 122452 79628 122492
rect 79670 122452 79710 122492
rect 79752 122452 79792 122492
rect 108424 124720 108464 124760
rect 108506 124720 108546 124760
rect 108588 124720 108628 124760
rect 108670 124720 108710 124760
rect 108752 124720 108792 124760
rect 123544 124720 123584 124760
rect 123626 124720 123666 124760
rect 123708 124720 123748 124760
rect 123790 124720 123830 124760
rect 123872 124720 123912 124760
rect 138664 124720 138704 124760
rect 138746 124720 138786 124760
rect 138828 124720 138868 124760
rect 138910 124720 138950 124760
rect 138992 124720 139032 124760
rect 94544 123964 94584 124004
rect 94626 123964 94666 124004
rect 94708 123964 94748 124004
rect 94790 123964 94830 124004
rect 94872 123964 94912 124004
rect 109664 123964 109704 124004
rect 109746 123964 109786 124004
rect 109828 123964 109868 124004
rect 109910 123964 109950 124004
rect 109992 123964 110032 124004
rect 124784 123964 124824 124004
rect 124866 123964 124906 124004
rect 124948 123964 124988 124004
rect 125030 123964 125070 124004
rect 125112 123964 125152 124004
rect 139904 123964 139944 124004
rect 139986 123964 140026 124004
rect 140068 123964 140108 124004
rect 140150 123964 140190 124004
rect 140232 123964 140272 124004
rect 108424 123208 108464 123248
rect 108506 123208 108546 123248
rect 108588 123208 108628 123248
rect 108670 123208 108710 123248
rect 108752 123208 108792 123248
rect 123544 123208 123584 123248
rect 123626 123208 123666 123248
rect 123708 123208 123748 123248
rect 123790 123208 123830 123248
rect 123872 123208 123912 123248
rect 138664 123208 138704 123248
rect 138746 123208 138786 123248
rect 138828 123208 138868 123248
rect 138910 123208 138950 123248
rect 138992 123208 139032 123248
rect 94544 122452 94584 122492
rect 94626 122452 94666 122492
rect 94708 122452 94748 122492
rect 94790 122452 94830 122492
rect 94872 122452 94912 122492
rect 109664 122452 109704 122492
rect 109746 122452 109786 122492
rect 109828 122452 109868 122492
rect 109910 122452 109950 122492
rect 109992 122452 110032 122492
rect 124784 122452 124824 122492
rect 124866 122452 124906 122492
rect 124948 122452 124988 122492
rect 125030 122452 125070 122492
rect 125112 122452 125152 122492
rect 139904 122452 139944 122492
rect 139986 122452 140026 122492
rect 140068 122452 140108 122492
rect 140150 122452 140190 122492
rect 140232 122452 140272 122492
rect 78184 121696 78224 121736
rect 78266 121696 78306 121736
rect 78348 121696 78388 121736
rect 78430 121696 78470 121736
rect 78512 121696 78552 121736
rect 93304 121696 93344 121736
rect 93386 121696 93426 121736
rect 93468 121696 93508 121736
rect 93550 121696 93590 121736
rect 93632 121696 93672 121736
rect 108424 121696 108464 121736
rect 108506 121696 108546 121736
rect 108588 121696 108628 121736
rect 108670 121696 108710 121736
rect 108752 121696 108792 121736
rect 123544 121696 123584 121736
rect 123626 121696 123666 121736
rect 123708 121696 123748 121736
rect 123790 121696 123830 121736
rect 123872 121696 123912 121736
rect 138664 121696 138704 121736
rect 138746 121696 138786 121736
rect 138828 121696 138868 121736
rect 138910 121696 138950 121736
rect 138992 121696 139032 121736
rect 79424 120940 79464 120980
rect 79506 120940 79546 120980
rect 79588 120940 79628 120980
rect 79670 120940 79710 120980
rect 79752 120940 79792 120980
rect 94544 120940 94584 120980
rect 94626 120940 94666 120980
rect 94708 120940 94748 120980
rect 94790 120940 94830 120980
rect 94872 120940 94912 120980
rect 109664 120940 109704 120980
rect 109746 120940 109786 120980
rect 109828 120940 109868 120980
rect 109910 120940 109950 120980
rect 109992 120940 110032 120980
rect 124784 120940 124824 120980
rect 124866 120940 124906 120980
rect 124948 120940 124988 120980
rect 125030 120940 125070 120980
rect 125112 120940 125152 120980
rect 139904 120940 139944 120980
rect 139986 120940 140026 120980
rect 140068 120940 140108 120980
rect 140150 120940 140190 120980
rect 140232 120940 140272 120980
rect 78184 120184 78224 120224
rect 78266 120184 78306 120224
rect 78348 120184 78388 120224
rect 78430 120184 78470 120224
rect 78512 120184 78552 120224
rect 93304 120184 93344 120224
rect 93386 120184 93426 120224
rect 93468 120184 93508 120224
rect 93550 120184 93590 120224
rect 93632 120184 93672 120224
rect 108424 120184 108464 120224
rect 108506 120184 108546 120224
rect 108588 120184 108628 120224
rect 108670 120184 108710 120224
rect 108752 120184 108792 120224
rect 123544 120184 123584 120224
rect 123626 120184 123666 120224
rect 123708 120184 123748 120224
rect 123790 120184 123830 120224
rect 123872 120184 123912 120224
rect 138664 120184 138704 120224
rect 138746 120184 138786 120224
rect 138828 120184 138868 120224
rect 138910 120184 138950 120224
rect 138992 120184 139032 120224
rect 79424 119428 79464 119468
rect 79506 119428 79546 119468
rect 79588 119428 79628 119468
rect 79670 119428 79710 119468
rect 79752 119428 79792 119468
rect 94544 119428 94584 119468
rect 94626 119428 94666 119468
rect 94708 119428 94748 119468
rect 94790 119428 94830 119468
rect 94872 119428 94912 119468
rect 109664 119428 109704 119468
rect 109746 119428 109786 119468
rect 109828 119428 109868 119468
rect 109910 119428 109950 119468
rect 109992 119428 110032 119468
rect 124784 119428 124824 119468
rect 124866 119428 124906 119468
rect 124948 119428 124988 119468
rect 125030 119428 125070 119468
rect 125112 119428 125152 119468
rect 139904 119428 139944 119468
rect 139986 119428 140026 119468
rect 140068 119428 140108 119468
rect 140150 119428 140190 119468
rect 140232 119428 140272 119468
rect 78184 118672 78224 118712
rect 78266 118672 78306 118712
rect 78348 118672 78388 118712
rect 78430 118672 78470 118712
rect 78512 118672 78552 118712
rect 93304 118672 93344 118712
rect 93386 118672 93426 118712
rect 93468 118672 93508 118712
rect 93550 118672 93590 118712
rect 93632 118672 93672 118712
rect 108424 118672 108464 118712
rect 108506 118672 108546 118712
rect 108588 118672 108628 118712
rect 108670 118672 108710 118712
rect 108752 118672 108792 118712
rect 123544 118672 123584 118712
rect 123626 118672 123666 118712
rect 123708 118672 123748 118712
rect 123790 118672 123830 118712
rect 123872 118672 123912 118712
rect 138664 118672 138704 118712
rect 138746 118672 138786 118712
rect 138828 118672 138868 118712
rect 138910 118672 138950 118712
rect 138992 118672 139032 118712
rect 79424 117916 79464 117956
rect 79506 117916 79546 117956
rect 79588 117916 79628 117956
rect 79670 117916 79710 117956
rect 79752 117916 79792 117956
rect 94544 117916 94584 117956
rect 94626 117916 94666 117956
rect 94708 117916 94748 117956
rect 94790 117916 94830 117956
rect 94872 117916 94912 117956
rect 109664 117916 109704 117956
rect 109746 117916 109786 117956
rect 109828 117916 109868 117956
rect 109910 117916 109950 117956
rect 109992 117916 110032 117956
rect 124784 117916 124824 117956
rect 124866 117916 124906 117956
rect 124948 117916 124988 117956
rect 125030 117916 125070 117956
rect 125112 117916 125152 117956
rect 139904 117916 139944 117956
rect 139986 117916 140026 117956
rect 140068 117916 140108 117956
rect 140150 117916 140190 117956
rect 140232 117916 140272 117956
rect 78184 117160 78224 117200
rect 78266 117160 78306 117200
rect 78348 117160 78388 117200
rect 78430 117160 78470 117200
rect 78512 117160 78552 117200
rect 93304 117160 93344 117200
rect 93386 117160 93426 117200
rect 93468 117160 93508 117200
rect 93550 117160 93590 117200
rect 93632 117160 93672 117200
rect 108424 117160 108464 117200
rect 108506 117160 108546 117200
rect 108588 117160 108628 117200
rect 108670 117160 108710 117200
rect 108752 117160 108792 117200
rect 123544 117160 123584 117200
rect 123626 117160 123666 117200
rect 123708 117160 123748 117200
rect 123790 117160 123830 117200
rect 123872 117160 123912 117200
rect 138664 117160 138704 117200
rect 138746 117160 138786 117200
rect 138828 117160 138868 117200
rect 138910 117160 138950 117200
rect 138992 117160 139032 117200
rect 79424 116404 79464 116444
rect 79506 116404 79546 116444
rect 79588 116404 79628 116444
rect 79670 116404 79710 116444
rect 79752 116404 79792 116444
rect 94544 116404 94584 116444
rect 94626 116404 94666 116444
rect 94708 116404 94748 116444
rect 94790 116404 94830 116444
rect 94872 116404 94912 116444
rect 109664 116404 109704 116444
rect 109746 116404 109786 116444
rect 109828 116404 109868 116444
rect 109910 116404 109950 116444
rect 109992 116404 110032 116444
rect 124784 116404 124824 116444
rect 124866 116404 124906 116444
rect 124948 116404 124988 116444
rect 125030 116404 125070 116444
rect 125112 116404 125152 116444
rect 139904 116404 139944 116444
rect 139986 116404 140026 116444
rect 140068 116404 140108 116444
rect 140150 116404 140190 116444
rect 140232 116404 140272 116444
rect 78184 115648 78224 115688
rect 78266 115648 78306 115688
rect 78348 115648 78388 115688
rect 78430 115648 78470 115688
rect 78512 115648 78552 115688
rect 93304 115648 93344 115688
rect 93386 115648 93426 115688
rect 93468 115648 93508 115688
rect 93550 115648 93590 115688
rect 93632 115648 93672 115688
rect 108424 115648 108464 115688
rect 108506 115648 108546 115688
rect 108588 115648 108628 115688
rect 108670 115648 108710 115688
rect 108752 115648 108792 115688
rect 123544 115648 123584 115688
rect 123626 115648 123666 115688
rect 123708 115648 123748 115688
rect 123790 115648 123830 115688
rect 123872 115648 123912 115688
rect 138664 115648 138704 115688
rect 138746 115648 138786 115688
rect 138828 115648 138868 115688
rect 138910 115648 138950 115688
rect 138992 115648 139032 115688
rect 79424 114892 79464 114932
rect 79506 114892 79546 114932
rect 79588 114892 79628 114932
rect 79670 114892 79710 114932
rect 79752 114892 79792 114932
rect 94544 114892 94584 114932
rect 94626 114892 94666 114932
rect 94708 114892 94748 114932
rect 94790 114892 94830 114932
rect 94872 114892 94912 114932
rect 109664 114892 109704 114932
rect 109746 114892 109786 114932
rect 109828 114892 109868 114932
rect 109910 114892 109950 114932
rect 109992 114892 110032 114932
rect 124784 114892 124824 114932
rect 124866 114892 124906 114932
rect 124948 114892 124988 114932
rect 125030 114892 125070 114932
rect 125112 114892 125152 114932
rect 139904 114892 139944 114932
rect 139986 114892 140026 114932
rect 140068 114892 140108 114932
rect 140150 114892 140190 114932
rect 140232 114892 140272 114932
rect 78184 114136 78224 114176
rect 78266 114136 78306 114176
rect 78348 114136 78388 114176
rect 78430 114136 78470 114176
rect 78512 114136 78552 114176
rect 93304 114136 93344 114176
rect 93386 114136 93426 114176
rect 93468 114136 93508 114176
rect 93550 114136 93590 114176
rect 93632 114136 93672 114176
rect 108424 114136 108464 114176
rect 108506 114136 108546 114176
rect 108588 114136 108628 114176
rect 108670 114136 108710 114176
rect 108752 114136 108792 114176
rect 123544 114136 123584 114176
rect 123626 114136 123666 114176
rect 123708 114136 123748 114176
rect 123790 114136 123830 114176
rect 123872 114136 123912 114176
rect 138664 114136 138704 114176
rect 138746 114136 138786 114176
rect 138828 114136 138868 114176
rect 138910 114136 138950 114176
rect 138992 114136 139032 114176
rect 79424 113380 79464 113420
rect 79506 113380 79546 113420
rect 79588 113380 79628 113420
rect 79670 113380 79710 113420
rect 79752 113380 79792 113420
rect 94544 113380 94584 113420
rect 94626 113380 94666 113420
rect 94708 113380 94748 113420
rect 94790 113380 94830 113420
rect 94872 113380 94912 113420
rect 109664 113380 109704 113420
rect 109746 113380 109786 113420
rect 109828 113380 109868 113420
rect 109910 113380 109950 113420
rect 109992 113380 110032 113420
rect 124784 113380 124824 113420
rect 124866 113380 124906 113420
rect 124948 113380 124988 113420
rect 125030 113380 125070 113420
rect 125112 113380 125152 113420
rect 139904 113380 139944 113420
rect 139986 113380 140026 113420
rect 140068 113380 140108 113420
rect 140150 113380 140190 113420
rect 140232 113380 140272 113420
rect 78184 112624 78224 112664
rect 78266 112624 78306 112664
rect 78348 112624 78388 112664
rect 78430 112624 78470 112664
rect 78512 112624 78552 112664
rect 93304 112624 93344 112664
rect 93386 112624 93426 112664
rect 93468 112624 93508 112664
rect 93550 112624 93590 112664
rect 93632 112624 93672 112664
rect 108424 112624 108464 112664
rect 108506 112624 108546 112664
rect 108588 112624 108628 112664
rect 108670 112624 108710 112664
rect 108752 112624 108792 112664
rect 123544 112624 123584 112664
rect 123626 112624 123666 112664
rect 123708 112624 123748 112664
rect 123790 112624 123830 112664
rect 123872 112624 123912 112664
rect 138664 112624 138704 112664
rect 138746 112624 138786 112664
rect 138828 112624 138868 112664
rect 138910 112624 138950 112664
rect 138992 112624 139032 112664
rect 79424 111868 79464 111908
rect 79506 111868 79546 111908
rect 79588 111868 79628 111908
rect 79670 111868 79710 111908
rect 79752 111868 79792 111908
rect 94544 111868 94584 111908
rect 94626 111868 94666 111908
rect 94708 111868 94748 111908
rect 94790 111868 94830 111908
rect 94872 111868 94912 111908
rect 109664 111868 109704 111908
rect 109746 111868 109786 111908
rect 109828 111868 109868 111908
rect 109910 111868 109950 111908
rect 109992 111868 110032 111908
rect 124784 111868 124824 111908
rect 124866 111868 124906 111908
rect 124948 111868 124988 111908
rect 125030 111868 125070 111908
rect 125112 111868 125152 111908
rect 139904 111868 139944 111908
rect 139986 111868 140026 111908
rect 140068 111868 140108 111908
rect 140150 111868 140190 111908
rect 140232 111868 140272 111908
rect 78184 111112 78224 111152
rect 78266 111112 78306 111152
rect 78348 111112 78388 111152
rect 78430 111112 78470 111152
rect 78512 111112 78552 111152
rect 93304 111112 93344 111152
rect 93386 111112 93426 111152
rect 93468 111112 93508 111152
rect 93550 111112 93590 111152
rect 93632 111112 93672 111152
rect 108424 111112 108464 111152
rect 108506 111112 108546 111152
rect 108588 111112 108628 111152
rect 108670 111112 108710 111152
rect 108752 111112 108792 111152
rect 123544 111112 123584 111152
rect 123626 111112 123666 111152
rect 123708 111112 123748 111152
rect 123790 111112 123830 111152
rect 123872 111112 123912 111152
rect 138664 111112 138704 111152
rect 138746 111112 138786 111152
rect 138828 111112 138868 111152
rect 138910 111112 138950 111152
rect 138992 111112 139032 111152
rect 79424 110356 79464 110396
rect 79506 110356 79546 110396
rect 79588 110356 79628 110396
rect 79670 110356 79710 110396
rect 79752 110356 79792 110396
rect 94544 110356 94584 110396
rect 94626 110356 94666 110396
rect 94708 110356 94748 110396
rect 94790 110356 94830 110396
rect 94872 110356 94912 110396
rect 109664 110356 109704 110396
rect 109746 110356 109786 110396
rect 109828 110356 109868 110396
rect 109910 110356 109950 110396
rect 109992 110356 110032 110396
rect 124784 110356 124824 110396
rect 124866 110356 124906 110396
rect 124948 110356 124988 110396
rect 125030 110356 125070 110396
rect 125112 110356 125152 110396
rect 139904 110356 139944 110396
rect 139986 110356 140026 110396
rect 140068 110356 140108 110396
rect 140150 110356 140190 110396
rect 140232 110356 140272 110396
rect 78184 109600 78224 109640
rect 78266 109600 78306 109640
rect 78348 109600 78388 109640
rect 78430 109600 78470 109640
rect 78512 109600 78552 109640
rect 93304 109600 93344 109640
rect 93386 109600 93426 109640
rect 93468 109600 93508 109640
rect 93550 109600 93590 109640
rect 93632 109600 93672 109640
rect 108424 109600 108464 109640
rect 108506 109600 108546 109640
rect 108588 109600 108628 109640
rect 108670 109600 108710 109640
rect 108752 109600 108792 109640
rect 123544 109600 123584 109640
rect 123626 109600 123666 109640
rect 123708 109600 123748 109640
rect 123790 109600 123830 109640
rect 123872 109600 123912 109640
rect 138664 109600 138704 109640
rect 138746 109600 138786 109640
rect 138828 109600 138868 109640
rect 138910 109600 138950 109640
rect 138992 109600 139032 109640
rect 79424 108844 79464 108884
rect 79506 108844 79546 108884
rect 79588 108844 79628 108884
rect 79670 108844 79710 108884
rect 79752 108844 79792 108884
rect 94544 108844 94584 108884
rect 94626 108844 94666 108884
rect 94708 108844 94748 108884
rect 94790 108844 94830 108884
rect 94872 108844 94912 108884
rect 109664 108844 109704 108884
rect 109746 108844 109786 108884
rect 109828 108844 109868 108884
rect 109910 108844 109950 108884
rect 109992 108844 110032 108884
rect 124784 108844 124824 108884
rect 124866 108844 124906 108884
rect 124948 108844 124988 108884
rect 125030 108844 125070 108884
rect 125112 108844 125152 108884
rect 139904 108844 139944 108884
rect 139986 108844 140026 108884
rect 140068 108844 140108 108884
rect 140150 108844 140190 108884
rect 140232 108844 140272 108884
rect 78184 108088 78224 108128
rect 78266 108088 78306 108128
rect 78348 108088 78388 108128
rect 78430 108088 78470 108128
rect 78512 108088 78552 108128
rect 93304 108088 93344 108128
rect 93386 108088 93426 108128
rect 93468 108088 93508 108128
rect 93550 108088 93590 108128
rect 93632 108088 93672 108128
rect 108424 108088 108464 108128
rect 108506 108088 108546 108128
rect 108588 108088 108628 108128
rect 108670 108088 108710 108128
rect 108752 108088 108792 108128
rect 123544 108088 123584 108128
rect 123626 108088 123666 108128
rect 123708 108088 123748 108128
rect 123790 108088 123830 108128
rect 123872 108088 123912 108128
rect 138664 108088 138704 108128
rect 138746 108088 138786 108128
rect 138828 108088 138868 108128
rect 138910 108088 138950 108128
rect 138992 108088 139032 108128
rect 79424 107332 79464 107372
rect 79506 107332 79546 107372
rect 79588 107332 79628 107372
rect 79670 107332 79710 107372
rect 79752 107332 79792 107372
rect 94544 107332 94584 107372
rect 94626 107332 94666 107372
rect 94708 107332 94748 107372
rect 94790 107332 94830 107372
rect 94872 107332 94912 107372
rect 109664 107332 109704 107372
rect 109746 107332 109786 107372
rect 109828 107332 109868 107372
rect 109910 107332 109950 107372
rect 109992 107332 110032 107372
rect 124784 107332 124824 107372
rect 124866 107332 124906 107372
rect 124948 107332 124988 107372
rect 125030 107332 125070 107372
rect 125112 107332 125152 107372
rect 139904 107332 139944 107372
rect 139986 107332 140026 107372
rect 140068 107332 140108 107372
rect 140150 107332 140190 107372
rect 140232 107332 140272 107372
rect 78184 106576 78224 106616
rect 78266 106576 78306 106616
rect 78348 106576 78388 106616
rect 78430 106576 78470 106616
rect 78512 106576 78552 106616
rect 93304 106576 93344 106616
rect 93386 106576 93426 106616
rect 93468 106576 93508 106616
rect 93550 106576 93590 106616
rect 93632 106576 93672 106616
rect 108424 106576 108464 106616
rect 108506 106576 108546 106616
rect 108588 106576 108628 106616
rect 108670 106576 108710 106616
rect 108752 106576 108792 106616
rect 123544 106576 123584 106616
rect 123626 106576 123666 106616
rect 123708 106576 123748 106616
rect 123790 106576 123830 106616
rect 123872 106576 123912 106616
rect 138664 106576 138704 106616
rect 138746 106576 138786 106616
rect 138828 106576 138868 106616
rect 138910 106576 138950 106616
rect 138992 106576 139032 106616
rect 79424 105820 79464 105860
rect 79506 105820 79546 105860
rect 79588 105820 79628 105860
rect 79670 105820 79710 105860
rect 79752 105820 79792 105860
rect 94544 105820 94584 105860
rect 94626 105820 94666 105860
rect 94708 105820 94748 105860
rect 94790 105820 94830 105860
rect 94872 105820 94912 105860
rect 109664 105820 109704 105860
rect 109746 105820 109786 105860
rect 109828 105820 109868 105860
rect 109910 105820 109950 105860
rect 109992 105820 110032 105860
rect 124784 105820 124824 105860
rect 124866 105820 124906 105860
rect 124948 105820 124988 105860
rect 125030 105820 125070 105860
rect 125112 105820 125152 105860
rect 139904 105820 139944 105860
rect 139986 105820 140026 105860
rect 140068 105820 140108 105860
rect 140150 105820 140190 105860
rect 140232 105820 140272 105860
rect 78184 105064 78224 105104
rect 78266 105064 78306 105104
rect 78348 105064 78388 105104
rect 78430 105064 78470 105104
rect 78512 105064 78552 105104
rect 93304 105064 93344 105104
rect 93386 105064 93426 105104
rect 93468 105064 93508 105104
rect 93550 105064 93590 105104
rect 93632 105064 93672 105104
rect 108424 105064 108464 105104
rect 108506 105064 108546 105104
rect 108588 105064 108628 105104
rect 108670 105064 108710 105104
rect 108752 105064 108792 105104
rect 123544 105064 123584 105104
rect 123626 105064 123666 105104
rect 123708 105064 123748 105104
rect 123790 105064 123830 105104
rect 123872 105064 123912 105104
rect 138664 105064 138704 105104
rect 138746 105064 138786 105104
rect 138828 105064 138868 105104
rect 138910 105064 138950 105104
rect 138992 105064 139032 105104
rect 79424 104308 79464 104348
rect 79506 104308 79546 104348
rect 79588 104308 79628 104348
rect 79670 104308 79710 104348
rect 79752 104308 79792 104348
rect 94544 104308 94584 104348
rect 94626 104308 94666 104348
rect 94708 104308 94748 104348
rect 94790 104308 94830 104348
rect 94872 104308 94912 104348
rect 109664 104308 109704 104348
rect 109746 104308 109786 104348
rect 109828 104308 109868 104348
rect 109910 104308 109950 104348
rect 109992 104308 110032 104348
rect 124784 104308 124824 104348
rect 124866 104308 124906 104348
rect 124948 104308 124988 104348
rect 125030 104308 125070 104348
rect 125112 104308 125152 104348
rect 139904 104308 139944 104348
rect 139986 104308 140026 104348
rect 140068 104308 140108 104348
rect 140150 104308 140190 104348
rect 140232 104308 140272 104348
rect 78184 103552 78224 103592
rect 78266 103552 78306 103592
rect 78348 103552 78388 103592
rect 78430 103552 78470 103592
rect 78512 103552 78552 103592
rect 93304 103552 93344 103592
rect 93386 103552 93426 103592
rect 93468 103552 93508 103592
rect 93550 103552 93590 103592
rect 93632 103552 93672 103592
rect 108424 103552 108464 103592
rect 108506 103552 108546 103592
rect 108588 103552 108628 103592
rect 108670 103552 108710 103592
rect 108752 103552 108792 103592
rect 123544 103552 123584 103592
rect 123626 103552 123666 103592
rect 123708 103552 123748 103592
rect 123790 103552 123830 103592
rect 123872 103552 123912 103592
rect 138664 103552 138704 103592
rect 138746 103552 138786 103592
rect 138828 103552 138868 103592
rect 138910 103552 138950 103592
rect 138992 103552 139032 103592
rect 79424 102796 79464 102836
rect 79506 102796 79546 102836
rect 79588 102796 79628 102836
rect 79670 102796 79710 102836
rect 79752 102796 79792 102836
rect 94544 102796 94584 102836
rect 94626 102796 94666 102836
rect 94708 102796 94748 102836
rect 94790 102796 94830 102836
rect 94872 102796 94912 102836
rect 109664 102796 109704 102836
rect 109746 102796 109786 102836
rect 109828 102796 109868 102836
rect 109910 102796 109950 102836
rect 109992 102796 110032 102836
rect 124784 102796 124824 102836
rect 124866 102796 124906 102836
rect 124948 102796 124988 102836
rect 125030 102796 125070 102836
rect 125112 102796 125152 102836
rect 139904 102796 139944 102836
rect 139986 102796 140026 102836
rect 140068 102796 140108 102836
rect 140150 102796 140190 102836
rect 140232 102796 140272 102836
rect 78184 102040 78224 102080
rect 78266 102040 78306 102080
rect 78348 102040 78388 102080
rect 78430 102040 78470 102080
rect 78512 102040 78552 102080
rect 93304 102040 93344 102080
rect 93386 102040 93426 102080
rect 93468 102040 93508 102080
rect 93550 102040 93590 102080
rect 93632 102040 93672 102080
rect 108424 102040 108464 102080
rect 108506 102040 108546 102080
rect 108588 102040 108628 102080
rect 108670 102040 108710 102080
rect 108752 102040 108792 102080
rect 123544 102040 123584 102080
rect 123626 102040 123666 102080
rect 123708 102040 123748 102080
rect 123790 102040 123830 102080
rect 123872 102040 123912 102080
rect 138664 102040 138704 102080
rect 138746 102040 138786 102080
rect 138828 102040 138868 102080
rect 138910 102040 138950 102080
rect 138992 102040 139032 102080
rect 79424 101284 79464 101324
rect 79506 101284 79546 101324
rect 79588 101284 79628 101324
rect 79670 101284 79710 101324
rect 79752 101284 79792 101324
rect 94544 101284 94584 101324
rect 94626 101284 94666 101324
rect 94708 101284 94748 101324
rect 94790 101284 94830 101324
rect 94872 101284 94912 101324
rect 109664 101284 109704 101324
rect 109746 101284 109786 101324
rect 109828 101284 109868 101324
rect 109910 101284 109950 101324
rect 109992 101284 110032 101324
rect 124784 101284 124824 101324
rect 124866 101284 124906 101324
rect 124948 101284 124988 101324
rect 125030 101284 125070 101324
rect 125112 101284 125152 101324
rect 139904 101284 139944 101324
rect 139986 101284 140026 101324
rect 140068 101284 140108 101324
rect 140150 101284 140190 101324
rect 140232 101284 140272 101324
rect 78184 100528 78224 100568
rect 78266 100528 78306 100568
rect 78348 100528 78388 100568
rect 78430 100528 78470 100568
rect 78512 100528 78552 100568
rect 93304 100528 93344 100568
rect 93386 100528 93426 100568
rect 93468 100528 93508 100568
rect 93550 100528 93590 100568
rect 93632 100528 93672 100568
rect 108424 100528 108464 100568
rect 108506 100528 108546 100568
rect 108588 100528 108628 100568
rect 108670 100528 108710 100568
rect 108752 100528 108792 100568
rect 123544 100528 123584 100568
rect 123626 100528 123666 100568
rect 123708 100528 123748 100568
rect 123790 100528 123830 100568
rect 123872 100528 123912 100568
rect 138664 100528 138704 100568
rect 138746 100528 138786 100568
rect 138828 100528 138868 100568
rect 138910 100528 138950 100568
rect 138992 100528 139032 100568
rect 79424 99772 79464 99812
rect 79506 99772 79546 99812
rect 79588 99772 79628 99812
rect 79670 99772 79710 99812
rect 79752 99772 79792 99812
rect 94544 99772 94584 99812
rect 94626 99772 94666 99812
rect 94708 99772 94748 99812
rect 94790 99772 94830 99812
rect 94872 99772 94912 99812
rect 109664 99772 109704 99812
rect 109746 99772 109786 99812
rect 109828 99772 109868 99812
rect 109910 99772 109950 99812
rect 109992 99772 110032 99812
rect 124784 99772 124824 99812
rect 124866 99772 124906 99812
rect 124948 99772 124988 99812
rect 125030 99772 125070 99812
rect 125112 99772 125152 99812
rect 139904 99772 139944 99812
rect 139986 99772 140026 99812
rect 140068 99772 140108 99812
rect 140150 99772 140190 99812
rect 140232 99772 140272 99812
rect 78184 99016 78224 99056
rect 78266 99016 78306 99056
rect 78348 99016 78388 99056
rect 78430 99016 78470 99056
rect 78512 99016 78552 99056
rect 93304 99016 93344 99056
rect 93386 99016 93426 99056
rect 93468 99016 93508 99056
rect 93550 99016 93590 99056
rect 93632 99016 93672 99056
rect 108424 99016 108464 99056
rect 108506 99016 108546 99056
rect 108588 99016 108628 99056
rect 108670 99016 108710 99056
rect 108752 99016 108792 99056
rect 123544 99016 123584 99056
rect 123626 99016 123666 99056
rect 123708 99016 123748 99056
rect 123790 99016 123830 99056
rect 123872 99016 123912 99056
rect 138664 99016 138704 99056
rect 138746 99016 138786 99056
rect 138828 99016 138868 99056
rect 138910 99016 138950 99056
rect 138992 99016 139032 99056
rect 79424 98260 79464 98300
rect 79506 98260 79546 98300
rect 79588 98260 79628 98300
rect 79670 98260 79710 98300
rect 79752 98260 79792 98300
rect 94544 98260 94584 98300
rect 94626 98260 94666 98300
rect 94708 98260 94748 98300
rect 94790 98260 94830 98300
rect 94872 98260 94912 98300
rect 109664 98260 109704 98300
rect 109746 98260 109786 98300
rect 109828 98260 109868 98300
rect 109910 98260 109950 98300
rect 109992 98260 110032 98300
rect 124784 98260 124824 98300
rect 124866 98260 124906 98300
rect 124948 98260 124988 98300
rect 125030 98260 125070 98300
rect 125112 98260 125152 98300
rect 139904 98260 139944 98300
rect 139986 98260 140026 98300
rect 140068 98260 140108 98300
rect 140150 98260 140190 98300
rect 140232 98260 140272 98300
rect 78184 97504 78224 97544
rect 78266 97504 78306 97544
rect 78348 97504 78388 97544
rect 78430 97504 78470 97544
rect 78512 97504 78552 97544
rect 93304 97504 93344 97544
rect 93386 97504 93426 97544
rect 93468 97504 93508 97544
rect 93550 97504 93590 97544
rect 93632 97504 93672 97544
rect 108424 97504 108464 97544
rect 108506 97504 108546 97544
rect 108588 97504 108628 97544
rect 108670 97504 108710 97544
rect 108752 97504 108792 97544
rect 123544 97504 123584 97544
rect 123626 97504 123666 97544
rect 123708 97504 123748 97544
rect 123790 97504 123830 97544
rect 123872 97504 123912 97544
rect 138664 97504 138704 97544
rect 138746 97504 138786 97544
rect 138828 97504 138868 97544
rect 138910 97504 138950 97544
rect 138992 97504 139032 97544
rect 79424 96748 79464 96788
rect 79506 96748 79546 96788
rect 79588 96748 79628 96788
rect 79670 96748 79710 96788
rect 79752 96748 79792 96788
rect 94544 96748 94584 96788
rect 94626 96748 94666 96788
rect 94708 96748 94748 96788
rect 94790 96748 94830 96788
rect 94872 96748 94912 96788
rect 109664 96748 109704 96788
rect 109746 96748 109786 96788
rect 109828 96748 109868 96788
rect 109910 96748 109950 96788
rect 109992 96748 110032 96788
rect 124784 96748 124824 96788
rect 124866 96748 124906 96788
rect 124948 96748 124988 96788
rect 125030 96748 125070 96788
rect 125112 96748 125152 96788
rect 139904 96748 139944 96788
rect 139986 96748 140026 96788
rect 140068 96748 140108 96788
rect 140150 96748 140190 96788
rect 140232 96748 140272 96788
rect 78184 95992 78224 96032
rect 78266 95992 78306 96032
rect 78348 95992 78388 96032
rect 78430 95992 78470 96032
rect 78512 95992 78552 96032
rect 93304 95992 93344 96032
rect 93386 95992 93426 96032
rect 93468 95992 93508 96032
rect 93550 95992 93590 96032
rect 93632 95992 93672 96032
rect 108424 95992 108464 96032
rect 108506 95992 108546 96032
rect 108588 95992 108628 96032
rect 108670 95992 108710 96032
rect 108752 95992 108792 96032
rect 123544 95992 123584 96032
rect 123626 95992 123666 96032
rect 123708 95992 123748 96032
rect 123790 95992 123830 96032
rect 123872 95992 123912 96032
rect 138664 95992 138704 96032
rect 138746 95992 138786 96032
rect 138828 95992 138868 96032
rect 138910 95992 138950 96032
rect 138992 95992 139032 96032
rect 79424 95236 79464 95276
rect 79506 95236 79546 95276
rect 79588 95236 79628 95276
rect 79670 95236 79710 95276
rect 79752 95236 79792 95276
rect 94544 95236 94584 95276
rect 94626 95236 94666 95276
rect 94708 95236 94748 95276
rect 94790 95236 94830 95276
rect 94872 95236 94912 95276
rect 109664 95236 109704 95276
rect 109746 95236 109786 95276
rect 109828 95236 109868 95276
rect 109910 95236 109950 95276
rect 109992 95236 110032 95276
rect 124784 95236 124824 95276
rect 124866 95236 124906 95276
rect 124948 95236 124988 95276
rect 125030 95236 125070 95276
rect 125112 95236 125152 95276
rect 139904 95236 139944 95276
rect 139986 95236 140026 95276
rect 140068 95236 140108 95276
rect 140150 95236 140190 95276
rect 140232 95236 140272 95276
rect 78184 94480 78224 94520
rect 78266 94480 78306 94520
rect 78348 94480 78388 94520
rect 78430 94480 78470 94520
rect 78512 94480 78552 94520
rect 93304 94480 93344 94520
rect 93386 94480 93426 94520
rect 93468 94480 93508 94520
rect 93550 94480 93590 94520
rect 93632 94480 93672 94520
rect 108424 94480 108464 94520
rect 108506 94480 108546 94520
rect 108588 94480 108628 94520
rect 108670 94480 108710 94520
rect 108752 94480 108792 94520
rect 123544 94480 123584 94520
rect 123626 94480 123666 94520
rect 123708 94480 123748 94520
rect 123790 94480 123830 94520
rect 123872 94480 123912 94520
rect 138664 94480 138704 94520
rect 138746 94480 138786 94520
rect 138828 94480 138868 94520
rect 138910 94480 138950 94520
rect 138992 94480 139032 94520
rect 79424 93724 79464 93764
rect 79506 93724 79546 93764
rect 79588 93724 79628 93764
rect 79670 93724 79710 93764
rect 79752 93724 79792 93764
rect 94544 93724 94584 93764
rect 94626 93724 94666 93764
rect 94708 93724 94748 93764
rect 94790 93724 94830 93764
rect 94872 93724 94912 93764
rect 109664 93724 109704 93764
rect 109746 93724 109786 93764
rect 109828 93724 109868 93764
rect 109910 93724 109950 93764
rect 109992 93724 110032 93764
rect 124784 93724 124824 93764
rect 124866 93724 124906 93764
rect 124948 93724 124988 93764
rect 125030 93724 125070 93764
rect 125112 93724 125152 93764
rect 139904 93724 139944 93764
rect 139986 93724 140026 93764
rect 140068 93724 140108 93764
rect 140150 93724 140190 93764
rect 140232 93724 140272 93764
rect 78184 92968 78224 93008
rect 78266 92968 78306 93008
rect 78348 92968 78388 93008
rect 78430 92968 78470 93008
rect 78512 92968 78552 93008
rect 93304 92968 93344 93008
rect 93386 92968 93426 93008
rect 93468 92968 93508 93008
rect 93550 92968 93590 93008
rect 93632 92968 93672 93008
rect 108424 92968 108464 93008
rect 108506 92968 108546 93008
rect 108588 92968 108628 93008
rect 108670 92968 108710 93008
rect 108752 92968 108792 93008
rect 123544 92968 123584 93008
rect 123626 92968 123666 93008
rect 123708 92968 123748 93008
rect 123790 92968 123830 93008
rect 123872 92968 123912 93008
rect 138664 92968 138704 93008
rect 138746 92968 138786 93008
rect 138828 92968 138868 93008
rect 138910 92968 138950 93008
rect 138992 92968 139032 93008
rect 79424 92212 79464 92252
rect 79506 92212 79546 92252
rect 79588 92212 79628 92252
rect 79670 92212 79710 92252
rect 79752 92212 79792 92252
rect 94544 92212 94584 92252
rect 94626 92212 94666 92252
rect 94708 92212 94748 92252
rect 94790 92212 94830 92252
rect 94872 92212 94912 92252
rect 109664 92212 109704 92252
rect 109746 92212 109786 92252
rect 109828 92212 109868 92252
rect 109910 92212 109950 92252
rect 109992 92212 110032 92252
rect 124784 92212 124824 92252
rect 124866 92212 124906 92252
rect 124948 92212 124988 92252
rect 125030 92212 125070 92252
rect 125112 92212 125152 92252
rect 139904 92212 139944 92252
rect 139986 92212 140026 92252
rect 140068 92212 140108 92252
rect 140150 92212 140190 92252
rect 140232 92212 140272 92252
rect 78184 91456 78224 91496
rect 78266 91456 78306 91496
rect 78348 91456 78388 91496
rect 78430 91456 78470 91496
rect 78512 91456 78552 91496
rect 93304 91456 93344 91496
rect 93386 91456 93426 91496
rect 93468 91456 93508 91496
rect 93550 91456 93590 91496
rect 93632 91456 93672 91496
rect 108424 91456 108464 91496
rect 108506 91456 108546 91496
rect 108588 91456 108628 91496
rect 108670 91456 108710 91496
rect 108752 91456 108792 91496
rect 123544 91456 123584 91496
rect 123626 91456 123666 91496
rect 123708 91456 123748 91496
rect 123790 91456 123830 91496
rect 123872 91456 123912 91496
rect 138664 91456 138704 91496
rect 138746 91456 138786 91496
rect 138828 91456 138868 91496
rect 138910 91456 138950 91496
rect 138992 91456 139032 91496
rect 79424 90700 79464 90740
rect 79506 90700 79546 90740
rect 79588 90700 79628 90740
rect 79670 90700 79710 90740
rect 79752 90700 79792 90740
rect 94544 90700 94584 90740
rect 94626 90700 94666 90740
rect 94708 90700 94748 90740
rect 94790 90700 94830 90740
rect 94872 90700 94912 90740
rect 109664 90700 109704 90740
rect 109746 90700 109786 90740
rect 109828 90700 109868 90740
rect 109910 90700 109950 90740
rect 109992 90700 110032 90740
rect 124784 90700 124824 90740
rect 124866 90700 124906 90740
rect 124948 90700 124988 90740
rect 125030 90700 125070 90740
rect 125112 90700 125152 90740
rect 139904 90700 139944 90740
rect 139986 90700 140026 90740
rect 140068 90700 140108 90740
rect 140150 90700 140190 90740
rect 140232 90700 140272 90740
rect 78184 89944 78224 89984
rect 78266 89944 78306 89984
rect 78348 89944 78388 89984
rect 78430 89944 78470 89984
rect 78512 89944 78552 89984
rect 93304 89944 93344 89984
rect 93386 89944 93426 89984
rect 93468 89944 93508 89984
rect 93550 89944 93590 89984
rect 93632 89944 93672 89984
rect 108424 89944 108464 89984
rect 108506 89944 108546 89984
rect 108588 89944 108628 89984
rect 108670 89944 108710 89984
rect 108752 89944 108792 89984
rect 123544 89944 123584 89984
rect 123626 89944 123666 89984
rect 123708 89944 123748 89984
rect 123790 89944 123830 89984
rect 123872 89944 123912 89984
rect 138664 89944 138704 89984
rect 138746 89944 138786 89984
rect 138828 89944 138868 89984
rect 138910 89944 138950 89984
rect 138992 89944 139032 89984
rect 79424 89188 79464 89228
rect 79506 89188 79546 89228
rect 79588 89188 79628 89228
rect 79670 89188 79710 89228
rect 79752 89188 79792 89228
rect 94544 89188 94584 89228
rect 94626 89188 94666 89228
rect 94708 89188 94748 89228
rect 94790 89188 94830 89228
rect 94872 89188 94912 89228
rect 109664 89188 109704 89228
rect 109746 89188 109786 89228
rect 109828 89188 109868 89228
rect 109910 89188 109950 89228
rect 109992 89188 110032 89228
rect 124784 89188 124824 89228
rect 124866 89188 124906 89228
rect 124948 89188 124988 89228
rect 125030 89188 125070 89228
rect 125112 89188 125152 89228
rect 139904 89188 139944 89228
rect 139986 89188 140026 89228
rect 140068 89188 140108 89228
rect 140150 89188 140190 89228
rect 140232 89188 140272 89228
rect 90700 89104 90740 89144
rect 92140 89104 92180 89144
rect 78184 88432 78224 88472
rect 78266 88432 78306 88472
rect 78348 88432 78388 88472
rect 78430 88432 78470 88472
rect 78512 88432 78552 88472
rect 93304 88432 93344 88472
rect 93386 88432 93426 88472
rect 93468 88432 93508 88472
rect 93550 88432 93590 88472
rect 93632 88432 93672 88472
rect 108424 88432 108464 88472
rect 108506 88432 108546 88472
rect 108588 88432 108628 88472
rect 108670 88432 108710 88472
rect 108752 88432 108792 88472
rect 123544 88432 123584 88472
rect 123626 88432 123666 88472
rect 123708 88432 123748 88472
rect 123790 88432 123830 88472
rect 123872 88432 123912 88472
rect 138664 88432 138704 88472
rect 138746 88432 138786 88472
rect 138828 88432 138868 88472
rect 138910 88432 138950 88472
rect 138992 88432 139032 88472
rect 79424 87676 79464 87716
rect 79506 87676 79546 87716
rect 79588 87676 79628 87716
rect 79670 87676 79710 87716
rect 79752 87676 79792 87716
rect 94544 87676 94584 87716
rect 94626 87676 94666 87716
rect 94708 87676 94748 87716
rect 94790 87676 94830 87716
rect 94872 87676 94912 87716
rect 109664 87676 109704 87716
rect 109746 87676 109786 87716
rect 109828 87676 109868 87716
rect 109910 87676 109950 87716
rect 109992 87676 110032 87716
rect 124784 87676 124824 87716
rect 124866 87676 124906 87716
rect 124948 87676 124988 87716
rect 125030 87676 125070 87716
rect 125112 87676 125152 87716
rect 139904 87676 139944 87716
rect 139986 87676 140026 87716
rect 140068 87676 140108 87716
rect 140150 87676 140190 87716
rect 140232 87676 140272 87716
rect 78184 86920 78224 86960
rect 78266 86920 78306 86960
rect 78348 86920 78388 86960
rect 78430 86920 78470 86960
rect 78512 86920 78552 86960
rect 93304 86920 93344 86960
rect 93386 86920 93426 86960
rect 93468 86920 93508 86960
rect 93550 86920 93590 86960
rect 93632 86920 93672 86960
rect 108424 86920 108464 86960
rect 108506 86920 108546 86960
rect 108588 86920 108628 86960
rect 108670 86920 108710 86960
rect 108752 86920 108792 86960
rect 123544 86920 123584 86960
rect 123626 86920 123666 86960
rect 123708 86920 123748 86960
rect 123790 86920 123830 86960
rect 123872 86920 123912 86960
rect 138664 86920 138704 86960
rect 138746 86920 138786 86960
rect 138828 86920 138868 86960
rect 138910 86920 138950 86960
rect 138992 86920 139032 86960
rect 79424 86164 79464 86204
rect 79506 86164 79546 86204
rect 79588 86164 79628 86204
rect 79670 86164 79710 86204
rect 79752 86164 79792 86204
rect 94544 86164 94584 86204
rect 94626 86164 94666 86204
rect 94708 86164 94748 86204
rect 94790 86164 94830 86204
rect 94872 86164 94912 86204
rect 109664 86164 109704 86204
rect 109746 86164 109786 86204
rect 109828 86164 109868 86204
rect 109910 86164 109950 86204
rect 109992 86164 110032 86204
rect 124784 86164 124824 86204
rect 124866 86164 124906 86204
rect 124948 86164 124988 86204
rect 125030 86164 125070 86204
rect 125112 86164 125152 86204
rect 139904 86164 139944 86204
rect 139986 86164 140026 86204
rect 140068 86164 140108 86204
rect 140150 86164 140190 86204
rect 140232 86164 140272 86204
rect 78184 85408 78224 85448
rect 78266 85408 78306 85448
rect 78348 85408 78388 85448
rect 78430 85408 78470 85448
rect 78512 85408 78552 85448
rect 93304 85408 93344 85448
rect 93386 85408 93426 85448
rect 93468 85408 93508 85448
rect 93550 85408 93590 85448
rect 93632 85408 93672 85448
rect 108424 85408 108464 85448
rect 108506 85408 108546 85448
rect 108588 85408 108628 85448
rect 108670 85408 108710 85448
rect 108752 85408 108792 85448
rect 123544 85408 123584 85448
rect 123626 85408 123666 85448
rect 123708 85408 123748 85448
rect 123790 85408 123830 85448
rect 123872 85408 123912 85448
rect 138664 85408 138704 85448
rect 138746 85408 138786 85448
rect 138828 85408 138868 85448
rect 138910 85408 138950 85448
rect 138992 85408 139032 85448
rect 79424 84652 79464 84692
rect 79506 84652 79546 84692
rect 79588 84652 79628 84692
rect 79670 84652 79710 84692
rect 79752 84652 79792 84692
rect 94544 84652 94584 84692
rect 94626 84652 94666 84692
rect 94708 84652 94748 84692
rect 94790 84652 94830 84692
rect 94872 84652 94912 84692
rect 109664 84652 109704 84692
rect 109746 84652 109786 84692
rect 109828 84652 109868 84692
rect 109910 84652 109950 84692
rect 109992 84652 110032 84692
rect 124784 84652 124824 84692
rect 124866 84652 124906 84692
rect 124948 84652 124988 84692
rect 125030 84652 125070 84692
rect 125112 84652 125152 84692
rect 139904 84652 139944 84692
rect 139986 84652 140026 84692
rect 140068 84652 140108 84692
rect 140150 84652 140190 84692
rect 140232 84652 140272 84692
rect 78184 83896 78224 83936
rect 78266 83896 78306 83936
rect 78348 83896 78388 83936
rect 78430 83896 78470 83936
rect 78512 83896 78552 83936
rect 93304 83896 93344 83936
rect 93386 83896 93426 83936
rect 93468 83896 93508 83936
rect 93550 83896 93590 83936
rect 93632 83896 93672 83936
rect 108424 83896 108464 83936
rect 108506 83896 108546 83936
rect 108588 83896 108628 83936
rect 108670 83896 108710 83936
rect 108752 83896 108792 83936
rect 123544 83896 123584 83936
rect 123626 83896 123666 83936
rect 123708 83896 123748 83936
rect 123790 83896 123830 83936
rect 123872 83896 123912 83936
rect 138664 83896 138704 83936
rect 138746 83896 138786 83936
rect 138828 83896 138868 83936
rect 138910 83896 138950 83936
rect 138992 83896 139032 83936
rect 79424 83140 79464 83180
rect 79506 83140 79546 83180
rect 79588 83140 79628 83180
rect 79670 83140 79710 83180
rect 79752 83140 79792 83180
rect 94544 83140 94584 83180
rect 94626 83140 94666 83180
rect 94708 83140 94748 83180
rect 94790 83140 94830 83180
rect 94872 83140 94912 83180
rect 109664 83140 109704 83180
rect 109746 83140 109786 83180
rect 109828 83140 109868 83180
rect 109910 83140 109950 83180
rect 109992 83140 110032 83180
rect 124784 83140 124824 83180
rect 124866 83140 124906 83180
rect 124948 83140 124988 83180
rect 125030 83140 125070 83180
rect 125112 83140 125152 83180
rect 139904 83140 139944 83180
rect 139986 83140 140026 83180
rect 140068 83140 140108 83180
rect 140150 83140 140190 83180
rect 140232 83140 140272 83180
rect 78184 82384 78224 82424
rect 78266 82384 78306 82424
rect 78348 82384 78388 82424
rect 78430 82384 78470 82424
rect 78512 82384 78552 82424
rect 93304 82384 93344 82424
rect 93386 82384 93426 82424
rect 93468 82384 93508 82424
rect 93550 82384 93590 82424
rect 93632 82384 93672 82424
rect 108424 82384 108464 82424
rect 108506 82384 108546 82424
rect 108588 82384 108628 82424
rect 108670 82384 108710 82424
rect 108752 82384 108792 82424
rect 123544 82384 123584 82424
rect 123626 82384 123666 82424
rect 123708 82384 123748 82424
rect 123790 82384 123830 82424
rect 123872 82384 123912 82424
rect 138664 82384 138704 82424
rect 138746 82384 138786 82424
rect 138828 82384 138868 82424
rect 138910 82384 138950 82424
rect 138992 82384 139032 82424
rect 79424 81628 79464 81668
rect 79506 81628 79546 81668
rect 79588 81628 79628 81668
rect 79670 81628 79710 81668
rect 79752 81628 79792 81668
rect 94544 81628 94584 81668
rect 94626 81628 94666 81668
rect 94708 81628 94748 81668
rect 94790 81628 94830 81668
rect 94872 81628 94912 81668
rect 109664 81628 109704 81668
rect 109746 81628 109786 81668
rect 109828 81628 109868 81668
rect 109910 81628 109950 81668
rect 109992 81628 110032 81668
rect 124784 81628 124824 81668
rect 124866 81628 124906 81668
rect 124948 81628 124988 81668
rect 125030 81628 125070 81668
rect 125112 81628 125152 81668
rect 139904 81628 139944 81668
rect 139986 81628 140026 81668
rect 140068 81628 140108 81668
rect 140150 81628 140190 81668
rect 140232 81628 140272 81668
rect 78184 80872 78224 80912
rect 78266 80872 78306 80912
rect 78348 80872 78388 80912
rect 78430 80872 78470 80912
rect 78512 80872 78552 80912
rect 93304 80872 93344 80912
rect 93386 80872 93426 80912
rect 93468 80872 93508 80912
rect 93550 80872 93590 80912
rect 93632 80872 93672 80912
rect 108424 80872 108464 80912
rect 108506 80872 108546 80912
rect 108588 80872 108628 80912
rect 108670 80872 108710 80912
rect 108752 80872 108792 80912
rect 123544 80872 123584 80912
rect 123626 80872 123666 80912
rect 123708 80872 123748 80912
rect 123790 80872 123830 80912
rect 123872 80872 123912 80912
rect 138664 80872 138704 80912
rect 138746 80872 138786 80912
rect 138828 80872 138868 80912
rect 138910 80872 138950 80912
rect 138992 80872 139032 80912
rect 79424 80116 79464 80156
rect 79506 80116 79546 80156
rect 79588 80116 79628 80156
rect 79670 80116 79710 80156
rect 79752 80116 79792 80156
rect 94544 80116 94584 80156
rect 94626 80116 94666 80156
rect 94708 80116 94748 80156
rect 94790 80116 94830 80156
rect 94872 80116 94912 80156
rect 109664 80116 109704 80156
rect 109746 80116 109786 80156
rect 109828 80116 109868 80156
rect 109910 80116 109950 80156
rect 109992 80116 110032 80156
rect 124784 80116 124824 80156
rect 124866 80116 124906 80156
rect 124948 80116 124988 80156
rect 125030 80116 125070 80156
rect 125112 80116 125152 80156
rect 139904 80116 139944 80156
rect 139986 80116 140026 80156
rect 140068 80116 140108 80156
rect 140150 80116 140190 80156
rect 140232 80116 140272 80156
rect 78184 79360 78224 79400
rect 78266 79360 78306 79400
rect 78348 79360 78388 79400
rect 78430 79360 78470 79400
rect 78512 79360 78552 79400
rect 93304 79360 93344 79400
rect 93386 79360 93426 79400
rect 93468 79360 93508 79400
rect 93550 79360 93590 79400
rect 93632 79360 93672 79400
rect 108424 79360 108464 79400
rect 108506 79360 108546 79400
rect 108588 79360 108628 79400
rect 108670 79360 108710 79400
rect 108752 79360 108792 79400
rect 123544 79360 123584 79400
rect 123626 79360 123666 79400
rect 123708 79360 123748 79400
rect 123790 79360 123830 79400
rect 123872 79360 123912 79400
rect 138664 79360 138704 79400
rect 138746 79360 138786 79400
rect 138828 79360 138868 79400
rect 138910 79360 138950 79400
rect 138992 79360 139032 79400
rect 79424 78604 79464 78644
rect 79506 78604 79546 78644
rect 79588 78604 79628 78644
rect 79670 78604 79710 78644
rect 79752 78604 79792 78644
rect 94544 78604 94584 78644
rect 94626 78604 94666 78644
rect 94708 78604 94748 78644
rect 94790 78604 94830 78644
rect 94872 78604 94912 78644
rect 109664 78604 109704 78644
rect 109746 78604 109786 78644
rect 109828 78604 109868 78644
rect 109910 78604 109950 78644
rect 109992 78604 110032 78644
rect 124784 78604 124824 78644
rect 124866 78604 124906 78644
rect 124948 78604 124988 78644
rect 125030 78604 125070 78644
rect 125112 78604 125152 78644
rect 139904 78604 139944 78644
rect 139986 78604 140026 78644
rect 140068 78604 140108 78644
rect 140150 78604 140190 78644
rect 140232 78604 140272 78644
rect 78184 77848 78224 77888
rect 78266 77848 78306 77888
rect 78348 77848 78388 77888
rect 78430 77848 78470 77888
rect 78512 77848 78552 77888
rect 93304 77848 93344 77888
rect 93386 77848 93426 77888
rect 93468 77848 93508 77888
rect 93550 77848 93590 77888
rect 93632 77848 93672 77888
rect 108424 77848 108464 77888
rect 108506 77848 108546 77888
rect 108588 77848 108628 77888
rect 108670 77848 108710 77888
rect 108752 77848 108792 77888
rect 123544 77848 123584 77888
rect 123626 77848 123666 77888
rect 123708 77848 123748 77888
rect 123790 77848 123830 77888
rect 123872 77848 123912 77888
rect 138664 77848 138704 77888
rect 138746 77848 138786 77888
rect 138828 77848 138868 77888
rect 138910 77848 138950 77888
rect 138992 77848 139032 77888
rect 79424 77092 79464 77132
rect 79506 77092 79546 77132
rect 79588 77092 79628 77132
rect 79670 77092 79710 77132
rect 79752 77092 79792 77132
rect 94544 77092 94584 77132
rect 94626 77092 94666 77132
rect 94708 77092 94748 77132
rect 94790 77092 94830 77132
rect 94872 77092 94912 77132
rect 109664 77092 109704 77132
rect 109746 77092 109786 77132
rect 109828 77092 109868 77132
rect 109910 77092 109950 77132
rect 109992 77092 110032 77132
rect 124784 77092 124824 77132
rect 124866 77092 124906 77132
rect 124948 77092 124988 77132
rect 125030 77092 125070 77132
rect 125112 77092 125152 77132
rect 139904 77092 139944 77132
rect 139986 77092 140026 77132
rect 140068 77092 140108 77132
rect 140150 77092 140190 77132
rect 140232 77092 140272 77132
rect 78184 76336 78224 76376
rect 78266 76336 78306 76376
rect 78348 76336 78388 76376
rect 78430 76336 78470 76376
rect 78512 76336 78552 76376
rect 93304 76336 93344 76376
rect 93386 76336 93426 76376
rect 93468 76336 93508 76376
rect 93550 76336 93590 76376
rect 93632 76336 93672 76376
rect 108424 76336 108464 76376
rect 108506 76336 108546 76376
rect 108588 76336 108628 76376
rect 108670 76336 108710 76376
rect 108752 76336 108792 76376
rect 123544 76336 123584 76376
rect 123626 76336 123666 76376
rect 123708 76336 123748 76376
rect 123790 76336 123830 76376
rect 123872 76336 123912 76376
rect 138664 76336 138704 76376
rect 138746 76336 138786 76376
rect 138828 76336 138868 76376
rect 138910 76336 138950 76376
rect 138992 76336 139032 76376
rect 79424 75580 79464 75620
rect 79506 75580 79546 75620
rect 79588 75580 79628 75620
rect 79670 75580 79710 75620
rect 79752 75580 79792 75620
rect 94544 75580 94584 75620
rect 94626 75580 94666 75620
rect 94708 75580 94748 75620
rect 94790 75580 94830 75620
rect 94872 75580 94912 75620
rect 109664 75580 109704 75620
rect 109746 75580 109786 75620
rect 109828 75580 109868 75620
rect 109910 75580 109950 75620
rect 109992 75580 110032 75620
rect 124784 75580 124824 75620
rect 124866 75580 124906 75620
rect 124948 75580 124988 75620
rect 125030 75580 125070 75620
rect 125112 75580 125152 75620
rect 139904 75580 139944 75620
rect 139986 75580 140026 75620
rect 140068 75580 140108 75620
rect 140150 75580 140190 75620
rect 140232 75580 140272 75620
rect 90700 71212 90740 71252
rect 92140 71212 92180 71252
<< metal5 >>
rect 79415 148196 79462 148238
rect 79586 148196 79630 148238
rect 79754 148196 79801 148238
rect 79415 148156 79424 148196
rect 79586 148156 79588 148196
rect 79628 148156 79630 148196
rect 79792 148156 79801 148196
rect 79415 148114 79462 148156
rect 79586 148114 79630 148156
rect 79754 148114 79801 148156
rect 94535 148196 94582 148238
rect 94706 148196 94750 148238
rect 94874 148196 94921 148238
rect 94535 148156 94544 148196
rect 94706 148156 94708 148196
rect 94748 148156 94750 148196
rect 94912 148156 94921 148196
rect 94535 148114 94582 148156
rect 94706 148114 94750 148156
rect 94874 148114 94921 148156
rect 109655 148196 109702 148238
rect 109826 148196 109870 148238
rect 109994 148196 110041 148238
rect 109655 148156 109664 148196
rect 109826 148156 109828 148196
rect 109868 148156 109870 148196
rect 110032 148156 110041 148196
rect 109655 148114 109702 148156
rect 109826 148114 109870 148156
rect 109994 148114 110041 148156
rect 124775 148196 124822 148238
rect 124946 148196 124990 148238
rect 125114 148196 125161 148238
rect 124775 148156 124784 148196
rect 124946 148156 124948 148196
rect 124988 148156 124990 148196
rect 125152 148156 125161 148196
rect 124775 148114 124822 148156
rect 124946 148114 124990 148156
rect 125114 148114 125161 148156
rect 139895 148196 139942 148238
rect 140066 148196 140110 148238
rect 140234 148196 140281 148238
rect 139895 148156 139904 148196
rect 140066 148156 140068 148196
rect 140108 148156 140110 148196
rect 140272 148156 140281 148196
rect 139895 148114 139942 148156
rect 140066 148114 140110 148156
rect 140234 148114 140281 148156
rect 78175 147440 78222 147482
rect 78346 147440 78390 147482
rect 78514 147440 78561 147482
rect 78175 147400 78184 147440
rect 78346 147400 78348 147440
rect 78388 147400 78390 147440
rect 78552 147400 78561 147440
rect 78175 147358 78222 147400
rect 78346 147358 78390 147400
rect 78514 147358 78561 147400
rect 93295 147440 93342 147482
rect 93466 147440 93510 147482
rect 93634 147440 93681 147482
rect 93295 147400 93304 147440
rect 93466 147400 93468 147440
rect 93508 147400 93510 147440
rect 93672 147400 93681 147440
rect 93295 147358 93342 147400
rect 93466 147358 93510 147400
rect 93634 147358 93681 147400
rect 108415 147440 108462 147482
rect 108586 147440 108630 147482
rect 108754 147440 108801 147482
rect 108415 147400 108424 147440
rect 108586 147400 108588 147440
rect 108628 147400 108630 147440
rect 108792 147400 108801 147440
rect 108415 147358 108462 147400
rect 108586 147358 108630 147400
rect 108754 147358 108801 147400
rect 123535 147440 123582 147482
rect 123706 147440 123750 147482
rect 123874 147440 123921 147482
rect 123535 147400 123544 147440
rect 123706 147400 123708 147440
rect 123748 147400 123750 147440
rect 123912 147400 123921 147440
rect 123535 147358 123582 147400
rect 123706 147358 123750 147400
rect 123874 147358 123921 147400
rect 138655 147440 138702 147482
rect 138826 147440 138870 147482
rect 138994 147440 139041 147482
rect 138655 147400 138664 147440
rect 138826 147400 138828 147440
rect 138868 147400 138870 147440
rect 139032 147400 139041 147440
rect 138655 147358 138702 147400
rect 138826 147358 138870 147400
rect 138994 147358 139041 147400
rect 79415 146684 79462 146726
rect 79586 146684 79630 146726
rect 79754 146684 79801 146726
rect 79415 146644 79424 146684
rect 79586 146644 79588 146684
rect 79628 146644 79630 146684
rect 79792 146644 79801 146684
rect 79415 146602 79462 146644
rect 79586 146602 79630 146644
rect 79754 146602 79801 146644
rect 94535 146684 94582 146726
rect 94706 146684 94750 146726
rect 94874 146684 94921 146726
rect 94535 146644 94544 146684
rect 94706 146644 94708 146684
rect 94748 146644 94750 146684
rect 94912 146644 94921 146684
rect 94535 146602 94582 146644
rect 94706 146602 94750 146644
rect 94874 146602 94921 146644
rect 109655 146684 109702 146726
rect 109826 146684 109870 146726
rect 109994 146684 110041 146726
rect 109655 146644 109664 146684
rect 109826 146644 109828 146684
rect 109868 146644 109870 146684
rect 110032 146644 110041 146684
rect 109655 146602 109702 146644
rect 109826 146602 109870 146644
rect 109994 146602 110041 146644
rect 124775 146684 124822 146726
rect 124946 146684 124990 146726
rect 125114 146684 125161 146726
rect 124775 146644 124784 146684
rect 124946 146644 124948 146684
rect 124988 146644 124990 146684
rect 125152 146644 125161 146684
rect 124775 146602 124822 146644
rect 124946 146602 124990 146644
rect 125114 146602 125161 146644
rect 139895 146684 139942 146726
rect 140066 146684 140110 146726
rect 140234 146684 140281 146726
rect 139895 146644 139904 146684
rect 140066 146644 140068 146684
rect 140108 146644 140110 146684
rect 140272 146644 140281 146684
rect 139895 146602 139942 146644
rect 140066 146602 140110 146644
rect 140234 146602 140281 146644
rect 78175 145928 78222 145970
rect 78346 145928 78390 145970
rect 78514 145928 78561 145970
rect 78175 145888 78184 145928
rect 78346 145888 78348 145928
rect 78388 145888 78390 145928
rect 78552 145888 78561 145928
rect 78175 145846 78222 145888
rect 78346 145846 78390 145888
rect 78514 145846 78561 145888
rect 93295 145928 93342 145970
rect 93466 145928 93510 145970
rect 93634 145928 93681 145970
rect 93295 145888 93304 145928
rect 93466 145888 93468 145928
rect 93508 145888 93510 145928
rect 93672 145888 93681 145928
rect 93295 145846 93342 145888
rect 93466 145846 93510 145888
rect 93634 145846 93681 145888
rect 108415 145928 108462 145970
rect 108586 145928 108630 145970
rect 108754 145928 108801 145970
rect 108415 145888 108424 145928
rect 108586 145888 108588 145928
rect 108628 145888 108630 145928
rect 108792 145888 108801 145928
rect 108415 145846 108462 145888
rect 108586 145846 108630 145888
rect 108754 145846 108801 145888
rect 123535 145928 123582 145970
rect 123706 145928 123750 145970
rect 123874 145928 123921 145970
rect 123535 145888 123544 145928
rect 123706 145888 123708 145928
rect 123748 145888 123750 145928
rect 123912 145888 123921 145928
rect 123535 145846 123582 145888
rect 123706 145846 123750 145888
rect 123874 145846 123921 145888
rect 138655 145928 138702 145970
rect 138826 145928 138870 145970
rect 138994 145928 139041 145970
rect 138655 145888 138664 145928
rect 138826 145888 138828 145928
rect 138868 145888 138870 145928
rect 139032 145888 139041 145928
rect 138655 145846 138702 145888
rect 138826 145846 138870 145888
rect 138994 145846 139041 145888
rect 79415 145172 79462 145214
rect 79586 145172 79630 145214
rect 79754 145172 79801 145214
rect 79415 145132 79424 145172
rect 79586 145132 79588 145172
rect 79628 145132 79630 145172
rect 79792 145132 79801 145172
rect 79415 145090 79462 145132
rect 79586 145090 79630 145132
rect 79754 145090 79801 145132
rect 94535 145172 94582 145214
rect 94706 145172 94750 145214
rect 94874 145172 94921 145214
rect 94535 145132 94544 145172
rect 94706 145132 94708 145172
rect 94748 145132 94750 145172
rect 94912 145132 94921 145172
rect 94535 145090 94582 145132
rect 94706 145090 94750 145132
rect 94874 145090 94921 145132
rect 109655 145172 109702 145214
rect 109826 145172 109870 145214
rect 109994 145172 110041 145214
rect 109655 145132 109664 145172
rect 109826 145132 109828 145172
rect 109868 145132 109870 145172
rect 110032 145132 110041 145172
rect 109655 145090 109702 145132
rect 109826 145090 109870 145132
rect 109994 145090 110041 145132
rect 124775 145172 124822 145214
rect 124946 145172 124990 145214
rect 125114 145172 125161 145214
rect 124775 145132 124784 145172
rect 124946 145132 124948 145172
rect 124988 145132 124990 145172
rect 125152 145132 125161 145172
rect 124775 145090 124822 145132
rect 124946 145090 124990 145132
rect 125114 145090 125161 145132
rect 139895 145172 139942 145214
rect 140066 145172 140110 145214
rect 140234 145172 140281 145214
rect 139895 145132 139904 145172
rect 140066 145132 140068 145172
rect 140108 145132 140110 145172
rect 140272 145132 140281 145172
rect 139895 145090 139942 145132
rect 140066 145090 140110 145132
rect 140234 145090 140281 145132
rect 78175 144416 78222 144458
rect 78346 144416 78390 144458
rect 78514 144416 78561 144458
rect 78175 144376 78184 144416
rect 78346 144376 78348 144416
rect 78388 144376 78390 144416
rect 78552 144376 78561 144416
rect 78175 144334 78222 144376
rect 78346 144334 78390 144376
rect 78514 144334 78561 144376
rect 93295 144416 93342 144458
rect 93466 144416 93510 144458
rect 93634 144416 93681 144458
rect 93295 144376 93304 144416
rect 93466 144376 93468 144416
rect 93508 144376 93510 144416
rect 93672 144376 93681 144416
rect 93295 144334 93342 144376
rect 93466 144334 93510 144376
rect 93634 144334 93681 144376
rect 108415 144416 108462 144458
rect 108586 144416 108630 144458
rect 108754 144416 108801 144458
rect 108415 144376 108424 144416
rect 108586 144376 108588 144416
rect 108628 144376 108630 144416
rect 108792 144376 108801 144416
rect 108415 144334 108462 144376
rect 108586 144334 108630 144376
rect 108754 144334 108801 144376
rect 123535 144416 123582 144458
rect 123706 144416 123750 144458
rect 123874 144416 123921 144458
rect 123535 144376 123544 144416
rect 123706 144376 123708 144416
rect 123748 144376 123750 144416
rect 123912 144376 123921 144416
rect 123535 144334 123582 144376
rect 123706 144334 123750 144376
rect 123874 144334 123921 144376
rect 138655 144416 138702 144458
rect 138826 144416 138870 144458
rect 138994 144416 139041 144458
rect 138655 144376 138664 144416
rect 138826 144376 138828 144416
rect 138868 144376 138870 144416
rect 139032 144376 139041 144416
rect 138655 144334 138702 144376
rect 138826 144334 138870 144376
rect 138994 144334 139041 144376
rect 79415 143660 79462 143702
rect 79586 143660 79630 143702
rect 79754 143660 79801 143702
rect 79415 143620 79424 143660
rect 79586 143620 79588 143660
rect 79628 143620 79630 143660
rect 79792 143620 79801 143660
rect 79415 143578 79462 143620
rect 79586 143578 79630 143620
rect 79754 143578 79801 143620
rect 94535 143660 94582 143702
rect 94706 143660 94750 143702
rect 94874 143660 94921 143702
rect 94535 143620 94544 143660
rect 94706 143620 94708 143660
rect 94748 143620 94750 143660
rect 94912 143620 94921 143660
rect 94535 143578 94582 143620
rect 94706 143578 94750 143620
rect 94874 143578 94921 143620
rect 109655 143660 109702 143702
rect 109826 143660 109870 143702
rect 109994 143660 110041 143702
rect 109655 143620 109664 143660
rect 109826 143620 109828 143660
rect 109868 143620 109870 143660
rect 110032 143620 110041 143660
rect 109655 143578 109702 143620
rect 109826 143578 109870 143620
rect 109994 143578 110041 143620
rect 124775 143660 124822 143702
rect 124946 143660 124990 143702
rect 125114 143660 125161 143702
rect 124775 143620 124784 143660
rect 124946 143620 124948 143660
rect 124988 143620 124990 143660
rect 125152 143620 125161 143660
rect 124775 143578 124822 143620
rect 124946 143578 124990 143620
rect 125114 143578 125161 143620
rect 139895 143660 139942 143702
rect 140066 143660 140110 143702
rect 140234 143660 140281 143702
rect 139895 143620 139904 143660
rect 140066 143620 140068 143660
rect 140108 143620 140110 143660
rect 140272 143620 140281 143660
rect 139895 143578 139942 143620
rect 140066 143578 140110 143620
rect 140234 143578 140281 143620
rect 78175 142904 78222 142946
rect 78346 142904 78390 142946
rect 78514 142904 78561 142946
rect 78175 142864 78184 142904
rect 78346 142864 78348 142904
rect 78388 142864 78390 142904
rect 78552 142864 78561 142904
rect 78175 142822 78222 142864
rect 78346 142822 78390 142864
rect 78514 142822 78561 142864
rect 93295 142904 93342 142946
rect 93466 142904 93510 142946
rect 93634 142904 93681 142946
rect 93295 142864 93304 142904
rect 93466 142864 93468 142904
rect 93508 142864 93510 142904
rect 93672 142864 93681 142904
rect 93295 142822 93342 142864
rect 93466 142822 93510 142864
rect 93634 142822 93681 142864
rect 108415 142904 108462 142946
rect 108586 142904 108630 142946
rect 108754 142904 108801 142946
rect 108415 142864 108424 142904
rect 108586 142864 108588 142904
rect 108628 142864 108630 142904
rect 108792 142864 108801 142904
rect 108415 142822 108462 142864
rect 108586 142822 108630 142864
rect 108754 142822 108801 142864
rect 123535 142904 123582 142946
rect 123706 142904 123750 142946
rect 123874 142904 123921 142946
rect 123535 142864 123544 142904
rect 123706 142864 123708 142904
rect 123748 142864 123750 142904
rect 123912 142864 123921 142904
rect 123535 142822 123582 142864
rect 123706 142822 123750 142864
rect 123874 142822 123921 142864
rect 138655 142904 138702 142946
rect 138826 142904 138870 142946
rect 138994 142904 139041 142946
rect 138655 142864 138664 142904
rect 138826 142864 138828 142904
rect 138868 142864 138870 142904
rect 139032 142864 139041 142904
rect 138655 142822 138702 142864
rect 138826 142822 138870 142864
rect 138994 142822 139041 142864
rect 79415 142148 79462 142190
rect 79586 142148 79630 142190
rect 79754 142148 79801 142190
rect 79415 142108 79424 142148
rect 79586 142108 79588 142148
rect 79628 142108 79630 142148
rect 79792 142108 79801 142148
rect 79415 142066 79462 142108
rect 79586 142066 79630 142108
rect 79754 142066 79801 142108
rect 94535 142148 94582 142190
rect 94706 142148 94750 142190
rect 94874 142148 94921 142190
rect 94535 142108 94544 142148
rect 94706 142108 94708 142148
rect 94748 142108 94750 142148
rect 94912 142108 94921 142148
rect 94535 142066 94582 142108
rect 94706 142066 94750 142108
rect 94874 142066 94921 142108
rect 109655 142148 109702 142190
rect 109826 142148 109870 142190
rect 109994 142148 110041 142190
rect 109655 142108 109664 142148
rect 109826 142108 109828 142148
rect 109868 142108 109870 142148
rect 110032 142108 110041 142148
rect 109655 142066 109702 142108
rect 109826 142066 109870 142108
rect 109994 142066 110041 142108
rect 124775 142148 124822 142190
rect 124946 142148 124990 142190
rect 125114 142148 125161 142190
rect 124775 142108 124784 142148
rect 124946 142108 124948 142148
rect 124988 142108 124990 142148
rect 125152 142108 125161 142148
rect 124775 142066 124822 142108
rect 124946 142066 124990 142108
rect 125114 142066 125161 142108
rect 139895 142148 139942 142190
rect 140066 142148 140110 142190
rect 140234 142148 140281 142190
rect 139895 142108 139904 142148
rect 140066 142108 140068 142148
rect 140108 142108 140110 142148
rect 140272 142108 140281 142148
rect 139895 142066 139942 142108
rect 140066 142066 140110 142108
rect 140234 142066 140281 142108
rect 78175 141392 78222 141434
rect 78346 141392 78390 141434
rect 78514 141392 78561 141434
rect 78175 141352 78184 141392
rect 78346 141352 78348 141392
rect 78388 141352 78390 141392
rect 78552 141352 78561 141392
rect 78175 141310 78222 141352
rect 78346 141310 78390 141352
rect 78514 141310 78561 141352
rect 93295 141392 93342 141434
rect 93466 141392 93510 141434
rect 93634 141392 93681 141434
rect 93295 141352 93304 141392
rect 93466 141352 93468 141392
rect 93508 141352 93510 141392
rect 93672 141352 93681 141392
rect 93295 141310 93342 141352
rect 93466 141310 93510 141352
rect 93634 141310 93681 141352
rect 108415 141392 108462 141434
rect 108586 141392 108630 141434
rect 108754 141392 108801 141434
rect 108415 141352 108424 141392
rect 108586 141352 108588 141392
rect 108628 141352 108630 141392
rect 108792 141352 108801 141392
rect 108415 141310 108462 141352
rect 108586 141310 108630 141352
rect 108754 141310 108801 141352
rect 123535 141392 123582 141434
rect 123706 141392 123750 141434
rect 123874 141392 123921 141434
rect 123535 141352 123544 141392
rect 123706 141352 123708 141392
rect 123748 141352 123750 141392
rect 123912 141352 123921 141392
rect 123535 141310 123582 141352
rect 123706 141310 123750 141352
rect 123874 141310 123921 141352
rect 138655 141392 138702 141434
rect 138826 141392 138870 141434
rect 138994 141392 139041 141434
rect 138655 141352 138664 141392
rect 138826 141352 138828 141392
rect 138868 141352 138870 141392
rect 139032 141352 139041 141392
rect 138655 141310 138702 141352
rect 138826 141310 138870 141352
rect 138994 141310 139041 141352
rect 79415 140636 79462 140678
rect 79586 140636 79630 140678
rect 79754 140636 79801 140678
rect 79415 140596 79424 140636
rect 79586 140596 79588 140636
rect 79628 140596 79630 140636
rect 79792 140596 79801 140636
rect 79415 140554 79462 140596
rect 79586 140554 79630 140596
rect 79754 140554 79801 140596
rect 94535 140636 94582 140678
rect 94706 140636 94750 140678
rect 94874 140636 94921 140678
rect 94535 140596 94544 140636
rect 94706 140596 94708 140636
rect 94748 140596 94750 140636
rect 94912 140596 94921 140636
rect 94535 140554 94582 140596
rect 94706 140554 94750 140596
rect 94874 140554 94921 140596
rect 109655 140636 109702 140678
rect 109826 140636 109870 140678
rect 109994 140636 110041 140678
rect 109655 140596 109664 140636
rect 109826 140596 109828 140636
rect 109868 140596 109870 140636
rect 110032 140596 110041 140636
rect 109655 140554 109702 140596
rect 109826 140554 109870 140596
rect 109994 140554 110041 140596
rect 124775 140636 124822 140678
rect 124946 140636 124990 140678
rect 125114 140636 125161 140678
rect 124775 140596 124784 140636
rect 124946 140596 124948 140636
rect 124988 140596 124990 140636
rect 125152 140596 125161 140636
rect 124775 140554 124822 140596
rect 124946 140554 124990 140596
rect 125114 140554 125161 140596
rect 139895 140636 139942 140678
rect 140066 140636 140110 140678
rect 140234 140636 140281 140678
rect 139895 140596 139904 140636
rect 140066 140596 140068 140636
rect 140108 140596 140110 140636
rect 140272 140596 140281 140636
rect 139895 140554 139942 140596
rect 140066 140554 140110 140596
rect 140234 140554 140281 140596
rect 78175 139880 78222 139922
rect 78346 139880 78390 139922
rect 78514 139880 78561 139922
rect 78175 139840 78184 139880
rect 78346 139840 78348 139880
rect 78388 139840 78390 139880
rect 78552 139840 78561 139880
rect 78175 139798 78222 139840
rect 78346 139798 78390 139840
rect 78514 139798 78561 139840
rect 93295 139880 93342 139922
rect 93466 139880 93510 139922
rect 93634 139880 93681 139922
rect 93295 139840 93304 139880
rect 93466 139840 93468 139880
rect 93508 139840 93510 139880
rect 93672 139840 93681 139880
rect 93295 139798 93342 139840
rect 93466 139798 93510 139840
rect 93634 139798 93681 139840
rect 108415 139880 108462 139922
rect 108586 139880 108630 139922
rect 108754 139880 108801 139922
rect 108415 139840 108424 139880
rect 108586 139840 108588 139880
rect 108628 139840 108630 139880
rect 108792 139840 108801 139880
rect 108415 139798 108462 139840
rect 108586 139798 108630 139840
rect 108754 139798 108801 139840
rect 123535 139880 123582 139922
rect 123706 139880 123750 139922
rect 123874 139880 123921 139922
rect 123535 139840 123544 139880
rect 123706 139840 123708 139880
rect 123748 139840 123750 139880
rect 123912 139840 123921 139880
rect 123535 139798 123582 139840
rect 123706 139798 123750 139840
rect 123874 139798 123921 139840
rect 138655 139880 138702 139922
rect 138826 139880 138870 139922
rect 138994 139880 139041 139922
rect 138655 139840 138664 139880
rect 138826 139840 138828 139880
rect 138868 139840 138870 139880
rect 139032 139840 139041 139880
rect 138655 139798 138702 139840
rect 138826 139798 138870 139840
rect 138994 139798 139041 139840
rect 79415 139124 79462 139166
rect 79586 139124 79630 139166
rect 79754 139124 79801 139166
rect 79415 139084 79424 139124
rect 79586 139084 79588 139124
rect 79628 139084 79630 139124
rect 79792 139084 79801 139124
rect 79415 139042 79462 139084
rect 79586 139042 79630 139084
rect 79754 139042 79801 139084
rect 94535 139124 94582 139166
rect 94706 139124 94750 139166
rect 94874 139124 94921 139166
rect 94535 139084 94544 139124
rect 94706 139084 94708 139124
rect 94748 139084 94750 139124
rect 94912 139084 94921 139124
rect 94535 139042 94582 139084
rect 94706 139042 94750 139084
rect 94874 139042 94921 139084
rect 109655 139124 109702 139166
rect 109826 139124 109870 139166
rect 109994 139124 110041 139166
rect 109655 139084 109664 139124
rect 109826 139084 109828 139124
rect 109868 139084 109870 139124
rect 110032 139084 110041 139124
rect 109655 139042 109702 139084
rect 109826 139042 109870 139084
rect 109994 139042 110041 139084
rect 124775 139124 124822 139166
rect 124946 139124 124990 139166
rect 125114 139124 125161 139166
rect 124775 139084 124784 139124
rect 124946 139084 124948 139124
rect 124988 139084 124990 139124
rect 125152 139084 125161 139124
rect 124775 139042 124822 139084
rect 124946 139042 124990 139084
rect 125114 139042 125161 139084
rect 139895 139124 139942 139166
rect 140066 139124 140110 139166
rect 140234 139124 140281 139166
rect 139895 139084 139904 139124
rect 140066 139084 140068 139124
rect 140108 139084 140110 139124
rect 140272 139084 140281 139124
rect 139895 139042 139942 139084
rect 140066 139042 140110 139084
rect 140234 139042 140281 139084
rect 78175 138368 78222 138410
rect 78346 138368 78390 138410
rect 78514 138368 78561 138410
rect 78175 138328 78184 138368
rect 78346 138328 78348 138368
rect 78388 138328 78390 138368
rect 78552 138328 78561 138368
rect 78175 138286 78222 138328
rect 78346 138286 78390 138328
rect 78514 138286 78561 138328
rect 93295 138368 93342 138410
rect 93466 138368 93510 138410
rect 93634 138368 93681 138410
rect 93295 138328 93304 138368
rect 93466 138328 93468 138368
rect 93508 138328 93510 138368
rect 93672 138328 93681 138368
rect 93295 138286 93342 138328
rect 93466 138286 93510 138328
rect 93634 138286 93681 138328
rect 108415 138368 108462 138410
rect 108586 138368 108630 138410
rect 108754 138368 108801 138410
rect 108415 138328 108424 138368
rect 108586 138328 108588 138368
rect 108628 138328 108630 138368
rect 108792 138328 108801 138368
rect 108415 138286 108462 138328
rect 108586 138286 108630 138328
rect 108754 138286 108801 138328
rect 123535 138368 123582 138410
rect 123706 138368 123750 138410
rect 123874 138368 123921 138410
rect 123535 138328 123544 138368
rect 123706 138328 123708 138368
rect 123748 138328 123750 138368
rect 123912 138328 123921 138368
rect 123535 138286 123582 138328
rect 123706 138286 123750 138328
rect 123874 138286 123921 138328
rect 138655 138368 138702 138410
rect 138826 138368 138870 138410
rect 138994 138368 139041 138410
rect 138655 138328 138664 138368
rect 138826 138328 138828 138368
rect 138868 138328 138870 138368
rect 139032 138328 139041 138368
rect 138655 138286 138702 138328
rect 138826 138286 138870 138328
rect 138994 138286 139041 138328
rect 79415 137612 79462 137654
rect 79586 137612 79630 137654
rect 79754 137612 79801 137654
rect 79415 137572 79424 137612
rect 79586 137572 79588 137612
rect 79628 137572 79630 137612
rect 79792 137572 79801 137612
rect 79415 137530 79462 137572
rect 79586 137530 79630 137572
rect 79754 137530 79801 137572
rect 94535 137612 94582 137654
rect 94706 137612 94750 137654
rect 94874 137612 94921 137654
rect 94535 137572 94544 137612
rect 94706 137572 94708 137612
rect 94748 137572 94750 137612
rect 94912 137572 94921 137612
rect 94535 137530 94582 137572
rect 94706 137530 94750 137572
rect 94874 137530 94921 137572
rect 109655 137612 109702 137654
rect 109826 137612 109870 137654
rect 109994 137612 110041 137654
rect 109655 137572 109664 137612
rect 109826 137572 109828 137612
rect 109868 137572 109870 137612
rect 110032 137572 110041 137612
rect 109655 137530 109702 137572
rect 109826 137530 109870 137572
rect 109994 137530 110041 137572
rect 124775 137612 124822 137654
rect 124946 137612 124990 137654
rect 125114 137612 125161 137654
rect 124775 137572 124784 137612
rect 124946 137572 124948 137612
rect 124988 137572 124990 137612
rect 125152 137572 125161 137612
rect 124775 137530 124822 137572
rect 124946 137530 124990 137572
rect 125114 137530 125161 137572
rect 139895 137612 139942 137654
rect 140066 137612 140110 137654
rect 140234 137612 140281 137654
rect 139895 137572 139904 137612
rect 140066 137572 140068 137612
rect 140108 137572 140110 137612
rect 140272 137572 140281 137612
rect 139895 137530 139942 137572
rect 140066 137530 140110 137572
rect 140234 137530 140281 137572
rect 78175 136856 78222 136898
rect 78346 136856 78390 136898
rect 78514 136856 78561 136898
rect 78175 136816 78184 136856
rect 78346 136816 78348 136856
rect 78388 136816 78390 136856
rect 78552 136816 78561 136856
rect 78175 136774 78222 136816
rect 78346 136774 78390 136816
rect 78514 136774 78561 136816
rect 93295 136856 93342 136898
rect 93466 136856 93510 136898
rect 93634 136856 93681 136898
rect 93295 136816 93304 136856
rect 93466 136816 93468 136856
rect 93508 136816 93510 136856
rect 93672 136816 93681 136856
rect 93295 136774 93342 136816
rect 93466 136774 93510 136816
rect 93634 136774 93681 136816
rect 108415 136856 108462 136898
rect 108586 136856 108630 136898
rect 108754 136856 108801 136898
rect 108415 136816 108424 136856
rect 108586 136816 108588 136856
rect 108628 136816 108630 136856
rect 108792 136816 108801 136856
rect 108415 136774 108462 136816
rect 108586 136774 108630 136816
rect 108754 136774 108801 136816
rect 123535 136856 123582 136898
rect 123706 136856 123750 136898
rect 123874 136856 123921 136898
rect 123535 136816 123544 136856
rect 123706 136816 123708 136856
rect 123748 136816 123750 136856
rect 123912 136816 123921 136856
rect 123535 136774 123582 136816
rect 123706 136774 123750 136816
rect 123874 136774 123921 136816
rect 138655 136856 138702 136898
rect 138826 136856 138870 136898
rect 138994 136856 139041 136898
rect 138655 136816 138664 136856
rect 138826 136816 138828 136856
rect 138868 136816 138870 136856
rect 139032 136816 139041 136856
rect 138655 136774 138702 136816
rect 138826 136774 138870 136816
rect 138994 136774 139041 136816
rect 79415 136100 79462 136142
rect 79586 136100 79630 136142
rect 79754 136100 79801 136142
rect 79415 136060 79424 136100
rect 79586 136060 79588 136100
rect 79628 136060 79630 136100
rect 79792 136060 79801 136100
rect 79415 136018 79462 136060
rect 79586 136018 79630 136060
rect 79754 136018 79801 136060
rect 94535 136100 94582 136142
rect 94706 136100 94750 136142
rect 94874 136100 94921 136142
rect 94535 136060 94544 136100
rect 94706 136060 94708 136100
rect 94748 136060 94750 136100
rect 94912 136060 94921 136100
rect 94535 136018 94582 136060
rect 94706 136018 94750 136060
rect 94874 136018 94921 136060
rect 109655 136100 109702 136142
rect 109826 136100 109870 136142
rect 109994 136100 110041 136142
rect 109655 136060 109664 136100
rect 109826 136060 109828 136100
rect 109868 136060 109870 136100
rect 110032 136060 110041 136100
rect 109655 136018 109702 136060
rect 109826 136018 109870 136060
rect 109994 136018 110041 136060
rect 124775 136100 124822 136142
rect 124946 136100 124990 136142
rect 125114 136100 125161 136142
rect 124775 136060 124784 136100
rect 124946 136060 124948 136100
rect 124988 136060 124990 136100
rect 125152 136060 125161 136100
rect 124775 136018 124822 136060
rect 124946 136018 124990 136060
rect 125114 136018 125161 136060
rect 139895 136100 139942 136142
rect 140066 136100 140110 136142
rect 140234 136100 140281 136142
rect 139895 136060 139904 136100
rect 140066 136060 140068 136100
rect 140108 136060 140110 136100
rect 140272 136060 140281 136100
rect 139895 136018 139942 136060
rect 140066 136018 140110 136060
rect 140234 136018 140281 136060
rect 78175 135344 78222 135386
rect 78346 135344 78390 135386
rect 78514 135344 78561 135386
rect 78175 135304 78184 135344
rect 78346 135304 78348 135344
rect 78388 135304 78390 135344
rect 78552 135304 78561 135344
rect 78175 135262 78222 135304
rect 78346 135262 78390 135304
rect 78514 135262 78561 135304
rect 93295 135344 93342 135386
rect 93466 135344 93510 135386
rect 93634 135344 93681 135386
rect 93295 135304 93304 135344
rect 93466 135304 93468 135344
rect 93508 135304 93510 135344
rect 93672 135304 93681 135344
rect 93295 135262 93342 135304
rect 93466 135262 93510 135304
rect 93634 135262 93681 135304
rect 108415 135344 108462 135386
rect 108586 135344 108630 135386
rect 108754 135344 108801 135386
rect 108415 135304 108424 135344
rect 108586 135304 108588 135344
rect 108628 135304 108630 135344
rect 108792 135304 108801 135344
rect 108415 135262 108462 135304
rect 108586 135262 108630 135304
rect 108754 135262 108801 135304
rect 123535 135344 123582 135386
rect 123706 135344 123750 135386
rect 123874 135344 123921 135386
rect 123535 135304 123544 135344
rect 123706 135304 123708 135344
rect 123748 135304 123750 135344
rect 123912 135304 123921 135344
rect 123535 135262 123582 135304
rect 123706 135262 123750 135304
rect 123874 135262 123921 135304
rect 138655 135344 138702 135386
rect 138826 135344 138870 135386
rect 138994 135344 139041 135386
rect 138655 135304 138664 135344
rect 138826 135304 138828 135344
rect 138868 135304 138870 135344
rect 139032 135304 139041 135344
rect 138655 135262 138702 135304
rect 138826 135262 138870 135304
rect 138994 135262 139041 135304
rect 79415 134588 79462 134630
rect 79586 134588 79630 134630
rect 79754 134588 79801 134630
rect 79415 134548 79424 134588
rect 79586 134548 79588 134588
rect 79628 134548 79630 134588
rect 79792 134548 79801 134588
rect 79415 134506 79462 134548
rect 79586 134506 79630 134548
rect 79754 134506 79801 134548
rect 94535 134588 94582 134630
rect 94706 134588 94750 134630
rect 94874 134588 94921 134630
rect 94535 134548 94544 134588
rect 94706 134548 94708 134588
rect 94748 134548 94750 134588
rect 94912 134548 94921 134588
rect 94535 134506 94582 134548
rect 94706 134506 94750 134548
rect 94874 134506 94921 134548
rect 109655 134588 109702 134630
rect 109826 134588 109870 134630
rect 109994 134588 110041 134630
rect 109655 134548 109664 134588
rect 109826 134548 109828 134588
rect 109868 134548 109870 134588
rect 110032 134548 110041 134588
rect 109655 134506 109702 134548
rect 109826 134506 109870 134548
rect 109994 134506 110041 134548
rect 124775 134588 124822 134630
rect 124946 134588 124990 134630
rect 125114 134588 125161 134630
rect 124775 134548 124784 134588
rect 124946 134548 124948 134588
rect 124988 134548 124990 134588
rect 125152 134548 125161 134588
rect 124775 134506 124822 134548
rect 124946 134506 124990 134548
rect 125114 134506 125161 134548
rect 139895 134588 139942 134630
rect 140066 134588 140110 134630
rect 140234 134588 140281 134630
rect 139895 134548 139904 134588
rect 140066 134548 140068 134588
rect 140108 134548 140110 134588
rect 140272 134548 140281 134588
rect 139895 134506 139942 134548
rect 140066 134506 140110 134548
rect 140234 134506 140281 134548
rect 78175 133832 78222 133874
rect 78346 133832 78390 133874
rect 78514 133832 78561 133874
rect 78175 133792 78184 133832
rect 78346 133792 78348 133832
rect 78388 133792 78390 133832
rect 78552 133792 78561 133832
rect 78175 133750 78222 133792
rect 78346 133750 78390 133792
rect 78514 133750 78561 133792
rect 93295 133832 93342 133874
rect 93466 133832 93510 133874
rect 93634 133832 93681 133874
rect 93295 133792 93304 133832
rect 93466 133792 93468 133832
rect 93508 133792 93510 133832
rect 93672 133792 93681 133832
rect 93295 133750 93342 133792
rect 93466 133750 93510 133792
rect 93634 133750 93681 133792
rect 108415 133832 108462 133874
rect 108586 133832 108630 133874
rect 108754 133832 108801 133874
rect 108415 133792 108424 133832
rect 108586 133792 108588 133832
rect 108628 133792 108630 133832
rect 108792 133792 108801 133832
rect 108415 133750 108462 133792
rect 108586 133750 108630 133792
rect 108754 133750 108801 133792
rect 123535 133832 123582 133874
rect 123706 133832 123750 133874
rect 123874 133832 123921 133874
rect 123535 133792 123544 133832
rect 123706 133792 123708 133832
rect 123748 133792 123750 133832
rect 123912 133792 123921 133832
rect 123535 133750 123582 133792
rect 123706 133750 123750 133792
rect 123874 133750 123921 133792
rect 138655 133832 138702 133874
rect 138826 133832 138870 133874
rect 138994 133832 139041 133874
rect 138655 133792 138664 133832
rect 138826 133792 138828 133832
rect 138868 133792 138870 133832
rect 139032 133792 139041 133832
rect 138655 133750 138702 133792
rect 138826 133750 138870 133792
rect 138994 133750 139041 133792
rect 79415 133076 79462 133118
rect 79586 133076 79630 133118
rect 79754 133076 79801 133118
rect 79415 133036 79424 133076
rect 79586 133036 79588 133076
rect 79628 133036 79630 133076
rect 79792 133036 79801 133076
rect 79415 132994 79462 133036
rect 79586 132994 79630 133036
rect 79754 132994 79801 133036
rect 94535 133076 94582 133118
rect 94706 133076 94750 133118
rect 94874 133076 94921 133118
rect 94535 133036 94544 133076
rect 94706 133036 94708 133076
rect 94748 133036 94750 133076
rect 94912 133036 94921 133076
rect 94535 132994 94582 133036
rect 94706 132994 94750 133036
rect 94874 132994 94921 133036
rect 109655 133076 109702 133118
rect 109826 133076 109870 133118
rect 109994 133076 110041 133118
rect 109655 133036 109664 133076
rect 109826 133036 109828 133076
rect 109868 133036 109870 133076
rect 110032 133036 110041 133076
rect 109655 132994 109702 133036
rect 109826 132994 109870 133036
rect 109994 132994 110041 133036
rect 124775 133076 124822 133118
rect 124946 133076 124990 133118
rect 125114 133076 125161 133118
rect 124775 133036 124784 133076
rect 124946 133036 124948 133076
rect 124988 133036 124990 133076
rect 125152 133036 125161 133076
rect 124775 132994 124822 133036
rect 124946 132994 124990 133036
rect 125114 132994 125161 133036
rect 139895 133076 139942 133118
rect 140066 133076 140110 133118
rect 140234 133076 140281 133118
rect 139895 133036 139904 133076
rect 140066 133036 140068 133076
rect 140108 133036 140110 133076
rect 140272 133036 140281 133076
rect 139895 132994 139942 133036
rect 140066 132994 140110 133036
rect 140234 132994 140281 133036
rect 78175 132320 78222 132362
rect 78346 132320 78390 132362
rect 78514 132320 78561 132362
rect 78175 132280 78184 132320
rect 78346 132280 78348 132320
rect 78388 132280 78390 132320
rect 78552 132280 78561 132320
rect 78175 132238 78222 132280
rect 78346 132238 78390 132280
rect 78514 132238 78561 132280
rect 93295 132320 93342 132362
rect 93466 132320 93510 132362
rect 93634 132320 93681 132362
rect 93295 132280 93304 132320
rect 93466 132280 93468 132320
rect 93508 132280 93510 132320
rect 93672 132280 93681 132320
rect 93295 132238 93342 132280
rect 93466 132238 93510 132280
rect 93634 132238 93681 132280
rect 108415 132320 108462 132362
rect 108586 132320 108630 132362
rect 108754 132320 108801 132362
rect 108415 132280 108424 132320
rect 108586 132280 108588 132320
rect 108628 132280 108630 132320
rect 108792 132280 108801 132320
rect 108415 132238 108462 132280
rect 108586 132238 108630 132280
rect 108754 132238 108801 132280
rect 123535 132320 123582 132362
rect 123706 132320 123750 132362
rect 123874 132320 123921 132362
rect 123535 132280 123544 132320
rect 123706 132280 123708 132320
rect 123748 132280 123750 132320
rect 123912 132280 123921 132320
rect 123535 132238 123582 132280
rect 123706 132238 123750 132280
rect 123874 132238 123921 132280
rect 138655 132320 138702 132362
rect 138826 132320 138870 132362
rect 138994 132320 139041 132362
rect 138655 132280 138664 132320
rect 138826 132280 138828 132320
rect 138868 132280 138870 132320
rect 139032 132280 139041 132320
rect 138655 132238 138702 132280
rect 138826 132238 138870 132280
rect 138994 132238 139041 132280
rect 79415 131564 79462 131606
rect 79586 131564 79630 131606
rect 79754 131564 79801 131606
rect 79415 131524 79424 131564
rect 79586 131524 79588 131564
rect 79628 131524 79630 131564
rect 79792 131524 79801 131564
rect 79415 131482 79462 131524
rect 79586 131482 79630 131524
rect 79754 131482 79801 131524
rect 94535 131564 94582 131606
rect 94706 131564 94750 131606
rect 94874 131564 94921 131606
rect 94535 131524 94544 131564
rect 94706 131524 94708 131564
rect 94748 131524 94750 131564
rect 94912 131524 94921 131564
rect 94535 131482 94582 131524
rect 94706 131482 94750 131524
rect 94874 131482 94921 131524
rect 109655 131564 109702 131606
rect 109826 131564 109870 131606
rect 109994 131564 110041 131606
rect 109655 131524 109664 131564
rect 109826 131524 109828 131564
rect 109868 131524 109870 131564
rect 110032 131524 110041 131564
rect 109655 131482 109702 131524
rect 109826 131482 109870 131524
rect 109994 131482 110041 131524
rect 124775 131564 124822 131606
rect 124946 131564 124990 131606
rect 125114 131564 125161 131606
rect 124775 131524 124784 131564
rect 124946 131524 124948 131564
rect 124988 131524 124990 131564
rect 125152 131524 125161 131564
rect 124775 131482 124822 131524
rect 124946 131482 124990 131524
rect 125114 131482 125161 131524
rect 139895 131564 139942 131606
rect 140066 131564 140110 131606
rect 140234 131564 140281 131606
rect 139895 131524 139904 131564
rect 140066 131524 140068 131564
rect 140108 131524 140110 131564
rect 140272 131524 140281 131564
rect 139895 131482 139942 131524
rect 140066 131482 140110 131524
rect 140234 131482 140281 131524
rect 78175 130808 78222 130850
rect 78346 130808 78390 130850
rect 78514 130808 78561 130850
rect 78175 130768 78184 130808
rect 78346 130768 78348 130808
rect 78388 130768 78390 130808
rect 78552 130768 78561 130808
rect 78175 130726 78222 130768
rect 78346 130726 78390 130768
rect 78514 130726 78561 130768
rect 93295 130808 93342 130850
rect 93466 130808 93510 130850
rect 93634 130808 93681 130850
rect 93295 130768 93304 130808
rect 93466 130768 93468 130808
rect 93508 130768 93510 130808
rect 93672 130768 93681 130808
rect 93295 130726 93342 130768
rect 93466 130726 93510 130768
rect 93634 130726 93681 130768
rect 108415 130808 108462 130850
rect 108586 130808 108630 130850
rect 108754 130808 108801 130850
rect 108415 130768 108424 130808
rect 108586 130768 108588 130808
rect 108628 130768 108630 130808
rect 108792 130768 108801 130808
rect 108415 130726 108462 130768
rect 108586 130726 108630 130768
rect 108754 130726 108801 130768
rect 123535 130808 123582 130850
rect 123706 130808 123750 130850
rect 123874 130808 123921 130850
rect 123535 130768 123544 130808
rect 123706 130768 123708 130808
rect 123748 130768 123750 130808
rect 123912 130768 123921 130808
rect 123535 130726 123582 130768
rect 123706 130726 123750 130768
rect 123874 130726 123921 130768
rect 138655 130808 138702 130850
rect 138826 130808 138870 130850
rect 138994 130808 139041 130850
rect 138655 130768 138664 130808
rect 138826 130768 138828 130808
rect 138868 130768 138870 130808
rect 139032 130768 139041 130808
rect 138655 130726 138702 130768
rect 138826 130726 138870 130768
rect 138994 130726 139041 130768
rect 79415 130052 79462 130094
rect 79586 130052 79630 130094
rect 79754 130052 79801 130094
rect 79415 130012 79424 130052
rect 79586 130012 79588 130052
rect 79628 130012 79630 130052
rect 79792 130012 79801 130052
rect 79415 129970 79462 130012
rect 79586 129970 79630 130012
rect 79754 129970 79801 130012
rect 94535 130052 94582 130094
rect 94706 130052 94750 130094
rect 94874 130052 94921 130094
rect 94535 130012 94544 130052
rect 94706 130012 94708 130052
rect 94748 130012 94750 130052
rect 94912 130012 94921 130052
rect 94535 129970 94582 130012
rect 94706 129970 94750 130012
rect 94874 129970 94921 130012
rect 109655 130052 109702 130094
rect 109826 130052 109870 130094
rect 109994 130052 110041 130094
rect 109655 130012 109664 130052
rect 109826 130012 109828 130052
rect 109868 130012 109870 130052
rect 110032 130012 110041 130052
rect 109655 129970 109702 130012
rect 109826 129970 109870 130012
rect 109994 129970 110041 130012
rect 124775 130052 124822 130094
rect 124946 130052 124990 130094
rect 125114 130052 125161 130094
rect 124775 130012 124784 130052
rect 124946 130012 124948 130052
rect 124988 130012 124990 130052
rect 125152 130012 125161 130052
rect 124775 129970 124822 130012
rect 124946 129970 124990 130012
rect 125114 129970 125161 130012
rect 139895 130052 139942 130094
rect 140066 130052 140110 130094
rect 140234 130052 140281 130094
rect 139895 130012 139904 130052
rect 140066 130012 140068 130052
rect 140108 130012 140110 130052
rect 140272 130012 140281 130052
rect 139895 129970 139942 130012
rect 140066 129970 140110 130012
rect 140234 129970 140281 130012
rect 78175 129296 78222 129338
rect 78346 129296 78390 129338
rect 78514 129296 78561 129338
rect 78175 129256 78184 129296
rect 78346 129256 78348 129296
rect 78388 129256 78390 129296
rect 78552 129256 78561 129296
rect 78175 129214 78222 129256
rect 78346 129214 78390 129256
rect 78514 129214 78561 129256
rect 93295 129296 93342 129338
rect 93466 129296 93510 129338
rect 93634 129296 93681 129338
rect 93295 129256 93304 129296
rect 93466 129256 93468 129296
rect 93508 129256 93510 129296
rect 93672 129256 93681 129296
rect 93295 129214 93342 129256
rect 93466 129214 93510 129256
rect 93634 129214 93681 129256
rect 108415 129296 108462 129338
rect 108586 129296 108630 129338
rect 108754 129296 108801 129338
rect 108415 129256 108424 129296
rect 108586 129256 108588 129296
rect 108628 129256 108630 129296
rect 108792 129256 108801 129296
rect 108415 129214 108462 129256
rect 108586 129214 108630 129256
rect 108754 129214 108801 129256
rect 123535 129296 123582 129338
rect 123706 129296 123750 129338
rect 123874 129296 123921 129338
rect 123535 129256 123544 129296
rect 123706 129256 123708 129296
rect 123748 129256 123750 129296
rect 123912 129256 123921 129296
rect 123535 129214 123582 129256
rect 123706 129214 123750 129256
rect 123874 129214 123921 129256
rect 138655 129296 138702 129338
rect 138826 129296 138870 129338
rect 138994 129296 139041 129338
rect 138655 129256 138664 129296
rect 138826 129256 138828 129296
rect 138868 129256 138870 129296
rect 139032 129256 139041 129296
rect 138655 129214 138702 129256
rect 138826 129214 138870 129256
rect 138994 129214 139041 129256
rect 79415 128540 79462 128582
rect 79586 128540 79630 128582
rect 79754 128540 79801 128582
rect 79415 128500 79424 128540
rect 79586 128500 79588 128540
rect 79628 128500 79630 128540
rect 79792 128500 79801 128540
rect 79415 128458 79462 128500
rect 79586 128458 79630 128500
rect 79754 128458 79801 128500
rect 94535 128540 94582 128582
rect 94706 128540 94750 128582
rect 94874 128540 94921 128582
rect 94535 128500 94544 128540
rect 94706 128500 94708 128540
rect 94748 128500 94750 128540
rect 94912 128500 94921 128540
rect 94535 128458 94582 128500
rect 94706 128458 94750 128500
rect 94874 128458 94921 128500
rect 109655 128540 109702 128582
rect 109826 128540 109870 128582
rect 109994 128540 110041 128582
rect 109655 128500 109664 128540
rect 109826 128500 109828 128540
rect 109868 128500 109870 128540
rect 110032 128500 110041 128540
rect 109655 128458 109702 128500
rect 109826 128458 109870 128500
rect 109994 128458 110041 128500
rect 124775 128540 124822 128582
rect 124946 128540 124990 128582
rect 125114 128540 125161 128582
rect 124775 128500 124784 128540
rect 124946 128500 124948 128540
rect 124988 128500 124990 128540
rect 125152 128500 125161 128540
rect 124775 128458 124822 128500
rect 124946 128458 124990 128500
rect 125114 128458 125161 128500
rect 139895 128540 139942 128582
rect 140066 128540 140110 128582
rect 140234 128540 140281 128582
rect 139895 128500 139904 128540
rect 140066 128500 140068 128540
rect 140108 128500 140110 128540
rect 140272 128500 140281 128540
rect 139895 128458 139942 128500
rect 140066 128458 140110 128500
rect 140234 128458 140281 128500
rect 78175 127784 78222 127826
rect 78346 127784 78390 127826
rect 78514 127784 78561 127826
rect 78175 127744 78184 127784
rect 78346 127744 78348 127784
rect 78388 127744 78390 127784
rect 78552 127744 78561 127784
rect 78175 127702 78222 127744
rect 78346 127702 78390 127744
rect 78514 127702 78561 127744
rect 93295 127784 93342 127826
rect 93466 127784 93510 127826
rect 93634 127784 93681 127826
rect 93295 127744 93304 127784
rect 93466 127744 93468 127784
rect 93508 127744 93510 127784
rect 93672 127744 93681 127784
rect 93295 127702 93342 127744
rect 93466 127702 93510 127744
rect 93634 127702 93681 127744
rect 108415 127784 108462 127826
rect 108586 127784 108630 127826
rect 108754 127784 108801 127826
rect 108415 127744 108424 127784
rect 108586 127744 108588 127784
rect 108628 127744 108630 127784
rect 108792 127744 108801 127784
rect 108415 127702 108462 127744
rect 108586 127702 108630 127744
rect 108754 127702 108801 127744
rect 123535 127784 123582 127826
rect 123706 127784 123750 127826
rect 123874 127784 123921 127826
rect 123535 127744 123544 127784
rect 123706 127744 123708 127784
rect 123748 127744 123750 127784
rect 123912 127744 123921 127784
rect 123535 127702 123582 127744
rect 123706 127702 123750 127744
rect 123874 127702 123921 127744
rect 138655 127784 138702 127826
rect 138826 127784 138870 127826
rect 138994 127784 139041 127826
rect 138655 127744 138664 127784
rect 138826 127744 138828 127784
rect 138868 127744 138870 127784
rect 139032 127744 139041 127784
rect 138655 127702 138702 127744
rect 138826 127702 138870 127744
rect 138994 127702 139041 127744
rect 79415 127028 79462 127070
rect 79586 127028 79630 127070
rect 79754 127028 79801 127070
rect 79415 126988 79424 127028
rect 79586 126988 79588 127028
rect 79628 126988 79630 127028
rect 79792 126988 79801 127028
rect 79415 126946 79462 126988
rect 79586 126946 79630 126988
rect 79754 126946 79801 126988
rect 94535 127028 94582 127070
rect 94706 127028 94750 127070
rect 94874 127028 94921 127070
rect 94535 126988 94544 127028
rect 94706 126988 94708 127028
rect 94748 126988 94750 127028
rect 94912 126988 94921 127028
rect 94535 126946 94582 126988
rect 94706 126946 94750 126988
rect 94874 126946 94921 126988
rect 109655 127028 109702 127070
rect 109826 127028 109870 127070
rect 109994 127028 110041 127070
rect 109655 126988 109664 127028
rect 109826 126988 109828 127028
rect 109868 126988 109870 127028
rect 110032 126988 110041 127028
rect 109655 126946 109702 126988
rect 109826 126946 109870 126988
rect 109994 126946 110041 126988
rect 124775 127028 124822 127070
rect 124946 127028 124990 127070
rect 125114 127028 125161 127070
rect 124775 126988 124784 127028
rect 124946 126988 124948 127028
rect 124988 126988 124990 127028
rect 125152 126988 125161 127028
rect 124775 126946 124822 126988
rect 124946 126946 124990 126988
rect 125114 126946 125161 126988
rect 139895 127028 139942 127070
rect 140066 127028 140110 127070
rect 140234 127028 140281 127070
rect 139895 126988 139904 127028
rect 140066 126988 140068 127028
rect 140108 126988 140110 127028
rect 140272 126988 140281 127028
rect 139895 126946 139942 126988
rect 140066 126946 140110 126988
rect 140234 126946 140281 126988
rect 78175 126272 78222 126314
rect 78346 126272 78390 126314
rect 78514 126272 78561 126314
rect 78175 126232 78184 126272
rect 78346 126232 78348 126272
rect 78388 126232 78390 126272
rect 78552 126232 78561 126272
rect 78175 126190 78222 126232
rect 78346 126190 78390 126232
rect 78514 126190 78561 126232
rect 93295 126272 93342 126314
rect 93466 126272 93510 126314
rect 93634 126272 93681 126314
rect 93295 126232 93304 126272
rect 93466 126232 93468 126272
rect 93508 126232 93510 126272
rect 93672 126232 93681 126272
rect 93295 126190 93342 126232
rect 93466 126190 93510 126232
rect 93634 126190 93681 126232
rect 108415 126272 108462 126314
rect 108586 126272 108630 126314
rect 108754 126272 108801 126314
rect 108415 126232 108424 126272
rect 108586 126232 108588 126272
rect 108628 126232 108630 126272
rect 108792 126232 108801 126272
rect 108415 126190 108462 126232
rect 108586 126190 108630 126232
rect 108754 126190 108801 126232
rect 123535 126272 123582 126314
rect 123706 126272 123750 126314
rect 123874 126272 123921 126314
rect 123535 126232 123544 126272
rect 123706 126232 123708 126272
rect 123748 126232 123750 126272
rect 123912 126232 123921 126272
rect 123535 126190 123582 126232
rect 123706 126190 123750 126232
rect 123874 126190 123921 126232
rect 138655 126272 138702 126314
rect 138826 126272 138870 126314
rect 138994 126272 139041 126314
rect 138655 126232 138664 126272
rect 138826 126232 138828 126272
rect 138868 126232 138870 126272
rect 139032 126232 139041 126272
rect 138655 126190 138702 126232
rect 138826 126190 138870 126232
rect 138994 126190 139041 126232
rect 79415 125516 79462 125558
rect 79586 125516 79630 125558
rect 79754 125516 79801 125558
rect 79415 125476 79424 125516
rect 79586 125476 79588 125516
rect 79628 125476 79630 125516
rect 79792 125476 79801 125516
rect 79415 125434 79462 125476
rect 79586 125434 79630 125476
rect 79754 125434 79801 125476
rect 94535 125516 94582 125558
rect 94706 125516 94750 125558
rect 94874 125516 94921 125558
rect 94535 125476 94544 125516
rect 94706 125476 94708 125516
rect 94748 125476 94750 125516
rect 94912 125476 94921 125516
rect 94535 125434 94582 125476
rect 94706 125434 94750 125476
rect 94874 125434 94921 125476
rect 109655 125516 109702 125558
rect 109826 125516 109870 125558
rect 109994 125516 110041 125558
rect 109655 125476 109664 125516
rect 109826 125476 109828 125516
rect 109868 125476 109870 125516
rect 110032 125476 110041 125516
rect 109655 125434 109702 125476
rect 109826 125434 109870 125476
rect 109994 125434 110041 125476
rect 124775 125516 124822 125558
rect 124946 125516 124990 125558
rect 125114 125516 125161 125558
rect 124775 125476 124784 125516
rect 124946 125476 124948 125516
rect 124988 125476 124990 125516
rect 125152 125476 125161 125516
rect 124775 125434 124822 125476
rect 124946 125434 124990 125476
rect 125114 125434 125161 125476
rect 139895 125516 139942 125558
rect 140066 125516 140110 125558
rect 140234 125516 140281 125558
rect 139895 125476 139904 125516
rect 140066 125476 140068 125516
rect 140108 125476 140110 125516
rect 140272 125476 140281 125516
rect 139895 125434 139942 125476
rect 140066 125434 140110 125476
rect 140234 125434 140281 125476
rect 78175 124760 78222 124802
rect 78346 124760 78390 124802
rect 78514 124760 78561 124802
rect 78175 124720 78184 124760
rect 78346 124720 78348 124760
rect 78388 124720 78390 124760
rect 78552 124720 78561 124760
rect 78175 124678 78222 124720
rect 78346 124678 78390 124720
rect 78514 124678 78561 124720
rect 93295 124760 93342 124802
rect 93466 124760 93510 124802
rect 93634 124760 93681 124802
rect 93295 124720 93304 124760
rect 93466 124720 93468 124760
rect 93508 124720 93510 124760
rect 93672 124720 93681 124760
rect 93295 124678 93342 124720
rect 93466 124678 93510 124720
rect 93634 124678 93681 124720
rect 108415 124760 108462 124802
rect 108586 124760 108630 124802
rect 108754 124760 108801 124802
rect 108415 124720 108424 124760
rect 108586 124720 108588 124760
rect 108628 124720 108630 124760
rect 108792 124720 108801 124760
rect 108415 124678 108462 124720
rect 108586 124678 108630 124720
rect 108754 124678 108801 124720
rect 123535 124760 123582 124802
rect 123706 124760 123750 124802
rect 123874 124760 123921 124802
rect 123535 124720 123544 124760
rect 123706 124720 123708 124760
rect 123748 124720 123750 124760
rect 123912 124720 123921 124760
rect 123535 124678 123582 124720
rect 123706 124678 123750 124720
rect 123874 124678 123921 124720
rect 138655 124760 138702 124802
rect 138826 124760 138870 124802
rect 138994 124760 139041 124802
rect 138655 124720 138664 124760
rect 138826 124720 138828 124760
rect 138868 124720 138870 124760
rect 139032 124720 139041 124760
rect 138655 124678 138702 124720
rect 138826 124678 138870 124720
rect 138994 124678 139041 124720
rect 79415 124004 79462 124046
rect 79586 124004 79630 124046
rect 79754 124004 79801 124046
rect 79415 123964 79424 124004
rect 79586 123964 79588 124004
rect 79628 123964 79630 124004
rect 79792 123964 79801 124004
rect 79415 123922 79462 123964
rect 79586 123922 79630 123964
rect 79754 123922 79801 123964
rect 94535 124004 94582 124046
rect 94706 124004 94750 124046
rect 94874 124004 94921 124046
rect 94535 123964 94544 124004
rect 94706 123964 94708 124004
rect 94748 123964 94750 124004
rect 94912 123964 94921 124004
rect 94535 123922 94582 123964
rect 94706 123922 94750 123964
rect 94874 123922 94921 123964
rect 109655 124004 109702 124046
rect 109826 124004 109870 124046
rect 109994 124004 110041 124046
rect 109655 123964 109664 124004
rect 109826 123964 109828 124004
rect 109868 123964 109870 124004
rect 110032 123964 110041 124004
rect 109655 123922 109702 123964
rect 109826 123922 109870 123964
rect 109994 123922 110041 123964
rect 124775 124004 124822 124046
rect 124946 124004 124990 124046
rect 125114 124004 125161 124046
rect 124775 123964 124784 124004
rect 124946 123964 124948 124004
rect 124988 123964 124990 124004
rect 125152 123964 125161 124004
rect 124775 123922 124822 123964
rect 124946 123922 124990 123964
rect 125114 123922 125161 123964
rect 139895 124004 139942 124046
rect 140066 124004 140110 124046
rect 140234 124004 140281 124046
rect 139895 123964 139904 124004
rect 140066 123964 140068 124004
rect 140108 123964 140110 124004
rect 140272 123964 140281 124004
rect 139895 123922 139942 123964
rect 140066 123922 140110 123964
rect 140234 123922 140281 123964
rect 78175 123248 78222 123290
rect 78346 123248 78390 123290
rect 78514 123248 78561 123290
rect 78175 123208 78184 123248
rect 78346 123208 78348 123248
rect 78388 123208 78390 123248
rect 78552 123208 78561 123248
rect 78175 123166 78222 123208
rect 78346 123166 78390 123208
rect 78514 123166 78561 123208
rect 93295 123248 93342 123290
rect 93466 123248 93510 123290
rect 93634 123248 93681 123290
rect 93295 123208 93304 123248
rect 93466 123208 93468 123248
rect 93508 123208 93510 123248
rect 93672 123208 93681 123248
rect 93295 123166 93342 123208
rect 93466 123166 93510 123208
rect 93634 123166 93681 123208
rect 108415 123248 108462 123290
rect 108586 123248 108630 123290
rect 108754 123248 108801 123290
rect 108415 123208 108424 123248
rect 108586 123208 108588 123248
rect 108628 123208 108630 123248
rect 108792 123208 108801 123248
rect 108415 123166 108462 123208
rect 108586 123166 108630 123208
rect 108754 123166 108801 123208
rect 123535 123248 123582 123290
rect 123706 123248 123750 123290
rect 123874 123248 123921 123290
rect 123535 123208 123544 123248
rect 123706 123208 123708 123248
rect 123748 123208 123750 123248
rect 123912 123208 123921 123248
rect 123535 123166 123582 123208
rect 123706 123166 123750 123208
rect 123874 123166 123921 123208
rect 138655 123248 138702 123290
rect 138826 123248 138870 123290
rect 138994 123248 139041 123290
rect 138655 123208 138664 123248
rect 138826 123208 138828 123248
rect 138868 123208 138870 123248
rect 139032 123208 139041 123248
rect 138655 123166 138702 123208
rect 138826 123166 138870 123208
rect 138994 123166 139041 123208
rect 79415 122492 79462 122534
rect 79586 122492 79630 122534
rect 79754 122492 79801 122534
rect 79415 122452 79424 122492
rect 79586 122452 79588 122492
rect 79628 122452 79630 122492
rect 79792 122452 79801 122492
rect 79415 122410 79462 122452
rect 79586 122410 79630 122452
rect 79754 122410 79801 122452
rect 94535 122492 94582 122534
rect 94706 122492 94750 122534
rect 94874 122492 94921 122534
rect 94535 122452 94544 122492
rect 94706 122452 94708 122492
rect 94748 122452 94750 122492
rect 94912 122452 94921 122492
rect 94535 122410 94582 122452
rect 94706 122410 94750 122452
rect 94874 122410 94921 122452
rect 109655 122492 109702 122534
rect 109826 122492 109870 122534
rect 109994 122492 110041 122534
rect 109655 122452 109664 122492
rect 109826 122452 109828 122492
rect 109868 122452 109870 122492
rect 110032 122452 110041 122492
rect 109655 122410 109702 122452
rect 109826 122410 109870 122452
rect 109994 122410 110041 122452
rect 124775 122492 124822 122534
rect 124946 122492 124990 122534
rect 125114 122492 125161 122534
rect 124775 122452 124784 122492
rect 124946 122452 124948 122492
rect 124988 122452 124990 122492
rect 125152 122452 125161 122492
rect 124775 122410 124822 122452
rect 124946 122410 124990 122452
rect 125114 122410 125161 122452
rect 139895 122492 139942 122534
rect 140066 122492 140110 122534
rect 140234 122492 140281 122534
rect 139895 122452 139904 122492
rect 140066 122452 140068 122492
rect 140108 122452 140110 122492
rect 140272 122452 140281 122492
rect 139895 122410 139942 122452
rect 140066 122410 140110 122452
rect 140234 122410 140281 122452
rect 78175 121736 78222 121778
rect 78346 121736 78390 121778
rect 78514 121736 78561 121778
rect 78175 121696 78184 121736
rect 78346 121696 78348 121736
rect 78388 121696 78390 121736
rect 78552 121696 78561 121736
rect 78175 121654 78222 121696
rect 78346 121654 78390 121696
rect 78514 121654 78561 121696
rect 93295 121736 93342 121778
rect 93466 121736 93510 121778
rect 93634 121736 93681 121778
rect 93295 121696 93304 121736
rect 93466 121696 93468 121736
rect 93508 121696 93510 121736
rect 93672 121696 93681 121736
rect 93295 121654 93342 121696
rect 93466 121654 93510 121696
rect 93634 121654 93681 121696
rect 108415 121736 108462 121778
rect 108586 121736 108630 121778
rect 108754 121736 108801 121778
rect 108415 121696 108424 121736
rect 108586 121696 108588 121736
rect 108628 121696 108630 121736
rect 108792 121696 108801 121736
rect 108415 121654 108462 121696
rect 108586 121654 108630 121696
rect 108754 121654 108801 121696
rect 123535 121736 123582 121778
rect 123706 121736 123750 121778
rect 123874 121736 123921 121778
rect 123535 121696 123544 121736
rect 123706 121696 123708 121736
rect 123748 121696 123750 121736
rect 123912 121696 123921 121736
rect 123535 121654 123582 121696
rect 123706 121654 123750 121696
rect 123874 121654 123921 121696
rect 138655 121736 138702 121778
rect 138826 121736 138870 121778
rect 138994 121736 139041 121778
rect 138655 121696 138664 121736
rect 138826 121696 138828 121736
rect 138868 121696 138870 121736
rect 139032 121696 139041 121736
rect 138655 121654 138702 121696
rect 138826 121654 138870 121696
rect 138994 121654 139041 121696
rect 79415 120980 79462 121022
rect 79586 120980 79630 121022
rect 79754 120980 79801 121022
rect 79415 120940 79424 120980
rect 79586 120940 79588 120980
rect 79628 120940 79630 120980
rect 79792 120940 79801 120980
rect 79415 120898 79462 120940
rect 79586 120898 79630 120940
rect 79754 120898 79801 120940
rect 94535 120980 94582 121022
rect 94706 120980 94750 121022
rect 94874 120980 94921 121022
rect 94535 120940 94544 120980
rect 94706 120940 94708 120980
rect 94748 120940 94750 120980
rect 94912 120940 94921 120980
rect 94535 120898 94582 120940
rect 94706 120898 94750 120940
rect 94874 120898 94921 120940
rect 109655 120980 109702 121022
rect 109826 120980 109870 121022
rect 109994 120980 110041 121022
rect 109655 120940 109664 120980
rect 109826 120940 109828 120980
rect 109868 120940 109870 120980
rect 110032 120940 110041 120980
rect 109655 120898 109702 120940
rect 109826 120898 109870 120940
rect 109994 120898 110041 120940
rect 124775 120980 124822 121022
rect 124946 120980 124990 121022
rect 125114 120980 125161 121022
rect 124775 120940 124784 120980
rect 124946 120940 124948 120980
rect 124988 120940 124990 120980
rect 125152 120940 125161 120980
rect 124775 120898 124822 120940
rect 124946 120898 124990 120940
rect 125114 120898 125161 120940
rect 139895 120980 139942 121022
rect 140066 120980 140110 121022
rect 140234 120980 140281 121022
rect 139895 120940 139904 120980
rect 140066 120940 140068 120980
rect 140108 120940 140110 120980
rect 140272 120940 140281 120980
rect 139895 120898 139942 120940
rect 140066 120898 140110 120940
rect 140234 120898 140281 120940
rect 78175 120224 78222 120266
rect 78346 120224 78390 120266
rect 78514 120224 78561 120266
rect 78175 120184 78184 120224
rect 78346 120184 78348 120224
rect 78388 120184 78390 120224
rect 78552 120184 78561 120224
rect 78175 120142 78222 120184
rect 78346 120142 78390 120184
rect 78514 120142 78561 120184
rect 93295 120224 93342 120266
rect 93466 120224 93510 120266
rect 93634 120224 93681 120266
rect 93295 120184 93304 120224
rect 93466 120184 93468 120224
rect 93508 120184 93510 120224
rect 93672 120184 93681 120224
rect 93295 120142 93342 120184
rect 93466 120142 93510 120184
rect 93634 120142 93681 120184
rect 108415 120224 108462 120266
rect 108586 120224 108630 120266
rect 108754 120224 108801 120266
rect 108415 120184 108424 120224
rect 108586 120184 108588 120224
rect 108628 120184 108630 120224
rect 108792 120184 108801 120224
rect 108415 120142 108462 120184
rect 108586 120142 108630 120184
rect 108754 120142 108801 120184
rect 123535 120224 123582 120266
rect 123706 120224 123750 120266
rect 123874 120224 123921 120266
rect 123535 120184 123544 120224
rect 123706 120184 123708 120224
rect 123748 120184 123750 120224
rect 123912 120184 123921 120224
rect 123535 120142 123582 120184
rect 123706 120142 123750 120184
rect 123874 120142 123921 120184
rect 138655 120224 138702 120266
rect 138826 120224 138870 120266
rect 138994 120224 139041 120266
rect 138655 120184 138664 120224
rect 138826 120184 138828 120224
rect 138868 120184 138870 120224
rect 139032 120184 139041 120224
rect 138655 120142 138702 120184
rect 138826 120142 138870 120184
rect 138994 120142 139041 120184
rect 79415 119468 79462 119510
rect 79586 119468 79630 119510
rect 79754 119468 79801 119510
rect 79415 119428 79424 119468
rect 79586 119428 79588 119468
rect 79628 119428 79630 119468
rect 79792 119428 79801 119468
rect 79415 119386 79462 119428
rect 79586 119386 79630 119428
rect 79754 119386 79801 119428
rect 94535 119468 94582 119510
rect 94706 119468 94750 119510
rect 94874 119468 94921 119510
rect 94535 119428 94544 119468
rect 94706 119428 94708 119468
rect 94748 119428 94750 119468
rect 94912 119428 94921 119468
rect 94535 119386 94582 119428
rect 94706 119386 94750 119428
rect 94874 119386 94921 119428
rect 109655 119468 109702 119510
rect 109826 119468 109870 119510
rect 109994 119468 110041 119510
rect 109655 119428 109664 119468
rect 109826 119428 109828 119468
rect 109868 119428 109870 119468
rect 110032 119428 110041 119468
rect 109655 119386 109702 119428
rect 109826 119386 109870 119428
rect 109994 119386 110041 119428
rect 124775 119468 124822 119510
rect 124946 119468 124990 119510
rect 125114 119468 125161 119510
rect 124775 119428 124784 119468
rect 124946 119428 124948 119468
rect 124988 119428 124990 119468
rect 125152 119428 125161 119468
rect 124775 119386 124822 119428
rect 124946 119386 124990 119428
rect 125114 119386 125161 119428
rect 139895 119468 139942 119510
rect 140066 119468 140110 119510
rect 140234 119468 140281 119510
rect 139895 119428 139904 119468
rect 140066 119428 140068 119468
rect 140108 119428 140110 119468
rect 140272 119428 140281 119468
rect 139895 119386 139942 119428
rect 140066 119386 140110 119428
rect 140234 119386 140281 119428
rect 78175 118712 78222 118754
rect 78346 118712 78390 118754
rect 78514 118712 78561 118754
rect 78175 118672 78184 118712
rect 78346 118672 78348 118712
rect 78388 118672 78390 118712
rect 78552 118672 78561 118712
rect 78175 118630 78222 118672
rect 78346 118630 78390 118672
rect 78514 118630 78561 118672
rect 93295 118712 93342 118754
rect 93466 118712 93510 118754
rect 93634 118712 93681 118754
rect 93295 118672 93304 118712
rect 93466 118672 93468 118712
rect 93508 118672 93510 118712
rect 93672 118672 93681 118712
rect 93295 118630 93342 118672
rect 93466 118630 93510 118672
rect 93634 118630 93681 118672
rect 108415 118712 108462 118754
rect 108586 118712 108630 118754
rect 108754 118712 108801 118754
rect 108415 118672 108424 118712
rect 108586 118672 108588 118712
rect 108628 118672 108630 118712
rect 108792 118672 108801 118712
rect 108415 118630 108462 118672
rect 108586 118630 108630 118672
rect 108754 118630 108801 118672
rect 123535 118712 123582 118754
rect 123706 118712 123750 118754
rect 123874 118712 123921 118754
rect 123535 118672 123544 118712
rect 123706 118672 123708 118712
rect 123748 118672 123750 118712
rect 123912 118672 123921 118712
rect 123535 118630 123582 118672
rect 123706 118630 123750 118672
rect 123874 118630 123921 118672
rect 138655 118712 138702 118754
rect 138826 118712 138870 118754
rect 138994 118712 139041 118754
rect 138655 118672 138664 118712
rect 138826 118672 138828 118712
rect 138868 118672 138870 118712
rect 139032 118672 139041 118712
rect 138655 118630 138702 118672
rect 138826 118630 138870 118672
rect 138994 118630 139041 118672
rect 79415 117956 79462 117998
rect 79586 117956 79630 117998
rect 79754 117956 79801 117998
rect 79415 117916 79424 117956
rect 79586 117916 79588 117956
rect 79628 117916 79630 117956
rect 79792 117916 79801 117956
rect 79415 117874 79462 117916
rect 79586 117874 79630 117916
rect 79754 117874 79801 117916
rect 94535 117956 94582 117998
rect 94706 117956 94750 117998
rect 94874 117956 94921 117998
rect 94535 117916 94544 117956
rect 94706 117916 94708 117956
rect 94748 117916 94750 117956
rect 94912 117916 94921 117956
rect 94535 117874 94582 117916
rect 94706 117874 94750 117916
rect 94874 117874 94921 117916
rect 109655 117956 109702 117998
rect 109826 117956 109870 117998
rect 109994 117956 110041 117998
rect 109655 117916 109664 117956
rect 109826 117916 109828 117956
rect 109868 117916 109870 117956
rect 110032 117916 110041 117956
rect 109655 117874 109702 117916
rect 109826 117874 109870 117916
rect 109994 117874 110041 117916
rect 124775 117956 124822 117998
rect 124946 117956 124990 117998
rect 125114 117956 125161 117998
rect 124775 117916 124784 117956
rect 124946 117916 124948 117956
rect 124988 117916 124990 117956
rect 125152 117916 125161 117956
rect 124775 117874 124822 117916
rect 124946 117874 124990 117916
rect 125114 117874 125161 117916
rect 139895 117956 139942 117998
rect 140066 117956 140110 117998
rect 140234 117956 140281 117998
rect 139895 117916 139904 117956
rect 140066 117916 140068 117956
rect 140108 117916 140110 117956
rect 140272 117916 140281 117956
rect 139895 117874 139942 117916
rect 140066 117874 140110 117916
rect 140234 117874 140281 117916
rect 78175 117200 78222 117242
rect 78346 117200 78390 117242
rect 78514 117200 78561 117242
rect 78175 117160 78184 117200
rect 78346 117160 78348 117200
rect 78388 117160 78390 117200
rect 78552 117160 78561 117200
rect 78175 117118 78222 117160
rect 78346 117118 78390 117160
rect 78514 117118 78561 117160
rect 93295 117200 93342 117242
rect 93466 117200 93510 117242
rect 93634 117200 93681 117242
rect 93295 117160 93304 117200
rect 93466 117160 93468 117200
rect 93508 117160 93510 117200
rect 93672 117160 93681 117200
rect 93295 117118 93342 117160
rect 93466 117118 93510 117160
rect 93634 117118 93681 117160
rect 108415 117200 108462 117242
rect 108586 117200 108630 117242
rect 108754 117200 108801 117242
rect 108415 117160 108424 117200
rect 108586 117160 108588 117200
rect 108628 117160 108630 117200
rect 108792 117160 108801 117200
rect 108415 117118 108462 117160
rect 108586 117118 108630 117160
rect 108754 117118 108801 117160
rect 123535 117200 123582 117242
rect 123706 117200 123750 117242
rect 123874 117200 123921 117242
rect 123535 117160 123544 117200
rect 123706 117160 123708 117200
rect 123748 117160 123750 117200
rect 123912 117160 123921 117200
rect 123535 117118 123582 117160
rect 123706 117118 123750 117160
rect 123874 117118 123921 117160
rect 138655 117200 138702 117242
rect 138826 117200 138870 117242
rect 138994 117200 139041 117242
rect 138655 117160 138664 117200
rect 138826 117160 138828 117200
rect 138868 117160 138870 117200
rect 139032 117160 139041 117200
rect 138655 117118 138702 117160
rect 138826 117118 138870 117160
rect 138994 117118 139041 117160
rect 79415 116444 79462 116486
rect 79586 116444 79630 116486
rect 79754 116444 79801 116486
rect 79415 116404 79424 116444
rect 79586 116404 79588 116444
rect 79628 116404 79630 116444
rect 79792 116404 79801 116444
rect 79415 116362 79462 116404
rect 79586 116362 79630 116404
rect 79754 116362 79801 116404
rect 94535 116444 94582 116486
rect 94706 116444 94750 116486
rect 94874 116444 94921 116486
rect 94535 116404 94544 116444
rect 94706 116404 94708 116444
rect 94748 116404 94750 116444
rect 94912 116404 94921 116444
rect 94535 116362 94582 116404
rect 94706 116362 94750 116404
rect 94874 116362 94921 116404
rect 109655 116444 109702 116486
rect 109826 116444 109870 116486
rect 109994 116444 110041 116486
rect 109655 116404 109664 116444
rect 109826 116404 109828 116444
rect 109868 116404 109870 116444
rect 110032 116404 110041 116444
rect 109655 116362 109702 116404
rect 109826 116362 109870 116404
rect 109994 116362 110041 116404
rect 124775 116444 124822 116486
rect 124946 116444 124990 116486
rect 125114 116444 125161 116486
rect 124775 116404 124784 116444
rect 124946 116404 124948 116444
rect 124988 116404 124990 116444
rect 125152 116404 125161 116444
rect 124775 116362 124822 116404
rect 124946 116362 124990 116404
rect 125114 116362 125161 116404
rect 139895 116444 139942 116486
rect 140066 116444 140110 116486
rect 140234 116444 140281 116486
rect 139895 116404 139904 116444
rect 140066 116404 140068 116444
rect 140108 116404 140110 116444
rect 140272 116404 140281 116444
rect 139895 116362 139942 116404
rect 140066 116362 140110 116404
rect 140234 116362 140281 116404
rect 78175 115688 78222 115730
rect 78346 115688 78390 115730
rect 78514 115688 78561 115730
rect 78175 115648 78184 115688
rect 78346 115648 78348 115688
rect 78388 115648 78390 115688
rect 78552 115648 78561 115688
rect 78175 115606 78222 115648
rect 78346 115606 78390 115648
rect 78514 115606 78561 115648
rect 93295 115688 93342 115730
rect 93466 115688 93510 115730
rect 93634 115688 93681 115730
rect 93295 115648 93304 115688
rect 93466 115648 93468 115688
rect 93508 115648 93510 115688
rect 93672 115648 93681 115688
rect 93295 115606 93342 115648
rect 93466 115606 93510 115648
rect 93634 115606 93681 115648
rect 108415 115688 108462 115730
rect 108586 115688 108630 115730
rect 108754 115688 108801 115730
rect 108415 115648 108424 115688
rect 108586 115648 108588 115688
rect 108628 115648 108630 115688
rect 108792 115648 108801 115688
rect 108415 115606 108462 115648
rect 108586 115606 108630 115648
rect 108754 115606 108801 115648
rect 123535 115688 123582 115730
rect 123706 115688 123750 115730
rect 123874 115688 123921 115730
rect 123535 115648 123544 115688
rect 123706 115648 123708 115688
rect 123748 115648 123750 115688
rect 123912 115648 123921 115688
rect 123535 115606 123582 115648
rect 123706 115606 123750 115648
rect 123874 115606 123921 115648
rect 138655 115688 138702 115730
rect 138826 115688 138870 115730
rect 138994 115688 139041 115730
rect 138655 115648 138664 115688
rect 138826 115648 138828 115688
rect 138868 115648 138870 115688
rect 139032 115648 139041 115688
rect 138655 115606 138702 115648
rect 138826 115606 138870 115648
rect 138994 115606 139041 115648
rect 79415 114932 79462 114974
rect 79586 114932 79630 114974
rect 79754 114932 79801 114974
rect 79415 114892 79424 114932
rect 79586 114892 79588 114932
rect 79628 114892 79630 114932
rect 79792 114892 79801 114932
rect 79415 114850 79462 114892
rect 79586 114850 79630 114892
rect 79754 114850 79801 114892
rect 94535 114932 94582 114974
rect 94706 114932 94750 114974
rect 94874 114932 94921 114974
rect 94535 114892 94544 114932
rect 94706 114892 94708 114932
rect 94748 114892 94750 114932
rect 94912 114892 94921 114932
rect 94535 114850 94582 114892
rect 94706 114850 94750 114892
rect 94874 114850 94921 114892
rect 109655 114932 109702 114974
rect 109826 114932 109870 114974
rect 109994 114932 110041 114974
rect 109655 114892 109664 114932
rect 109826 114892 109828 114932
rect 109868 114892 109870 114932
rect 110032 114892 110041 114932
rect 109655 114850 109702 114892
rect 109826 114850 109870 114892
rect 109994 114850 110041 114892
rect 124775 114932 124822 114974
rect 124946 114932 124990 114974
rect 125114 114932 125161 114974
rect 124775 114892 124784 114932
rect 124946 114892 124948 114932
rect 124988 114892 124990 114932
rect 125152 114892 125161 114932
rect 124775 114850 124822 114892
rect 124946 114850 124990 114892
rect 125114 114850 125161 114892
rect 139895 114932 139942 114974
rect 140066 114932 140110 114974
rect 140234 114932 140281 114974
rect 139895 114892 139904 114932
rect 140066 114892 140068 114932
rect 140108 114892 140110 114932
rect 140272 114892 140281 114932
rect 139895 114850 139942 114892
rect 140066 114850 140110 114892
rect 140234 114850 140281 114892
rect 78175 114176 78222 114218
rect 78346 114176 78390 114218
rect 78514 114176 78561 114218
rect 78175 114136 78184 114176
rect 78346 114136 78348 114176
rect 78388 114136 78390 114176
rect 78552 114136 78561 114176
rect 78175 114094 78222 114136
rect 78346 114094 78390 114136
rect 78514 114094 78561 114136
rect 93295 114176 93342 114218
rect 93466 114176 93510 114218
rect 93634 114176 93681 114218
rect 93295 114136 93304 114176
rect 93466 114136 93468 114176
rect 93508 114136 93510 114176
rect 93672 114136 93681 114176
rect 93295 114094 93342 114136
rect 93466 114094 93510 114136
rect 93634 114094 93681 114136
rect 108415 114176 108462 114218
rect 108586 114176 108630 114218
rect 108754 114176 108801 114218
rect 108415 114136 108424 114176
rect 108586 114136 108588 114176
rect 108628 114136 108630 114176
rect 108792 114136 108801 114176
rect 108415 114094 108462 114136
rect 108586 114094 108630 114136
rect 108754 114094 108801 114136
rect 123535 114176 123582 114218
rect 123706 114176 123750 114218
rect 123874 114176 123921 114218
rect 123535 114136 123544 114176
rect 123706 114136 123708 114176
rect 123748 114136 123750 114176
rect 123912 114136 123921 114176
rect 123535 114094 123582 114136
rect 123706 114094 123750 114136
rect 123874 114094 123921 114136
rect 138655 114176 138702 114218
rect 138826 114176 138870 114218
rect 138994 114176 139041 114218
rect 138655 114136 138664 114176
rect 138826 114136 138828 114176
rect 138868 114136 138870 114176
rect 139032 114136 139041 114176
rect 138655 114094 138702 114136
rect 138826 114094 138870 114136
rect 138994 114094 139041 114136
rect 79415 113420 79462 113462
rect 79586 113420 79630 113462
rect 79754 113420 79801 113462
rect 79415 113380 79424 113420
rect 79586 113380 79588 113420
rect 79628 113380 79630 113420
rect 79792 113380 79801 113420
rect 79415 113338 79462 113380
rect 79586 113338 79630 113380
rect 79754 113338 79801 113380
rect 94535 113420 94582 113462
rect 94706 113420 94750 113462
rect 94874 113420 94921 113462
rect 94535 113380 94544 113420
rect 94706 113380 94708 113420
rect 94748 113380 94750 113420
rect 94912 113380 94921 113420
rect 94535 113338 94582 113380
rect 94706 113338 94750 113380
rect 94874 113338 94921 113380
rect 109655 113420 109702 113462
rect 109826 113420 109870 113462
rect 109994 113420 110041 113462
rect 109655 113380 109664 113420
rect 109826 113380 109828 113420
rect 109868 113380 109870 113420
rect 110032 113380 110041 113420
rect 109655 113338 109702 113380
rect 109826 113338 109870 113380
rect 109994 113338 110041 113380
rect 124775 113420 124822 113462
rect 124946 113420 124990 113462
rect 125114 113420 125161 113462
rect 124775 113380 124784 113420
rect 124946 113380 124948 113420
rect 124988 113380 124990 113420
rect 125152 113380 125161 113420
rect 124775 113338 124822 113380
rect 124946 113338 124990 113380
rect 125114 113338 125161 113380
rect 139895 113420 139942 113462
rect 140066 113420 140110 113462
rect 140234 113420 140281 113462
rect 139895 113380 139904 113420
rect 140066 113380 140068 113420
rect 140108 113380 140110 113420
rect 140272 113380 140281 113420
rect 139895 113338 139942 113380
rect 140066 113338 140110 113380
rect 140234 113338 140281 113380
rect 78175 112664 78222 112706
rect 78346 112664 78390 112706
rect 78514 112664 78561 112706
rect 78175 112624 78184 112664
rect 78346 112624 78348 112664
rect 78388 112624 78390 112664
rect 78552 112624 78561 112664
rect 78175 112582 78222 112624
rect 78346 112582 78390 112624
rect 78514 112582 78561 112624
rect 93295 112664 93342 112706
rect 93466 112664 93510 112706
rect 93634 112664 93681 112706
rect 93295 112624 93304 112664
rect 93466 112624 93468 112664
rect 93508 112624 93510 112664
rect 93672 112624 93681 112664
rect 93295 112582 93342 112624
rect 93466 112582 93510 112624
rect 93634 112582 93681 112624
rect 108415 112664 108462 112706
rect 108586 112664 108630 112706
rect 108754 112664 108801 112706
rect 108415 112624 108424 112664
rect 108586 112624 108588 112664
rect 108628 112624 108630 112664
rect 108792 112624 108801 112664
rect 108415 112582 108462 112624
rect 108586 112582 108630 112624
rect 108754 112582 108801 112624
rect 123535 112664 123582 112706
rect 123706 112664 123750 112706
rect 123874 112664 123921 112706
rect 123535 112624 123544 112664
rect 123706 112624 123708 112664
rect 123748 112624 123750 112664
rect 123912 112624 123921 112664
rect 123535 112582 123582 112624
rect 123706 112582 123750 112624
rect 123874 112582 123921 112624
rect 138655 112664 138702 112706
rect 138826 112664 138870 112706
rect 138994 112664 139041 112706
rect 138655 112624 138664 112664
rect 138826 112624 138828 112664
rect 138868 112624 138870 112664
rect 139032 112624 139041 112664
rect 138655 112582 138702 112624
rect 138826 112582 138870 112624
rect 138994 112582 139041 112624
rect 79415 111908 79462 111950
rect 79586 111908 79630 111950
rect 79754 111908 79801 111950
rect 79415 111868 79424 111908
rect 79586 111868 79588 111908
rect 79628 111868 79630 111908
rect 79792 111868 79801 111908
rect 79415 111826 79462 111868
rect 79586 111826 79630 111868
rect 79754 111826 79801 111868
rect 94535 111908 94582 111950
rect 94706 111908 94750 111950
rect 94874 111908 94921 111950
rect 94535 111868 94544 111908
rect 94706 111868 94708 111908
rect 94748 111868 94750 111908
rect 94912 111868 94921 111908
rect 94535 111826 94582 111868
rect 94706 111826 94750 111868
rect 94874 111826 94921 111868
rect 109655 111908 109702 111950
rect 109826 111908 109870 111950
rect 109994 111908 110041 111950
rect 109655 111868 109664 111908
rect 109826 111868 109828 111908
rect 109868 111868 109870 111908
rect 110032 111868 110041 111908
rect 109655 111826 109702 111868
rect 109826 111826 109870 111868
rect 109994 111826 110041 111868
rect 124775 111908 124822 111950
rect 124946 111908 124990 111950
rect 125114 111908 125161 111950
rect 124775 111868 124784 111908
rect 124946 111868 124948 111908
rect 124988 111868 124990 111908
rect 125152 111868 125161 111908
rect 124775 111826 124822 111868
rect 124946 111826 124990 111868
rect 125114 111826 125161 111868
rect 139895 111908 139942 111950
rect 140066 111908 140110 111950
rect 140234 111908 140281 111950
rect 139895 111868 139904 111908
rect 140066 111868 140068 111908
rect 140108 111868 140110 111908
rect 140272 111868 140281 111908
rect 139895 111826 139942 111868
rect 140066 111826 140110 111868
rect 140234 111826 140281 111868
rect 78175 111152 78222 111194
rect 78346 111152 78390 111194
rect 78514 111152 78561 111194
rect 78175 111112 78184 111152
rect 78346 111112 78348 111152
rect 78388 111112 78390 111152
rect 78552 111112 78561 111152
rect 78175 111070 78222 111112
rect 78346 111070 78390 111112
rect 78514 111070 78561 111112
rect 93295 111152 93342 111194
rect 93466 111152 93510 111194
rect 93634 111152 93681 111194
rect 93295 111112 93304 111152
rect 93466 111112 93468 111152
rect 93508 111112 93510 111152
rect 93672 111112 93681 111152
rect 93295 111070 93342 111112
rect 93466 111070 93510 111112
rect 93634 111070 93681 111112
rect 108415 111152 108462 111194
rect 108586 111152 108630 111194
rect 108754 111152 108801 111194
rect 108415 111112 108424 111152
rect 108586 111112 108588 111152
rect 108628 111112 108630 111152
rect 108792 111112 108801 111152
rect 108415 111070 108462 111112
rect 108586 111070 108630 111112
rect 108754 111070 108801 111112
rect 123535 111152 123582 111194
rect 123706 111152 123750 111194
rect 123874 111152 123921 111194
rect 123535 111112 123544 111152
rect 123706 111112 123708 111152
rect 123748 111112 123750 111152
rect 123912 111112 123921 111152
rect 123535 111070 123582 111112
rect 123706 111070 123750 111112
rect 123874 111070 123921 111112
rect 138655 111152 138702 111194
rect 138826 111152 138870 111194
rect 138994 111152 139041 111194
rect 138655 111112 138664 111152
rect 138826 111112 138828 111152
rect 138868 111112 138870 111152
rect 139032 111112 139041 111152
rect 138655 111070 138702 111112
rect 138826 111070 138870 111112
rect 138994 111070 139041 111112
rect 79415 110396 79462 110438
rect 79586 110396 79630 110438
rect 79754 110396 79801 110438
rect 79415 110356 79424 110396
rect 79586 110356 79588 110396
rect 79628 110356 79630 110396
rect 79792 110356 79801 110396
rect 79415 110314 79462 110356
rect 79586 110314 79630 110356
rect 79754 110314 79801 110356
rect 94535 110396 94582 110438
rect 94706 110396 94750 110438
rect 94874 110396 94921 110438
rect 94535 110356 94544 110396
rect 94706 110356 94708 110396
rect 94748 110356 94750 110396
rect 94912 110356 94921 110396
rect 94535 110314 94582 110356
rect 94706 110314 94750 110356
rect 94874 110314 94921 110356
rect 109655 110396 109702 110438
rect 109826 110396 109870 110438
rect 109994 110396 110041 110438
rect 109655 110356 109664 110396
rect 109826 110356 109828 110396
rect 109868 110356 109870 110396
rect 110032 110356 110041 110396
rect 109655 110314 109702 110356
rect 109826 110314 109870 110356
rect 109994 110314 110041 110356
rect 124775 110396 124822 110438
rect 124946 110396 124990 110438
rect 125114 110396 125161 110438
rect 124775 110356 124784 110396
rect 124946 110356 124948 110396
rect 124988 110356 124990 110396
rect 125152 110356 125161 110396
rect 124775 110314 124822 110356
rect 124946 110314 124990 110356
rect 125114 110314 125161 110356
rect 139895 110396 139942 110438
rect 140066 110396 140110 110438
rect 140234 110396 140281 110438
rect 139895 110356 139904 110396
rect 140066 110356 140068 110396
rect 140108 110356 140110 110396
rect 140272 110356 140281 110396
rect 139895 110314 139942 110356
rect 140066 110314 140110 110356
rect 140234 110314 140281 110356
rect 78175 109640 78222 109682
rect 78346 109640 78390 109682
rect 78514 109640 78561 109682
rect 78175 109600 78184 109640
rect 78346 109600 78348 109640
rect 78388 109600 78390 109640
rect 78552 109600 78561 109640
rect 78175 109558 78222 109600
rect 78346 109558 78390 109600
rect 78514 109558 78561 109600
rect 93295 109640 93342 109682
rect 93466 109640 93510 109682
rect 93634 109640 93681 109682
rect 93295 109600 93304 109640
rect 93466 109600 93468 109640
rect 93508 109600 93510 109640
rect 93672 109600 93681 109640
rect 93295 109558 93342 109600
rect 93466 109558 93510 109600
rect 93634 109558 93681 109600
rect 108415 109640 108462 109682
rect 108586 109640 108630 109682
rect 108754 109640 108801 109682
rect 108415 109600 108424 109640
rect 108586 109600 108588 109640
rect 108628 109600 108630 109640
rect 108792 109600 108801 109640
rect 108415 109558 108462 109600
rect 108586 109558 108630 109600
rect 108754 109558 108801 109600
rect 123535 109640 123582 109682
rect 123706 109640 123750 109682
rect 123874 109640 123921 109682
rect 123535 109600 123544 109640
rect 123706 109600 123708 109640
rect 123748 109600 123750 109640
rect 123912 109600 123921 109640
rect 123535 109558 123582 109600
rect 123706 109558 123750 109600
rect 123874 109558 123921 109600
rect 138655 109640 138702 109682
rect 138826 109640 138870 109682
rect 138994 109640 139041 109682
rect 138655 109600 138664 109640
rect 138826 109600 138828 109640
rect 138868 109600 138870 109640
rect 139032 109600 139041 109640
rect 138655 109558 138702 109600
rect 138826 109558 138870 109600
rect 138994 109558 139041 109600
rect 79415 108884 79462 108926
rect 79586 108884 79630 108926
rect 79754 108884 79801 108926
rect 79415 108844 79424 108884
rect 79586 108844 79588 108884
rect 79628 108844 79630 108884
rect 79792 108844 79801 108884
rect 79415 108802 79462 108844
rect 79586 108802 79630 108844
rect 79754 108802 79801 108844
rect 94535 108884 94582 108926
rect 94706 108884 94750 108926
rect 94874 108884 94921 108926
rect 94535 108844 94544 108884
rect 94706 108844 94708 108884
rect 94748 108844 94750 108884
rect 94912 108844 94921 108884
rect 94535 108802 94582 108844
rect 94706 108802 94750 108844
rect 94874 108802 94921 108844
rect 109655 108884 109702 108926
rect 109826 108884 109870 108926
rect 109994 108884 110041 108926
rect 109655 108844 109664 108884
rect 109826 108844 109828 108884
rect 109868 108844 109870 108884
rect 110032 108844 110041 108884
rect 109655 108802 109702 108844
rect 109826 108802 109870 108844
rect 109994 108802 110041 108844
rect 124775 108884 124822 108926
rect 124946 108884 124990 108926
rect 125114 108884 125161 108926
rect 124775 108844 124784 108884
rect 124946 108844 124948 108884
rect 124988 108844 124990 108884
rect 125152 108844 125161 108884
rect 124775 108802 124822 108844
rect 124946 108802 124990 108844
rect 125114 108802 125161 108844
rect 139895 108884 139942 108926
rect 140066 108884 140110 108926
rect 140234 108884 140281 108926
rect 139895 108844 139904 108884
rect 140066 108844 140068 108884
rect 140108 108844 140110 108884
rect 140272 108844 140281 108884
rect 139895 108802 139942 108844
rect 140066 108802 140110 108844
rect 140234 108802 140281 108844
rect 78175 108128 78222 108170
rect 78346 108128 78390 108170
rect 78514 108128 78561 108170
rect 78175 108088 78184 108128
rect 78346 108088 78348 108128
rect 78388 108088 78390 108128
rect 78552 108088 78561 108128
rect 78175 108046 78222 108088
rect 78346 108046 78390 108088
rect 78514 108046 78561 108088
rect 93295 108128 93342 108170
rect 93466 108128 93510 108170
rect 93634 108128 93681 108170
rect 93295 108088 93304 108128
rect 93466 108088 93468 108128
rect 93508 108088 93510 108128
rect 93672 108088 93681 108128
rect 93295 108046 93342 108088
rect 93466 108046 93510 108088
rect 93634 108046 93681 108088
rect 108415 108128 108462 108170
rect 108586 108128 108630 108170
rect 108754 108128 108801 108170
rect 108415 108088 108424 108128
rect 108586 108088 108588 108128
rect 108628 108088 108630 108128
rect 108792 108088 108801 108128
rect 108415 108046 108462 108088
rect 108586 108046 108630 108088
rect 108754 108046 108801 108088
rect 123535 108128 123582 108170
rect 123706 108128 123750 108170
rect 123874 108128 123921 108170
rect 123535 108088 123544 108128
rect 123706 108088 123708 108128
rect 123748 108088 123750 108128
rect 123912 108088 123921 108128
rect 123535 108046 123582 108088
rect 123706 108046 123750 108088
rect 123874 108046 123921 108088
rect 138655 108128 138702 108170
rect 138826 108128 138870 108170
rect 138994 108128 139041 108170
rect 138655 108088 138664 108128
rect 138826 108088 138828 108128
rect 138868 108088 138870 108128
rect 139032 108088 139041 108128
rect 138655 108046 138702 108088
rect 138826 108046 138870 108088
rect 138994 108046 139041 108088
rect 79415 107372 79462 107414
rect 79586 107372 79630 107414
rect 79754 107372 79801 107414
rect 79415 107332 79424 107372
rect 79586 107332 79588 107372
rect 79628 107332 79630 107372
rect 79792 107332 79801 107372
rect 79415 107290 79462 107332
rect 79586 107290 79630 107332
rect 79754 107290 79801 107332
rect 94535 107372 94582 107414
rect 94706 107372 94750 107414
rect 94874 107372 94921 107414
rect 94535 107332 94544 107372
rect 94706 107332 94708 107372
rect 94748 107332 94750 107372
rect 94912 107332 94921 107372
rect 94535 107290 94582 107332
rect 94706 107290 94750 107332
rect 94874 107290 94921 107332
rect 109655 107372 109702 107414
rect 109826 107372 109870 107414
rect 109994 107372 110041 107414
rect 109655 107332 109664 107372
rect 109826 107332 109828 107372
rect 109868 107332 109870 107372
rect 110032 107332 110041 107372
rect 109655 107290 109702 107332
rect 109826 107290 109870 107332
rect 109994 107290 110041 107332
rect 124775 107372 124822 107414
rect 124946 107372 124990 107414
rect 125114 107372 125161 107414
rect 124775 107332 124784 107372
rect 124946 107332 124948 107372
rect 124988 107332 124990 107372
rect 125152 107332 125161 107372
rect 124775 107290 124822 107332
rect 124946 107290 124990 107332
rect 125114 107290 125161 107332
rect 139895 107372 139942 107414
rect 140066 107372 140110 107414
rect 140234 107372 140281 107414
rect 139895 107332 139904 107372
rect 140066 107332 140068 107372
rect 140108 107332 140110 107372
rect 140272 107332 140281 107372
rect 139895 107290 139942 107332
rect 140066 107290 140110 107332
rect 140234 107290 140281 107332
rect 78175 106616 78222 106658
rect 78346 106616 78390 106658
rect 78514 106616 78561 106658
rect 78175 106576 78184 106616
rect 78346 106576 78348 106616
rect 78388 106576 78390 106616
rect 78552 106576 78561 106616
rect 78175 106534 78222 106576
rect 78346 106534 78390 106576
rect 78514 106534 78561 106576
rect 93295 106616 93342 106658
rect 93466 106616 93510 106658
rect 93634 106616 93681 106658
rect 93295 106576 93304 106616
rect 93466 106576 93468 106616
rect 93508 106576 93510 106616
rect 93672 106576 93681 106616
rect 93295 106534 93342 106576
rect 93466 106534 93510 106576
rect 93634 106534 93681 106576
rect 108415 106616 108462 106658
rect 108586 106616 108630 106658
rect 108754 106616 108801 106658
rect 108415 106576 108424 106616
rect 108586 106576 108588 106616
rect 108628 106576 108630 106616
rect 108792 106576 108801 106616
rect 108415 106534 108462 106576
rect 108586 106534 108630 106576
rect 108754 106534 108801 106576
rect 123535 106616 123582 106658
rect 123706 106616 123750 106658
rect 123874 106616 123921 106658
rect 123535 106576 123544 106616
rect 123706 106576 123708 106616
rect 123748 106576 123750 106616
rect 123912 106576 123921 106616
rect 123535 106534 123582 106576
rect 123706 106534 123750 106576
rect 123874 106534 123921 106576
rect 138655 106616 138702 106658
rect 138826 106616 138870 106658
rect 138994 106616 139041 106658
rect 138655 106576 138664 106616
rect 138826 106576 138828 106616
rect 138868 106576 138870 106616
rect 139032 106576 139041 106616
rect 138655 106534 138702 106576
rect 138826 106534 138870 106576
rect 138994 106534 139041 106576
rect 79415 105860 79462 105902
rect 79586 105860 79630 105902
rect 79754 105860 79801 105902
rect 79415 105820 79424 105860
rect 79586 105820 79588 105860
rect 79628 105820 79630 105860
rect 79792 105820 79801 105860
rect 79415 105778 79462 105820
rect 79586 105778 79630 105820
rect 79754 105778 79801 105820
rect 94535 105860 94582 105902
rect 94706 105860 94750 105902
rect 94874 105860 94921 105902
rect 94535 105820 94544 105860
rect 94706 105820 94708 105860
rect 94748 105820 94750 105860
rect 94912 105820 94921 105860
rect 94535 105778 94582 105820
rect 94706 105778 94750 105820
rect 94874 105778 94921 105820
rect 109655 105860 109702 105902
rect 109826 105860 109870 105902
rect 109994 105860 110041 105902
rect 109655 105820 109664 105860
rect 109826 105820 109828 105860
rect 109868 105820 109870 105860
rect 110032 105820 110041 105860
rect 109655 105778 109702 105820
rect 109826 105778 109870 105820
rect 109994 105778 110041 105820
rect 124775 105860 124822 105902
rect 124946 105860 124990 105902
rect 125114 105860 125161 105902
rect 124775 105820 124784 105860
rect 124946 105820 124948 105860
rect 124988 105820 124990 105860
rect 125152 105820 125161 105860
rect 124775 105778 124822 105820
rect 124946 105778 124990 105820
rect 125114 105778 125161 105820
rect 139895 105860 139942 105902
rect 140066 105860 140110 105902
rect 140234 105860 140281 105902
rect 139895 105820 139904 105860
rect 140066 105820 140068 105860
rect 140108 105820 140110 105860
rect 140272 105820 140281 105860
rect 139895 105778 139942 105820
rect 140066 105778 140110 105820
rect 140234 105778 140281 105820
rect 78175 105104 78222 105146
rect 78346 105104 78390 105146
rect 78514 105104 78561 105146
rect 78175 105064 78184 105104
rect 78346 105064 78348 105104
rect 78388 105064 78390 105104
rect 78552 105064 78561 105104
rect 78175 105022 78222 105064
rect 78346 105022 78390 105064
rect 78514 105022 78561 105064
rect 93295 105104 93342 105146
rect 93466 105104 93510 105146
rect 93634 105104 93681 105146
rect 93295 105064 93304 105104
rect 93466 105064 93468 105104
rect 93508 105064 93510 105104
rect 93672 105064 93681 105104
rect 93295 105022 93342 105064
rect 93466 105022 93510 105064
rect 93634 105022 93681 105064
rect 108415 105104 108462 105146
rect 108586 105104 108630 105146
rect 108754 105104 108801 105146
rect 108415 105064 108424 105104
rect 108586 105064 108588 105104
rect 108628 105064 108630 105104
rect 108792 105064 108801 105104
rect 108415 105022 108462 105064
rect 108586 105022 108630 105064
rect 108754 105022 108801 105064
rect 123535 105104 123582 105146
rect 123706 105104 123750 105146
rect 123874 105104 123921 105146
rect 123535 105064 123544 105104
rect 123706 105064 123708 105104
rect 123748 105064 123750 105104
rect 123912 105064 123921 105104
rect 123535 105022 123582 105064
rect 123706 105022 123750 105064
rect 123874 105022 123921 105064
rect 138655 105104 138702 105146
rect 138826 105104 138870 105146
rect 138994 105104 139041 105146
rect 138655 105064 138664 105104
rect 138826 105064 138828 105104
rect 138868 105064 138870 105104
rect 139032 105064 139041 105104
rect 138655 105022 138702 105064
rect 138826 105022 138870 105064
rect 138994 105022 139041 105064
rect 79415 104348 79462 104390
rect 79586 104348 79630 104390
rect 79754 104348 79801 104390
rect 79415 104308 79424 104348
rect 79586 104308 79588 104348
rect 79628 104308 79630 104348
rect 79792 104308 79801 104348
rect 79415 104266 79462 104308
rect 79586 104266 79630 104308
rect 79754 104266 79801 104308
rect 94535 104348 94582 104390
rect 94706 104348 94750 104390
rect 94874 104348 94921 104390
rect 94535 104308 94544 104348
rect 94706 104308 94708 104348
rect 94748 104308 94750 104348
rect 94912 104308 94921 104348
rect 94535 104266 94582 104308
rect 94706 104266 94750 104308
rect 94874 104266 94921 104308
rect 109655 104348 109702 104390
rect 109826 104348 109870 104390
rect 109994 104348 110041 104390
rect 109655 104308 109664 104348
rect 109826 104308 109828 104348
rect 109868 104308 109870 104348
rect 110032 104308 110041 104348
rect 109655 104266 109702 104308
rect 109826 104266 109870 104308
rect 109994 104266 110041 104308
rect 124775 104348 124822 104390
rect 124946 104348 124990 104390
rect 125114 104348 125161 104390
rect 124775 104308 124784 104348
rect 124946 104308 124948 104348
rect 124988 104308 124990 104348
rect 125152 104308 125161 104348
rect 124775 104266 124822 104308
rect 124946 104266 124990 104308
rect 125114 104266 125161 104308
rect 139895 104348 139942 104390
rect 140066 104348 140110 104390
rect 140234 104348 140281 104390
rect 139895 104308 139904 104348
rect 140066 104308 140068 104348
rect 140108 104308 140110 104348
rect 140272 104308 140281 104348
rect 139895 104266 139942 104308
rect 140066 104266 140110 104308
rect 140234 104266 140281 104308
rect 78175 103592 78222 103634
rect 78346 103592 78390 103634
rect 78514 103592 78561 103634
rect 78175 103552 78184 103592
rect 78346 103552 78348 103592
rect 78388 103552 78390 103592
rect 78552 103552 78561 103592
rect 78175 103510 78222 103552
rect 78346 103510 78390 103552
rect 78514 103510 78561 103552
rect 93295 103592 93342 103634
rect 93466 103592 93510 103634
rect 93634 103592 93681 103634
rect 93295 103552 93304 103592
rect 93466 103552 93468 103592
rect 93508 103552 93510 103592
rect 93672 103552 93681 103592
rect 93295 103510 93342 103552
rect 93466 103510 93510 103552
rect 93634 103510 93681 103552
rect 108415 103592 108462 103634
rect 108586 103592 108630 103634
rect 108754 103592 108801 103634
rect 108415 103552 108424 103592
rect 108586 103552 108588 103592
rect 108628 103552 108630 103592
rect 108792 103552 108801 103592
rect 108415 103510 108462 103552
rect 108586 103510 108630 103552
rect 108754 103510 108801 103552
rect 123535 103592 123582 103634
rect 123706 103592 123750 103634
rect 123874 103592 123921 103634
rect 123535 103552 123544 103592
rect 123706 103552 123708 103592
rect 123748 103552 123750 103592
rect 123912 103552 123921 103592
rect 123535 103510 123582 103552
rect 123706 103510 123750 103552
rect 123874 103510 123921 103552
rect 138655 103592 138702 103634
rect 138826 103592 138870 103634
rect 138994 103592 139041 103634
rect 138655 103552 138664 103592
rect 138826 103552 138828 103592
rect 138868 103552 138870 103592
rect 139032 103552 139041 103592
rect 138655 103510 138702 103552
rect 138826 103510 138870 103552
rect 138994 103510 139041 103552
rect 79415 102836 79462 102878
rect 79586 102836 79630 102878
rect 79754 102836 79801 102878
rect 79415 102796 79424 102836
rect 79586 102796 79588 102836
rect 79628 102796 79630 102836
rect 79792 102796 79801 102836
rect 79415 102754 79462 102796
rect 79586 102754 79630 102796
rect 79754 102754 79801 102796
rect 94535 102836 94582 102878
rect 94706 102836 94750 102878
rect 94874 102836 94921 102878
rect 94535 102796 94544 102836
rect 94706 102796 94708 102836
rect 94748 102796 94750 102836
rect 94912 102796 94921 102836
rect 94535 102754 94582 102796
rect 94706 102754 94750 102796
rect 94874 102754 94921 102796
rect 109655 102836 109702 102878
rect 109826 102836 109870 102878
rect 109994 102836 110041 102878
rect 109655 102796 109664 102836
rect 109826 102796 109828 102836
rect 109868 102796 109870 102836
rect 110032 102796 110041 102836
rect 109655 102754 109702 102796
rect 109826 102754 109870 102796
rect 109994 102754 110041 102796
rect 124775 102836 124822 102878
rect 124946 102836 124990 102878
rect 125114 102836 125161 102878
rect 124775 102796 124784 102836
rect 124946 102796 124948 102836
rect 124988 102796 124990 102836
rect 125152 102796 125161 102836
rect 124775 102754 124822 102796
rect 124946 102754 124990 102796
rect 125114 102754 125161 102796
rect 139895 102836 139942 102878
rect 140066 102836 140110 102878
rect 140234 102836 140281 102878
rect 139895 102796 139904 102836
rect 140066 102796 140068 102836
rect 140108 102796 140110 102836
rect 140272 102796 140281 102836
rect 139895 102754 139942 102796
rect 140066 102754 140110 102796
rect 140234 102754 140281 102796
rect 78175 102080 78222 102122
rect 78346 102080 78390 102122
rect 78514 102080 78561 102122
rect 78175 102040 78184 102080
rect 78346 102040 78348 102080
rect 78388 102040 78390 102080
rect 78552 102040 78561 102080
rect 78175 101998 78222 102040
rect 78346 101998 78390 102040
rect 78514 101998 78561 102040
rect 93295 102080 93342 102122
rect 93466 102080 93510 102122
rect 93634 102080 93681 102122
rect 93295 102040 93304 102080
rect 93466 102040 93468 102080
rect 93508 102040 93510 102080
rect 93672 102040 93681 102080
rect 93295 101998 93342 102040
rect 93466 101998 93510 102040
rect 93634 101998 93681 102040
rect 108415 102080 108462 102122
rect 108586 102080 108630 102122
rect 108754 102080 108801 102122
rect 108415 102040 108424 102080
rect 108586 102040 108588 102080
rect 108628 102040 108630 102080
rect 108792 102040 108801 102080
rect 108415 101998 108462 102040
rect 108586 101998 108630 102040
rect 108754 101998 108801 102040
rect 123535 102080 123582 102122
rect 123706 102080 123750 102122
rect 123874 102080 123921 102122
rect 123535 102040 123544 102080
rect 123706 102040 123708 102080
rect 123748 102040 123750 102080
rect 123912 102040 123921 102080
rect 123535 101998 123582 102040
rect 123706 101998 123750 102040
rect 123874 101998 123921 102040
rect 138655 102080 138702 102122
rect 138826 102080 138870 102122
rect 138994 102080 139041 102122
rect 138655 102040 138664 102080
rect 138826 102040 138828 102080
rect 138868 102040 138870 102080
rect 139032 102040 139041 102080
rect 138655 101998 138702 102040
rect 138826 101998 138870 102040
rect 138994 101998 139041 102040
rect 79415 101324 79462 101366
rect 79586 101324 79630 101366
rect 79754 101324 79801 101366
rect 79415 101284 79424 101324
rect 79586 101284 79588 101324
rect 79628 101284 79630 101324
rect 79792 101284 79801 101324
rect 79415 101242 79462 101284
rect 79586 101242 79630 101284
rect 79754 101242 79801 101284
rect 94535 101324 94582 101366
rect 94706 101324 94750 101366
rect 94874 101324 94921 101366
rect 94535 101284 94544 101324
rect 94706 101284 94708 101324
rect 94748 101284 94750 101324
rect 94912 101284 94921 101324
rect 94535 101242 94582 101284
rect 94706 101242 94750 101284
rect 94874 101242 94921 101284
rect 109655 101324 109702 101366
rect 109826 101324 109870 101366
rect 109994 101324 110041 101366
rect 109655 101284 109664 101324
rect 109826 101284 109828 101324
rect 109868 101284 109870 101324
rect 110032 101284 110041 101324
rect 109655 101242 109702 101284
rect 109826 101242 109870 101284
rect 109994 101242 110041 101284
rect 124775 101324 124822 101366
rect 124946 101324 124990 101366
rect 125114 101324 125161 101366
rect 124775 101284 124784 101324
rect 124946 101284 124948 101324
rect 124988 101284 124990 101324
rect 125152 101284 125161 101324
rect 124775 101242 124822 101284
rect 124946 101242 124990 101284
rect 125114 101242 125161 101284
rect 139895 101324 139942 101366
rect 140066 101324 140110 101366
rect 140234 101324 140281 101366
rect 139895 101284 139904 101324
rect 140066 101284 140068 101324
rect 140108 101284 140110 101324
rect 140272 101284 140281 101324
rect 139895 101242 139942 101284
rect 140066 101242 140110 101284
rect 140234 101242 140281 101284
rect 78175 100568 78222 100610
rect 78346 100568 78390 100610
rect 78514 100568 78561 100610
rect 78175 100528 78184 100568
rect 78346 100528 78348 100568
rect 78388 100528 78390 100568
rect 78552 100528 78561 100568
rect 78175 100486 78222 100528
rect 78346 100486 78390 100528
rect 78514 100486 78561 100528
rect 93295 100568 93342 100610
rect 93466 100568 93510 100610
rect 93634 100568 93681 100610
rect 93295 100528 93304 100568
rect 93466 100528 93468 100568
rect 93508 100528 93510 100568
rect 93672 100528 93681 100568
rect 93295 100486 93342 100528
rect 93466 100486 93510 100528
rect 93634 100486 93681 100528
rect 108415 100568 108462 100610
rect 108586 100568 108630 100610
rect 108754 100568 108801 100610
rect 108415 100528 108424 100568
rect 108586 100528 108588 100568
rect 108628 100528 108630 100568
rect 108792 100528 108801 100568
rect 108415 100486 108462 100528
rect 108586 100486 108630 100528
rect 108754 100486 108801 100528
rect 123535 100568 123582 100610
rect 123706 100568 123750 100610
rect 123874 100568 123921 100610
rect 123535 100528 123544 100568
rect 123706 100528 123708 100568
rect 123748 100528 123750 100568
rect 123912 100528 123921 100568
rect 123535 100486 123582 100528
rect 123706 100486 123750 100528
rect 123874 100486 123921 100528
rect 138655 100568 138702 100610
rect 138826 100568 138870 100610
rect 138994 100568 139041 100610
rect 138655 100528 138664 100568
rect 138826 100528 138828 100568
rect 138868 100528 138870 100568
rect 139032 100528 139041 100568
rect 138655 100486 138702 100528
rect 138826 100486 138870 100528
rect 138994 100486 139041 100528
rect 79415 99812 79462 99854
rect 79586 99812 79630 99854
rect 79754 99812 79801 99854
rect 79415 99772 79424 99812
rect 79586 99772 79588 99812
rect 79628 99772 79630 99812
rect 79792 99772 79801 99812
rect 79415 99730 79462 99772
rect 79586 99730 79630 99772
rect 79754 99730 79801 99772
rect 94535 99812 94582 99854
rect 94706 99812 94750 99854
rect 94874 99812 94921 99854
rect 94535 99772 94544 99812
rect 94706 99772 94708 99812
rect 94748 99772 94750 99812
rect 94912 99772 94921 99812
rect 94535 99730 94582 99772
rect 94706 99730 94750 99772
rect 94874 99730 94921 99772
rect 109655 99812 109702 99854
rect 109826 99812 109870 99854
rect 109994 99812 110041 99854
rect 109655 99772 109664 99812
rect 109826 99772 109828 99812
rect 109868 99772 109870 99812
rect 110032 99772 110041 99812
rect 109655 99730 109702 99772
rect 109826 99730 109870 99772
rect 109994 99730 110041 99772
rect 124775 99812 124822 99854
rect 124946 99812 124990 99854
rect 125114 99812 125161 99854
rect 124775 99772 124784 99812
rect 124946 99772 124948 99812
rect 124988 99772 124990 99812
rect 125152 99772 125161 99812
rect 124775 99730 124822 99772
rect 124946 99730 124990 99772
rect 125114 99730 125161 99772
rect 139895 99812 139942 99854
rect 140066 99812 140110 99854
rect 140234 99812 140281 99854
rect 139895 99772 139904 99812
rect 140066 99772 140068 99812
rect 140108 99772 140110 99812
rect 140272 99772 140281 99812
rect 139895 99730 139942 99772
rect 140066 99730 140110 99772
rect 140234 99730 140281 99772
rect 78175 99056 78222 99098
rect 78346 99056 78390 99098
rect 78514 99056 78561 99098
rect 78175 99016 78184 99056
rect 78346 99016 78348 99056
rect 78388 99016 78390 99056
rect 78552 99016 78561 99056
rect 78175 98974 78222 99016
rect 78346 98974 78390 99016
rect 78514 98974 78561 99016
rect 93295 99056 93342 99098
rect 93466 99056 93510 99098
rect 93634 99056 93681 99098
rect 93295 99016 93304 99056
rect 93466 99016 93468 99056
rect 93508 99016 93510 99056
rect 93672 99016 93681 99056
rect 93295 98974 93342 99016
rect 93466 98974 93510 99016
rect 93634 98974 93681 99016
rect 108415 99056 108462 99098
rect 108586 99056 108630 99098
rect 108754 99056 108801 99098
rect 108415 99016 108424 99056
rect 108586 99016 108588 99056
rect 108628 99016 108630 99056
rect 108792 99016 108801 99056
rect 108415 98974 108462 99016
rect 108586 98974 108630 99016
rect 108754 98974 108801 99016
rect 123535 99056 123582 99098
rect 123706 99056 123750 99098
rect 123874 99056 123921 99098
rect 123535 99016 123544 99056
rect 123706 99016 123708 99056
rect 123748 99016 123750 99056
rect 123912 99016 123921 99056
rect 123535 98974 123582 99016
rect 123706 98974 123750 99016
rect 123874 98974 123921 99016
rect 138655 99056 138702 99098
rect 138826 99056 138870 99098
rect 138994 99056 139041 99098
rect 138655 99016 138664 99056
rect 138826 99016 138828 99056
rect 138868 99016 138870 99056
rect 139032 99016 139041 99056
rect 138655 98974 138702 99016
rect 138826 98974 138870 99016
rect 138994 98974 139041 99016
rect 79415 98300 79462 98342
rect 79586 98300 79630 98342
rect 79754 98300 79801 98342
rect 79415 98260 79424 98300
rect 79586 98260 79588 98300
rect 79628 98260 79630 98300
rect 79792 98260 79801 98300
rect 79415 98218 79462 98260
rect 79586 98218 79630 98260
rect 79754 98218 79801 98260
rect 94535 98300 94582 98342
rect 94706 98300 94750 98342
rect 94874 98300 94921 98342
rect 94535 98260 94544 98300
rect 94706 98260 94708 98300
rect 94748 98260 94750 98300
rect 94912 98260 94921 98300
rect 94535 98218 94582 98260
rect 94706 98218 94750 98260
rect 94874 98218 94921 98260
rect 109655 98300 109702 98342
rect 109826 98300 109870 98342
rect 109994 98300 110041 98342
rect 109655 98260 109664 98300
rect 109826 98260 109828 98300
rect 109868 98260 109870 98300
rect 110032 98260 110041 98300
rect 109655 98218 109702 98260
rect 109826 98218 109870 98260
rect 109994 98218 110041 98260
rect 124775 98300 124822 98342
rect 124946 98300 124990 98342
rect 125114 98300 125161 98342
rect 124775 98260 124784 98300
rect 124946 98260 124948 98300
rect 124988 98260 124990 98300
rect 125152 98260 125161 98300
rect 124775 98218 124822 98260
rect 124946 98218 124990 98260
rect 125114 98218 125161 98260
rect 139895 98300 139942 98342
rect 140066 98300 140110 98342
rect 140234 98300 140281 98342
rect 139895 98260 139904 98300
rect 140066 98260 140068 98300
rect 140108 98260 140110 98300
rect 140272 98260 140281 98300
rect 139895 98218 139942 98260
rect 140066 98218 140110 98260
rect 140234 98218 140281 98260
rect 78175 97544 78222 97586
rect 78346 97544 78390 97586
rect 78514 97544 78561 97586
rect 78175 97504 78184 97544
rect 78346 97504 78348 97544
rect 78388 97504 78390 97544
rect 78552 97504 78561 97544
rect 78175 97462 78222 97504
rect 78346 97462 78390 97504
rect 78514 97462 78561 97504
rect 93295 97544 93342 97586
rect 93466 97544 93510 97586
rect 93634 97544 93681 97586
rect 93295 97504 93304 97544
rect 93466 97504 93468 97544
rect 93508 97504 93510 97544
rect 93672 97504 93681 97544
rect 93295 97462 93342 97504
rect 93466 97462 93510 97504
rect 93634 97462 93681 97504
rect 108415 97544 108462 97586
rect 108586 97544 108630 97586
rect 108754 97544 108801 97586
rect 108415 97504 108424 97544
rect 108586 97504 108588 97544
rect 108628 97504 108630 97544
rect 108792 97504 108801 97544
rect 108415 97462 108462 97504
rect 108586 97462 108630 97504
rect 108754 97462 108801 97504
rect 123535 97544 123582 97586
rect 123706 97544 123750 97586
rect 123874 97544 123921 97586
rect 123535 97504 123544 97544
rect 123706 97504 123708 97544
rect 123748 97504 123750 97544
rect 123912 97504 123921 97544
rect 123535 97462 123582 97504
rect 123706 97462 123750 97504
rect 123874 97462 123921 97504
rect 138655 97544 138702 97586
rect 138826 97544 138870 97586
rect 138994 97544 139041 97586
rect 138655 97504 138664 97544
rect 138826 97504 138828 97544
rect 138868 97504 138870 97544
rect 139032 97504 139041 97544
rect 138655 97462 138702 97504
rect 138826 97462 138870 97504
rect 138994 97462 139041 97504
rect 79415 96788 79462 96830
rect 79586 96788 79630 96830
rect 79754 96788 79801 96830
rect 79415 96748 79424 96788
rect 79586 96748 79588 96788
rect 79628 96748 79630 96788
rect 79792 96748 79801 96788
rect 79415 96706 79462 96748
rect 79586 96706 79630 96748
rect 79754 96706 79801 96748
rect 94535 96788 94582 96830
rect 94706 96788 94750 96830
rect 94874 96788 94921 96830
rect 94535 96748 94544 96788
rect 94706 96748 94708 96788
rect 94748 96748 94750 96788
rect 94912 96748 94921 96788
rect 94535 96706 94582 96748
rect 94706 96706 94750 96748
rect 94874 96706 94921 96748
rect 109655 96788 109702 96830
rect 109826 96788 109870 96830
rect 109994 96788 110041 96830
rect 109655 96748 109664 96788
rect 109826 96748 109828 96788
rect 109868 96748 109870 96788
rect 110032 96748 110041 96788
rect 109655 96706 109702 96748
rect 109826 96706 109870 96748
rect 109994 96706 110041 96748
rect 124775 96788 124822 96830
rect 124946 96788 124990 96830
rect 125114 96788 125161 96830
rect 124775 96748 124784 96788
rect 124946 96748 124948 96788
rect 124988 96748 124990 96788
rect 125152 96748 125161 96788
rect 124775 96706 124822 96748
rect 124946 96706 124990 96748
rect 125114 96706 125161 96748
rect 139895 96788 139942 96830
rect 140066 96788 140110 96830
rect 140234 96788 140281 96830
rect 139895 96748 139904 96788
rect 140066 96748 140068 96788
rect 140108 96748 140110 96788
rect 140272 96748 140281 96788
rect 139895 96706 139942 96748
rect 140066 96706 140110 96748
rect 140234 96706 140281 96748
rect 78175 96032 78222 96074
rect 78346 96032 78390 96074
rect 78514 96032 78561 96074
rect 78175 95992 78184 96032
rect 78346 95992 78348 96032
rect 78388 95992 78390 96032
rect 78552 95992 78561 96032
rect 78175 95950 78222 95992
rect 78346 95950 78390 95992
rect 78514 95950 78561 95992
rect 93295 96032 93342 96074
rect 93466 96032 93510 96074
rect 93634 96032 93681 96074
rect 93295 95992 93304 96032
rect 93466 95992 93468 96032
rect 93508 95992 93510 96032
rect 93672 95992 93681 96032
rect 93295 95950 93342 95992
rect 93466 95950 93510 95992
rect 93634 95950 93681 95992
rect 108415 96032 108462 96074
rect 108586 96032 108630 96074
rect 108754 96032 108801 96074
rect 108415 95992 108424 96032
rect 108586 95992 108588 96032
rect 108628 95992 108630 96032
rect 108792 95992 108801 96032
rect 108415 95950 108462 95992
rect 108586 95950 108630 95992
rect 108754 95950 108801 95992
rect 123535 96032 123582 96074
rect 123706 96032 123750 96074
rect 123874 96032 123921 96074
rect 123535 95992 123544 96032
rect 123706 95992 123708 96032
rect 123748 95992 123750 96032
rect 123912 95992 123921 96032
rect 123535 95950 123582 95992
rect 123706 95950 123750 95992
rect 123874 95950 123921 95992
rect 138655 96032 138702 96074
rect 138826 96032 138870 96074
rect 138994 96032 139041 96074
rect 138655 95992 138664 96032
rect 138826 95992 138828 96032
rect 138868 95992 138870 96032
rect 139032 95992 139041 96032
rect 138655 95950 138702 95992
rect 138826 95950 138870 95992
rect 138994 95950 139041 95992
rect 79415 95276 79462 95318
rect 79586 95276 79630 95318
rect 79754 95276 79801 95318
rect 79415 95236 79424 95276
rect 79586 95236 79588 95276
rect 79628 95236 79630 95276
rect 79792 95236 79801 95276
rect 79415 95194 79462 95236
rect 79586 95194 79630 95236
rect 79754 95194 79801 95236
rect 94535 95276 94582 95318
rect 94706 95276 94750 95318
rect 94874 95276 94921 95318
rect 94535 95236 94544 95276
rect 94706 95236 94708 95276
rect 94748 95236 94750 95276
rect 94912 95236 94921 95276
rect 94535 95194 94582 95236
rect 94706 95194 94750 95236
rect 94874 95194 94921 95236
rect 109655 95276 109702 95318
rect 109826 95276 109870 95318
rect 109994 95276 110041 95318
rect 109655 95236 109664 95276
rect 109826 95236 109828 95276
rect 109868 95236 109870 95276
rect 110032 95236 110041 95276
rect 109655 95194 109702 95236
rect 109826 95194 109870 95236
rect 109994 95194 110041 95236
rect 124775 95276 124822 95318
rect 124946 95276 124990 95318
rect 125114 95276 125161 95318
rect 124775 95236 124784 95276
rect 124946 95236 124948 95276
rect 124988 95236 124990 95276
rect 125152 95236 125161 95276
rect 124775 95194 124822 95236
rect 124946 95194 124990 95236
rect 125114 95194 125161 95236
rect 139895 95276 139942 95318
rect 140066 95276 140110 95318
rect 140234 95276 140281 95318
rect 139895 95236 139904 95276
rect 140066 95236 140068 95276
rect 140108 95236 140110 95276
rect 140272 95236 140281 95276
rect 139895 95194 139942 95236
rect 140066 95194 140110 95236
rect 140234 95194 140281 95236
rect 78175 94520 78222 94562
rect 78346 94520 78390 94562
rect 78514 94520 78561 94562
rect 78175 94480 78184 94520
rect 78346 94480 78348 94520
rect 78388 94480 78390 94520
rect 78552 94480 78561 94520
rect 78175 94438 78222 94480
rect 78346 94438 78390 94480
rect 78514 94438 78561 94480
rect 93295 94520 93342 94562
rect 93466 94520 93510 94562
rect 93634 94520 93681 94562
rect 93295 94480 93304 94520
rect 93466 94480 93468 94520
rect 93508 94480 93510 94520
rect 93672 94480 93681 94520
rect 93295 94438 93342 94480
rect 93466 94438 93510 94480
rect 93634 94438 93681 94480
rect 108415 94520 108462 94562
rect 108586 94520 108630 94562
rect 108754 94520 108801 94562
rect 108415 94480 108424 94520
rect 108586 94480 108588 94520
rect 108628 94480 108630 94520
rect 108792 94480 108801 94520
rect 108415 94438 108462 94480
rect 108586 94438 108630 94480
rect 108754 94438 108801 94480
rect 123535 94520 123582 94562
rect 123706 94520 123750 94562
rect 123874 94520 123921 94562
rect 123535 94480 123544 94520
rect 123706 94480 123708 94520
rect 123748 94480 123750 94520
rect 123912 94480 123921 94520
rect 123535 94438 123582 94480
rect 123706 94438 123750 94480
rect 123874 94438 123921 94480
rect 138655 94520 138702 94562
rect 138826 94520 138870 94562
rect 138994 94520 139041 94562
rect 138655 94480 138664 94520
rect 138826 94480 138828 94520
rect 138868 94480 138870 94520
rect 139032 94480 139041 94520
rect 138655 94438 138702 94480
rect 138826 94438 138870 94480
rect 138994 94438 139041 94480
rect 79415 93764 79462 93806
rect 79586 93764 79630 93806
rect 79754 93764 79801 93806
rect 79415 93724 79424 93764
rect 79586 93724 79588 93764
rect 79628 93724 79630 93764
rect 79792 93724 79801 93764
rect 79415 93682 79462 93724
rect 79586 93682 79630 93724
rect 79754 93682 79801 93724
rect 94535 93764 94582 93806
rect 94706 93764 94750 93806
rect 94874 93764 94921 93806
rect 94535 93724 94544 93764
rect 94706 93724 94708 93764
rect 94748 93724 94750 93764
rect 94912 93724 94921 93764
rect 94535 93682 94582 93724
rect 94706 93682 94750 93724
rect 94874 93682 94921 93724
rect 109655 93764 109702 93806
rect 109826 93764 109870 93806
rect 109994 93764 110041 93806
rect 109655 93724 109664 93764
rect 109826 93724 109828 93764
rect 109868 93724 109870 93764
rect 110032 93724 110041 93764
rect 109655 93682 109702 93724
rect 109826 93682 109870 93724
rect 109994 93682 110041 93724
rect 124775 93764 124822 93806
rect 124946 93764 124990 93806
rect 125114 93764 125161 93806
rect 124775 93724 124784 93764
rect 124946 93724 124948 93764
rect 124988 93724 124990 93764
rect 125152 93724 125161 93764
rect 124775 93682 124822 93724
rect 124946 93682 124990 93724
rect 125114 93682 125161 93724
rect 139895 93764 139942 93806
rect 140066 93764 140110 93806
rect 140234 93764 140281 93806
rect 139895 93724 139904 93764
rect 140066 93724 140068 93764
rect 140108 93724 140110 93764
rect 140272 93724 140281 93764
rect 139895 93682 139942 93724
rect 140066 93682 140110 93724
rect 140234 93682 140281 93724
rect 78175 93008 78222 93050
rect 78346 93008 78390 93050
rect 78514 93008 78561 93050
rect 78175 92968 78184 93008
rect 78346 92968 78348 93008
rect 78388 92968 78390 93008
rect 78552 92968 78561 93008
rect 78175 92926 78222 92968
rect 78346 92926 78390 92968
rect 78514 92926 78561 92968
rect 93295 93008 93342 93050
rect 93466 93008 93510 93050
rect 93634 93008 93681 93050
rect 93295 92968 93304 93008
rect 93466 92968 93468 93008
rect 93508 92968 93510 93008
rect 93672 92968 93681 93008
rect 93295 92926 93342 92968
rect 93466 92926 93510 92968
rect 93634 92926 93681 92968
rect 108415 93008 108462 93050
rect 108586 93008 108630 93050
rect 108754 93008 108801 93050
rect 108415 92968 108424 93008
rect 108586 92968 108588 93008
rect 108628 92968 108630 93008
rect 108792 92968 108801 93008
rect 108415 92926 108462 92968
rect 108586 92926 108630 92968
rect 108754 92926 108801 92968
rect 123535 93008 123582 93050
rect 123706 93008 123750 93050
rect 123874 93008 123921 93050
rect 123535 92968 123544 93008
rect 123706 92968 123708 93008
rect 123748 92968 123750 93008
rect 123912 92968 123921 93008
rect 123535 92926 123582 92968
rect 123706 92926 123750 92968
rect 123874 92926 123921 92968
rect 138655 93008 138702 93050
rect 138826 93008 138870 93050
rect 138994 93008 139041 93050
rect 138655 92968 138664 93008
rect 138826 92968 138828 93008
rect 138868 92968 138870 93008
rect 139032 92968 139041 93008
rect 138655 92926 138702 92968
rect 138826 92926 138870 92968
rect 138994 92926 139041 92968
rect 79415 92252 79462 92294
rect 79586 92252 79630 92294
rect 79754 92252 79801 92294
rect 79415 92212 79424 92252
rect 79586 92212 79588 92252
rect 79628 92212 79630 92252
rect 79792 92212 79801 92252
rect 79415 92170 79462 92212
rect 79586 92170 79630 92212
rect 79754 92170 79801 92212
rect 94535 92252 94582 92294
rect 94706 92252 94750 92294
rect 94874 92252 94921 92294
rect 94535 92212 94544 92252
rect 94706 92212 94708 92252
rect 94748 92212 94750 92252
rect 94912 92212 94921 92252
rect 94535 92170 94582 92212
rect 94706 92170 94750 92212
rect 94874 92170 94921 92212
rect 109655 92252 109702 92294
rect 109826 92252 109870 92294
rect 109994 92252 110041 92294
rect 109655 92212 109664 92252
rect 109826 92212 109828 92252
rect 109868 92212 109870 92252
rect 110032 92212 110041 92252
rect 109655 92170 109702 92212
rect 109826 92170 109870 92212
rect 109994 92170 110041 92212
rect 124775 92252 124822 92294
rect 124946 92252 124990 92294
rect 125114 92252 125161 92294
rect 124775 92212 124784 92252
rect 124946 92212 124948 92252
rect 124988 92212 124990 92252
rect 125152 92212 125161 92252
rect 124775 92170 124822 92212
rect 124946 92170 124990 92212
rect 125114 92170 125161 92212
rect 139895 92252 139942 92294
rect 140066 92252 140110 92294
rect 140234 92252 140281 92294
rect 139895 92212 139904 92252
rect 140066 92212 140068 92252
rect 140108 92212 140110 92252
rect 140272 92212 140281 92252
rect 139895 92170 139942 92212
rect 140066 92170 140110 92212
rect 140234 92170 140281 92212
rect 78175 91496 78222 91538
rect 78346 91496 78390 91538
rect 78514 91496 78561 91538
rect 78175 91456 78184 91496
rect 78346 91456 78348 91496
rect 78388 91456 78390 91496
rect 78552 91456 78561 91496
rect 78175 91414 78222 91456
rect 78346 91414 78390 91456
rect 78514 91414 78561 91456
rect 93295 91496 93342 91538
rect 93466 91496 93510 91538
rect 93634 91496 93681 91538
rect 93295 91456 93304 91496
rect 93466 91456 93468 91496
rect 93508 91456 93510 91496
rect 93672 91456 93681 91496
rect 93295 91414 93342 91456
rect 93466 91414 93510 91456
rect 93634 91414 93681 91456
rect 108415 91496 108462 91538
rect 108586 91496 108630 91538
rect 108754 91496 108801 91538
rect 108415 91456 108424 91496
rect 108586 91456 108588 91496
rect 108628 91456 108630 91496
rect 108792 91456 108801 91496
rect 108415 91414 108462 91456
rect 108586 91414 108630 91456
rect 108754 91414 108801 91456
rect 123535 91496 123582 91538
rect 123706 91496 123750 91538
rect 123874 91496 123921 91538
rect 123535 91456 123544 91496
rect 123706 91456 123708 91496
rect 123748 91456 123750 91496
rect 123912 91456 123921 91496
rect 123535 91414 123582 91456
rect 123706 91414 123750 91456
rect 123874 91414 123921 91456
rect 138655 91496 138702 91538
rect 138826 91496 138870 91538
rect 138994 91496 139041 91538
rect 138655 91456 138664 91496
rect 138826 91456 138828 91496
rect 138868 91456 138870 91496
rect 139032 91456 139041 91496
rect 138655 91414 138702 91456
rect 138826 91414 138870 91456
rect 138994 91414 139041 91456
rect 79415 90740 79462 90782
rect 79586 90740 79630 90782
rect 79754 90740 79801 90782
rect 79415 90700 79424 90740
rect 79586 90700 79588 90740
rect 79628 90700 79630 90740
rect 79792 90700 79801 90740
rect 79415 90658 79462 90700
rect 79586 90658 79630 90700
rect 79754 90658 79801 90700
rect 94535 90740 94582 90782
rect 94706 90740 94750 90782
rect 94874 90740 94921 90782
rect 94535 90700 94544 90740
rect 94706 90700 94708 90740
rect 94748 90700 94750 90740
rect 94912 90700 94921 90740
rect 94535 90658 94582 90700
rect 94706 90658 94750 90700
rect 94874 90658 94921 90700
rect 109655 90740 109702 90782
rect 109826 90740 109870 90782
rect 109994 90740 110041 90782
rect 109655 90700 109664 90740
rect 109826 90700 109828 90740
rect 109868 90700 109870 90740
rect 110032 90700 110041 90740
rect 109655 90658 109702 90700
rect 109826 90658 109870 90700
rect 109994 90658 110041 90700
rect 124775 90740 124822 90782
rect 124946 90740 124990 90782
rect 125114 90740 125161 90782
rect 124775 90700 124784 90740
rect 124946 90700 124948 90740
rect 124988 90700 124990 90740
rect 125152 90700 125161 90740
rect 124775 90658 124822 90700
rect 124946 90658 124990 90700
rect 125114 90658 125161 90700
rect 139895 90740 139942 90782
rect 140066 90740 140110 90782
rect 140234 90740 140281 90782
rect 139895 90700 139904 90740
rect 140066 90700 140068 90740
rect 140108 90700 140110 90740
rect 140272 90700 140281 90740
rect 139895 90658 139942 90700
rect 140066 90658 140110 90700
rect 140234 90658 140281 90700
rect 78175 89984 78222 90026
rect 78346 89984 78390 90026
rect 78514 89984 78561 90026
rect 78175 89944 78184 89984
rect 78346 89944 78348 89984
rect 78388 89944 78390 89984
rect 78552 89944 78561 89984
rect 78175 89902 78222 89944
rect 78346 89902 78390 89944
rect 78514 89902 78561 89944
rect 93295 89984 93342 90026
rect 93466 89984 93510 90026
rect 93634 89984 93681 90026
rect 93295 89944 93304 89984
rect 93466 89944 93468 89984
rect 93508 89944 93510 89984
rect 93672 89944 93681 89984
rect 93295 89902 93342 89944
rect 93466 89902 93510 89944
rect 93634 89902 93681 89944
rect 108415 89984 108462 90026
rect 108586 89984 108630 90026
rect 108754 89984 108801 90026
rect 108415 89944 108424 89984
rect 108586 89944 108588 89984
rect 108628 89944 108630 89984
rect 108792 89944 108801 89984
rect 108415 89902 108462 89944
rect 108586 89902 108630 89944
rect 108754 89902 108801 89944
rect 123535 89984 123582 90026
rect 123706 89984 123750 90026
rect 123874 89984 123921 90026
rect 123535 89944 123544 89984
rect 123706 89944 123708 89984
rect 123748 89944 123750 89984
rect 123912 89944 123921 89984
rect 123535 89902 123582 89944
rect 123706 89902 123750 89944
rect 123874 89902 123921 89944
rect 138655 89984 138702 90026
rect 138826 89984 138870 90026
rect 138994 89984 139041 90026
rect 138655 89944 138664 89984
rect 138826 89944 138828 89984
rect 138868 89944 138870 89984
rect 139032 89944 139041 89984
rect 138655 89902 138702 89944
rect 138826 89902 138870 89944
rect 138994 89902 139041 89944
rect 79415 89228 79462 89270
rect 79586 89228 79630 89270
rect 79754 89228 79801 89270
rect 79415 89188 79424 89228
rect 79586 89188 79588 89228
rect 79628 89188 79630 89228
rect 79792 89188 79801 89228
rect 79415 89146 79462 89188
rect 79586 89146 79630 89188
rect 79754 89146 79801 89188
rect 94535 89228 94582 89270
rect 94706 89228 94750 89270
rect 94874 89228 94921 89270
rect 94535 89188 94544 89228
rect 94706 89188 94708 89228
rect 94748 89188 94750 89228
rect 94912 89188 94921 89228
rect 94535 89146 94582 89188
rect 94706 89146 94750 89188
rect 94874 89146 94921 89188
rect 109655 89228 109702 89270
rect 109826 89228 109870 89270
rect 109994 89228 110041 89270
rect 109655 89188 109664 89228
rect 109826 89188 109828 89228
rect 109868 89188 109870 89228
rect 110032 89188 110041 89228
rect 109655 89146 109702 89188
rect 109826 89146 109870 89188
rect 109994 89146 110041 89188
rect 124775 89228 124822 89270
rect 124946 89228 124990 89270
rect 125114 89228 125161 89270
rect 124775 89188 124784 89228
rect 124946 89188 124948 89228
rect 124988 89188 124990 89228
rect 125152 89188 125161 89228
rect 124775 89146 124822 89188
rect 124946 89146 124990 89188
rect 125114 89146 125161 89188
rect 139895 89228 139942 89270
rect 140066 89228 140110 89270
rect 140234 89228 140281 89270
rect 139895 89188 139904 89228
rect 140066 89188 140068 89228
rect 140108 89188 140110 89228
rect 140272 89188 140281 89228
rect 139895 89146 139942 89188
rect 140066 89146 140110 89188
rect 140234 89146 140281 89188
rect 90691 89104 90700 89144
rect 90740 89104 92140 89144
rect 92180 89104 92189 89144
rect 78175 88472 78222 88514
rect 78346 88472 78390 88514
rect 78514 88472 78561 88514
rect 78175 88432 78184 88472
rect 78346 88432 78348 88472
rect 78388 88432 78390 88472
rect 78552 88432 78561 88472
rect 78175 88390 78222 88432
rect 78346 88390 78390 88432
rect 78514 88390 78561 88432
rect 93295 88472 93342 88514
rect 93466 88472 93510 88514
rect 93634 88472 93681 88514
rect 93295 88432 93304 88472
rect 93466 88432 93468 88472
rect 93508 88432 93510 88472
rect 93672 88432 93681 88472
rect 93295 88390 93342 88432
rect 93466 88390 93510 88432
rect 93634 88390 93681 88432
rect 108415 88472 108462 88514
rect 108586 88472 108630 88514
rect 108754 88472 108801 88514
rect 108415 88432 108424 88472
rect 108586 88432 108588 88472
rect 108628 88432 108630 88472
rect 108792 88432 108801 88472
rect 108415 88390 108462 88432
rect 108586 88390 108630 88432
rect 108754 88390 108801 88432
rect 123535 88472 123582 88514
rect 123706 88472 123750 88514
rect 123874 88472 123921 88514
rect 123535 88432 123544 88472
rect 123706 88432 123708 88472
rect 123748 88432 123750 88472
rect 123912 88432 123921 88472
rect 123535 88390 123582 88432
rect 123706 88390 123750 88432
rect 123874 88390 123921 88432
rect 138655 88472 138702 88514
rect 138826 88472 138870 88514
rect 138994 88472 139041 88514
rect 138655 88432 138664 88472
rect 138826 88432 138828 88472
rect 138868 88432 138870 88472
rect 139032 88432 139041 88472
rect 138655 88390 138702 88432
rect 138826 88390 138870 88432
rect 138994 88390 139041 88432
rect 79415 87716 79462 87758
rect 79586 87716 79630 87758
rect 79754 87716 79801 87758
rect 79415 87676 79424 87716
rect 79586 87676 79588 87716
rect 79628 87676 79630 87716
rect 79792 87676 79801 87716
rect 79415 87634 79462 87676
rect 79586 87634 79630 87676
rect 79754 87634 79801 87676
rect 94535 87716 94582 87758
rect 94706 87716 94750 87758
rect 94874 87716 94921 87758
rect 94535 87676 94544 87716
rect 94706 87676 94708 87716
rect 94748 87676 94750 87716
rect 94912 87676 94921 87716
rect 94535 87634 94582 87676
rect 94706 87634 94750 87676
rect 94874 87634 94921 87676
rect 109655 87716 109702 87758
rect 109826 87716 109870 87758
rect 109994 87716 110041 87758
rect 109655 87676 109664 87716
rect 109826 87676 109828 87716
rect 109868 87676 109870 87716
rect 110032 87676 110041 87716
rect 109655 87634 109702 87676
rect 109826 87634 109870 87676
rect 109994 87634 110041 87676
rect 124775 87716 124822 87758
rect 124946 87716 124990 87758
rect 125114 87716 125161 87758
rect 124775 87676 124784 87716
rect 124946 87676 124948 87716
rect 124988 87676 124990 87716
rect 125152 87676 125161 87716
rect 124775 87634 124822 87676
rect 124946 87634 124990 87676
rect 125114 87634 125161 87676
rect 139895 87716 139942 87758
rect 140066 87716 140110 87758
rect 140234 87716 140281 87758
rect 139895 87676 139904 87716
rect 140066 87676 140068 87716
rect 140108 87676 140110 87716
rect 140272 87676 140281 87716
rect 139895 87634 139942 87676
rect 140066 87634 140110 87676
rect 140234 87634 140281 87676
rect 78175 86960 78222 87002
rect 78346 86960 78390 87002
rect 78514 86960 78561 87002
rect 78175 86920 78184 86960
rect 78346 86920 78348 86960
rect 78388 86920 78390 86960
rect 78552 86920 78561 86960
rect 78175 86878 78222 86920
rect 78346 86878 78390 86920
rect 78514 86878 78561 86920
rect 93295 86960 93342 87002
rect 93466 86960 93510 87002
rect 93634 86960 93681 87002
rect 93295 86920 93304 86960
rect 93466 86920 93468 86960
rect 93508 86920 93510 86960
rect 93672 86920 93681 86960
rect 93295 86878 93342 86920
rect 93466 86878 93510 86920
rect 93634 86878 93681 86920
rect 108415 86960 108462 87002
rect 108586 86960 108630 87002
rect 108754 86960 108801 87002
rect 108415 86920 108424 86960
rect 108586 86920 108588 86960
rect 108628 86920 108630 86960
rect 108792 86920 108801 86960
rect 108415 86878 108462 86920
rect 108586 86878 108630 86920
rect 108754 86878 108801 86920
rect 123535 86960 123582 87002
rect 123706 86960 123750 87002
rect 123874 86960 123921 87002
rect 123535 86920 123544 86960
rect 123706 86920 123708 86960
rect 123748 86920 123750 86960
rect 123912 86920 123921 86960
rect 123535 86878 123582 86920
rect 123706 86878 123750 86920
rect 123874 86878 123921 86920
rect 138655 86960 138702 87002
rect 138826 86960 138870 87002
rect 138994 86960 139041 87002
rect 138655 86920 138664 86960
rect 138826 86920 138828 86960
rect 138868 86920 138870 86960
rect 139032 86920 139041 86960
rect 138655 86878 138702 86920
rect 138826 86878 138870 86920
rect 138994 86878 139041 86920
rect 79415 86204 79462 86246
rect 79586 86204 79630 86246
rect 79754 86204 79801 86246
rect 79415 86164 79424 86204
rect 79586 86164 79588 86204
rect 79628 86164 79630 86204
rect 79792 86164 79801 86204
rect 79415 86122 79462 86164
rect 79586 86122 79630 86164
rect 79754 86122 79801 86164
rect 94535 86204 94582 86246
rect 94706 86204 94750 86246
rect 94874 86204 94921 86246
rect 94535 86164 94544 86204
rect 94706 86164 94708 86204
rect 94748 86164 94750 86204
rect 94912 86164 94921 86204
rect 94535 86122 94582 86164
rect 94706 86122 94750 86164
rect 94874 86122 94921 86164
rect 109655 86204 109702 86246
rect 109826 86204 109870 86246
rect 109994 86204 110041 86246
rect 109655 86164 109664 86204
rect 109826 86164 109828 86204
rect 109868 86164 109870 86204
rect 110032 86164 110041 86204
rect 109655 86122 109702 86164
rect 109826 86122 109870 86164
rect 109994 86122 110041 86164
rect 124775 86204 124822 86246
rect 124946 86204 124990 86246
rect 125114 86204 125161 86246
rect 124775 86164 124784 86204
rect 124946 86164 124948 86204
rect 124988 86164 124990 86204
rect 125152 86164 125161 86204
rect 124775 86122 124822 86164
rect 124946 86122 124990 86164
rect 125114 86122 125161 86164
rect 139895 86204 139942 86246
rect 140066 86204 140110 86246
rect 140234 86204 140281 86246
rect 139895 86164 139904 86204
rect 140066 86164 140068 86204
rect 140108 86164 140110 86204
rect 140272 86164 140281 86204
rect 139895 86122 139942 86164
rect 140066 86122 140110 86164
rect 140234 86122 140281 86164
rect 78175 85448 78222 85490
rect 78346 85448 78390 85490
rect 78514 85448 78561 85490
rect 78175 85408 78184 85448
rect 78346 85408 78348 85448
rect 78388 85408 78390 85448
rect 78552 85408 78561 85448
rect 78175 85366 78222 85408
rect 78346 85366 78390 85408
rect 78514 85366 78561 85408
rect 93295 85448 93342 85490
rect 93466 85448 93510 85490
rect 93634 85448 93681 85490
rect 93295 85408 93304 85448
rect 93466 85408 93468 85448
rect 93508 85408 93510 85448
rect 93672 85408 93681 85448
rect 93295 85366 93342 85408
rect 93466 85366 93510 85408
rect 93634 85366 93681 85408
rect 108415 85448 108462 85490
rect 108586 85448 108630 85490
rect 108754 85448 108801 85490
rect 108415 85408 108424 85448
rect 108586 85408 108588 85448
rect 108628 85408 108630 85448
rect 108792 85408 108801 85448
rect 108415 85366 108462 85408
rect 108586 85366 108630 85408
rect 108754 85366 108801 85408
rect 123535 85448 123582 85490
rect 123706 85448 123750 85490
rect 123874 85448 123921 85490
rect 123535 85408 123544 85448
rect 123706 85408 123708 85448
rect 123748 85408 123750 85448
rect 123912 85408 123921 85448
rect 123535 85366 123582 85408
rect 123706 85366 123750 85408
rect 123874 85366 123921 85408
rect 138655 85448 138702 85490
rect 138826 85448 138870 85490
rect 138994 85448 139041 85490
rect 138655 85408 138664 85448
rect 138826 85408 138828 85448
rect 138868 85408 138870 85448
rect 139032 85408 139041 85448
rect 138655 85366 138702 85408
rect 138826 85366 138870 85408
rect 138994 85366 139041 85408
rect 79415 84692 79462 84734
rect 79586 84692 79630 84734
rect 79754 84692 79801 84734
rect 79415 84652 79424 84692
rect 79586 84652 79588 84692
rect 79628 84652 79630 84692
rect 79792 84652 79801 84692
rect 79415 84610 79462 84652
rect 79586 84610 79630 84652
rect 79754 84610 79801 84652
rect 94535 84692 94582 84734
rect 94706 84692 94750 84734
rect 94874 84692 94921 84734
rect 94535 84652 94544 84692
rect 94706 84652 94708 84692
rect 94748 84652 94750 84692
rect 94912 84652 94921 84692
rect 94535 84610 94582 84652
rect 94706 84610 94750 84652
rect 94874 84610 94921 84652
rect 109655 84692 109702 84734
rect 109826 84692 109870 84734
rect 109994 84692 110041 84734
rect 109655 84652 109664 84692
rect 109826 84652 109828 84692
rect 109868 84652 109870 84692
rect 110032 84652 110041 84692
rect 109655 84610 109702 84652
rect 109826 84610 109870 84652
rect 109994 84610 110041 84652
rect 124775 84692 124822 84734
rect 124946 84692 124990 84734
rect 125114 84692 125161 84734
rect 124775 84652 124784 84692
rect 124946 84652 124948 84692
rect 124988 84652 124990 84692
rect 125152 84652 125161 84692
rect 124775 84610 124822 84652
rect 124946 84610 124990 84652
rect 125114 84610 125161 84652
rect 139895 84692 139942 84734
rect 140066 84692 140110 84734
rect 140234 84692 140281 84734
rect 139895 84652 139904 84692
rect 140066 84652 140068 84692
rect 140108 84652 140110 84692
rect 140272 84652 140281 84692
rect 139895 84610 139942 84652
rect 140066 84610 140110 84652
rect 140234 84610 140281 84652
rect 78175 83936 78222 83978
rect 78346 83936 78390 83978
rect 78514 83936 78561 83978
rect 78175 83896 78184 83936
rect 78346 83896 78348 83936
rect 78388 83896 78390 83936
rect 78552 83896 78561 83936
rect 78175 83854 78222 83896
rect 78346 83854 78390 83896
rect 78514 83854 78561 83896
rect 93295 83936 93342 83978
rect 93466 83936 93510 83978
rect 93634 83936 93681 83978
rect 93295 83896 93304 83936
rect 93466 83896 93468 83936
rect 93508 83896 93510 83936
rect 93672 83896 93681 83936
rect 93295 83854 93342 83896
rect 93466 83854 93510 83896
rect 93634 83854 93681 83896
rect 108415 83936 108462 83978
rect 108586 83936 108630 83978
rect 108754 83936 108801 83978
rect 108415 83896 108424 83936
rect 108586 83896 108588 83936
rect 108628 83896 108630 83936
rect 108792 83896 108801 83936
rect 108415 83854 108462 83896
rect 108586 83854 108630 83896
rect 108754 83854 108801 83896
rect 123535 83936 123582 83978
rect 123706 83936 123750 83978
rect 123874 83936 123921 83978
rect 123535 83896 123544 83936
rect 123706 83896 123708 83936
rect 123748 83896 123750 83936
rect 123912 83896 123921 83936
rect 123535 83854 123582 83896
rect 123706 83854 123750 83896
rect 123874 83854 123921 83896
rect 138655 83936 138702 83978
rect 138826 83936 138870 83978
rect 138994 83936 139041 83978
rect 138655 83896 138664 83936
rect 138826 83896 138828 83936
rect 138868 83896 138870 83936
rect 139032 83896 139041 83936
rect 138655 83854 138702 83896
rect 138826 83854 138870 83896
rect 138994 83854 139041 83896
rect 79415 83180 79462 83222
rect 79586 83180 79630 83222
rect 79754 83180 79801 83222
rect 79415 83140 79424 83180
rect 79586 83140 79588 83180
rect 79628 83140 79630 83180
rect 79792 83140 79801 83180
rect 79415 83098 79462 83140
rect 79586 83098 79630 83140
rect 79754 83098 79801 83140
rect 94535 83180 94582 83222
rect 94706 83180 94750 83222
rect 94874 83180 94921 83222
rect 94535 83140 94544 83180
rect 94706 83140 94708 83180
rect 94748 83140 94750 83180
rect 94912 83140 94921 83180
rect 94535 83098 94582 83140
rect 94706 83098 94750 83140
rect 94874 83098 94921 83140
rect 109655 83180 109702 83222
rect 109826 83180 109870 83222
rect 109994 83180 110041 83222
rect 109655 83140 109664 83180
rect 109826 83140 109828 83180
rect 109868 83140 109870 83180
rect 110032 83140 110041 83180
rect 109655 83098 109702 83140
rect 109826 83098 109870 83140
rect 109994 83098 110041 83140
rect 124775 83180 124822 83222
rect 124946 83180 124990 83222
rect 125114 83180 125161 83222
rect 124775 83140 124784 83180
rect 124946 83140 124948 83180
rect 124988 83140 124990 83180
rect 125152 83140 125161 83180
rect 124775 83098 124822 83140
rect 124946 83098 124990 83140
rect 125114 83098 125161 83140
rect 139895 83180 139942 83222
rect 140066 83180 140110 83222
rect 140234 83180 140281 83222
rect 139895 83140 139904 83180
rect 140066 83140 140068 83180
rect 140108 83140 140110 83180
rect 140272 83140 140281 83180
rect 139895 83098 139942 83140
rect 140066 83098 140110 83140
rect 140234 83098 140281 83140
rect 78175 82424 78222 82466
rect 78346 82424 78390 82466
rect 78514 82424 78561 82466
rect 78175 82384 78184 82424
rect 78346 82384 78348 82424
rect 78388 82384 78390 82424
rect 78552 82384 78561 82424
rect 78175 82342 78222 82384
rect 78346 82342 78390 82384
rect 78514 82342 78561 82384
rect 93295 82424 93342 82466
rect 93466 82424 93510 82466
rect 93634 82424 93681 82466
rect 93295 82384 93304 82424
rect 93466 82384 93468 82424
rect 93508 82384 93510 82424
rect 93672 82384 93681 82424
rect 93295 82342 93342 82384
rect 93466 82342 93510 82384
rect 93634 82342 93681 82384
rect 108415 82424 108462 82466
rect 108586 82424 108630 82466
rect 108754 82424 108801 82466
rect 108415 82384 108424 82424
rect 108586 82384 108588 82424
rect 108628 82384 108630 82424
rect 108792 82384 108801 82424
rect 108415 82342 108462 82384
rect 108586 82342 108630 82384
rect 108754 82342 108801 82384
rect 123535 82424 123582 82466
rect 123706 82424 123750 82466
rect 123874 82424 123921 82466
rect 123535 82384 123544 82424
rect 123706 82384 123708 82424
rect 123748 82384 123750 82424
rect 123912 82384 123921 82424
rect 123535 82342 123582 82384
rect 123706 82342 123750 82384
rect 123874 82342 123921 82384
rect 138655 82424 138702 82466
rect 138826 82424 138870 82466
rect 138994 82424 139041 82466
rect 138655 82384 138664 82424
rect 138826 82384 138828 82424
rect 138868 82384 138870 82424
rect 139032 82384 139041 82424
rect 138655 82342 138702 82384
rect 138826 82342 138870 82384
rect 138994 82342 139041 82384
rect 79415 81668 79462 81710
rect 79586 81668 79630 81710
rect 79754 81668 79801 81710
rect 79415 81628 79424 81668
rect 79586 81628 79588 81668
rect 79628 81628 79630 81668
rect 79792 81628 79801 81668
rect 79415 81586 79462 81628
rect 79586 81586 79630 81628
rect 79754 81586 79801 81628
rect 94535 81668 94582 81710
rect 94706 81668 94750 81710
rect 94874 81668 94921 81710
rect 94535 81628 94544 81668
rect 94706 81628 94708 81668
rect 94748 81628 94750 81668
rect 94912 81628 94921 81668
rect 94535 81586 94582 81628
rect 94706 81586 94750 81628
rect 94874 81586 94921 81628
rect 109655 81668 109702 81710
rect 109826 81668 109870 81710
rect 109994 81668 110041 81710
rect 109655 81628 109664 81668
rect 109826 81628 109828 81668
rect 109868 81628 109870 81668
rect 110032 81628 110041 81668
rect 109655 81586 109702 81628
rect 109826 81586 109870 81628
rect 109994 81586 110041 81628
rect 124775 81668 124822 81710
rect 124946 81668 124990 81710
rect 125114 81668 125161 81710
rect 124775 81628 124784 81668
rect 124946 81628 124948 81668
rect 124988 81628 124990 81668
rect 125152 81628 125161 81668
rect 124775 81586 124822 81628
rect 124946 81586 124990 81628
rect 125114 81586 125161 81628
rect 139895 81668 139942 81710
rect 140066 81668 140110 81710
rect 140234 81668 140281 81710
rect 139895 81628 139904 81668
rect 140066 81628 140068 81668
rect 140108 81628 140110 81668
rect 140272 81628 140281 81668
rect 139895 81586 139942 81628
rect 140066 81586 140110 81628
rect 140234 81586 140281 81628
rect 78175 80912 78222 80954
rect 78346 80912 78390 80954
rect 78514 80912 78561 80954
rect 78175 80872 78184 80912
rect 78346 80872 78348 80912
rect 78388 80872 78390 80912
rect 78552 80872 78561 80912
rect 78175 80830 78222 80872
rect 78346 80830 78390 80872
rect 78514 80830 78561 80872
rect 93295 80912 93342 80954
rect 93466 80912 93510 80954
rect 93634 80912 93681 80954
rect 93295 80872 93304 80912
rect 93466 80872 93468 80912
rect 93508 80872 93510 80912
rect 93672 80872 93681 80912
rect 93295 80830 93342 80872
rect 93466 80830 93510 80872
rect 93634 80830 93681 80872
rect 108415 80912 108462 80954
rect 108586 80912 108630 80954
rect 108754 80912 108801 80954
rect 108415 80872 108424 80912
rect 108586 80872 108588 80912
rect 108628 80872 108630 80912
rect 108792 80872 108801 80912
rect 108415 80830 108462 80872
rect 108586 80830 108630 80872
rect 108754 80830 108801 80872
rect 123535 80912 123582 80954
rect 123706 80912 123750 80954
rect 123874 80912 123921 80954
rect 123535 80872 123544 80912
rect 123706 80872 123708 80912
rect 123748 80872 123750 80912
rect 123912 80872 123921 80912
rect 123535 80830 123582 80872
rect 123706 80830 123750 80872
rect 123874 80830 123921 80872
rect 138655 80912 138702 80954
rect 138826 80912 138870 80954
rect 138994 80912 139041 80954
rect 138655 80872 138664 80912
rect 138826 80872 138828 80912
rect 138868 80872 138870 80912
rect 139032 80872 139041 80912
rect 138655 80830 138702 80872
rect 138826 80830 138870 80872
rect 138994 80830 139041 80872
rect 79415 80156 79462 80198
rect 79586 80156 79630 80198
rect 79754 80156 79801 80198
rect 79415 80116 79424 80156
rect 79586 80116 79588 80156
rect 79628 80116 79630 80156
rect 79792 80116 79801 80156
rect 79415 80074 79462 80116
rect 79586 80074 79630 80116
rect 79754 80074 79801 80116
rect 94535 80156 94582 80198
rect 94706 80156 94750 80198
rect 94874 80156 94921 80198
rect 94535 80116 94544 80156
rect 94706 80116 94708 80156
rect 94748 80116 94750 80156
rect 94912 80116 94921 80156
rect 94535 80074 94582 80116
rect 94706 80074 94750 80116
rect 94874 80074 94921 80116
rect 109655 80156 109702 80198
rect 109826 80156 109870 80198
rect 109994 80156 110041 80198
rect 109655 80116 109664 80156
rect 109826 80116 109828 80156
rect 109868 80116 109870 80156
rect 110032 80116 110041 80156
rect 109655 80074 109702 80116
rect 109826 80074 109870 80116
rect 109994 80074 110041 80116
rect 124775 80156 124822 80198
rect 124946 80156 124990 80198
rect 125114 80156 125161 80198
rect 124775 80116 124784 80156
rect 124946 80116 124948 80156
rect 124988 80116 124990 80156
rect 125152 80116 125161 80156
rect 124775 80074 124822 80116
rect 124946 80074 124990 80116
rect 125114 80074 125161 80116
rect 139895 80156 139942 80198
rect 140066 80156 140110 80198
rect 140234 80156 140281 80198
rect 139895 80116 139904 80156
rect 140066 80116 140068 80156
rect 140108 80116 140110 80156
rect 140272 80116 140281 80156
rect 139895 80074 139942 80116
rect 140066 80074 140110 80116
rect 140234 80074 140281 80116
rect 78175 79400 78222 79442
rect 78346 79400 78390 79442
rect 78514 79400 78561 79442
rect 78175 79360 78184 79400
rect 78346 79360 78348 79400
rect 78388 79360 78390 79400
rect 78552 79360 78561 79400
rect 78175 79318 78222 79360
rect 78346 79318 78390 79360
rect 78514 79318 78561 79360
rect 93295 79400 93342 79442
rect 93466 79400 93510 79442
rect 93634 79400 93681 79442
rect 93295 79360 93304 79400
rect 93466 79360 93468 79400
rect 93508 79360 93510 79400
rect 93672 79360 93681 79400
rect 93295 79318 93342 79360
rect 93466 79318 93510 79360
rect 93634 79318 93681 79360
rect 108415 79400 108462 79442
rect 108586 79400 108630 79442
rect 108754 79400 108801 79442
rect 108415 79360 108424 79400
rect 108586 79360 108588 79400
rect 108628 79360 108630 79400
rect 108792 79360 108801 79400
rect 108415 79318 108462 79360
rect 108586 79318 108630 79360
rect 108754 79318 108801 79360
rect 123535 79400 123582 79442
rect 123706 79400 123750 79442
rect 123874 79400 123921 79442
rect 123535 79360 123544 79400
rect 123706 79360 123708 79400
rect 123748 79360 123750 79400
rect 123912 79360 123921 79400
rect 123535 79318 123582 79360
rect 123706 79318 123750 79360
rect 123874 79318 123921 79360
rect 138655 79400 138702 79442
rect 138826 79400 138870 79442
rect 138994 79400 139041 79442
rect 138655 79360 138664 79400
rect 138826 79360 138828 79400
rect 138868 79360 138870 79400
rect 139032 79360 139041 79400
rect 138655 79318 138702 79360
rect 138826 79318 138870 79360
rect 138994 79318 139041 79360
rect 79415 78644 79462 78686
rect 79586 78644 79630 78686
rect 79754 78644 79801 78686
rect 79415 78604 79424 78644
rect 79586 78604 79588 78644
rect 79628 78604 79630 78644
rect 79792 78604 79801 78644
rect 79415 78562 79462 78604
rect 79586 78562 79630 78604
rect 79754 78562 79801 78604
rect 94535 78644 94582 78686
rect 94706 78644 94750 78686
rect 94874 78644 94921 78686
rect 94535 78604 94544 78644
rect 94706 78604 94708 78644
rect 94748 78604 94750 78644
rect 94912 78604 94921 78644
rect 94535 78562 94582 78604
rect 94706 78562 94750 78604
rect 94874 78562 94921 78604
rect 109655 78644 109702 78686
rect 109826 78644 109870 78686
rect 109994 78644 110041 78686
rect 109655 78604 109664 78644
rect 109826 78604 109828 78644
rect 109868 78604 109870 78644
rect 110032 78604 110041 78644
rect 109655 78562 109702 78604
rect 109826 78562 109870 78604
rect 109994 78562 110041 78604
rect 124775 78644 124822 78686
rect 124946 78644 124990 78686
rect 125114 78644 125161 78686
rect 124775 78604 124784 78644
rect 124946 78604 124948 78644
rect 124988 78604 124990 78644
rect 125152 78604 125161 78644
rect 124775 78562 124822 78604
rect 124946 78562 124990 78604
rect 125114 78562 125161 78604
rect 139895 78644 139942 78686
rect 140066 78644 140110 78686
rect 140234 78644 140281 78686
rect 139895 78604 139904 78644
rect 140066 78604 140068 78644
rect 140108 78604 140110 78644
rect 140272 78604 140281 78644
rect 139895 78562 139942 78604
rect 140066 78562 140110 78604
rect 140234 78562 140281 78604
rect 78175 77888 78222 77930
rect 78346 77888 78390 77930
rect 78514 77888 78561 77930
rect 78175 77848 78184 77888
rect 78346 77848 78348 77888
rect 78388 77848 78390 77888
rect 78552 77848 78561 77888
rect 78175 77806 78222 77848
rect 78346 77806 78390 77848
rect 78514 77806 78561 77848
rect 93295 77888 93342 77930
rect 93466 77888 93510 77930
rect 93634 77888 93681 77930
rect 93295 77848 93304 77888
rect 93466 77848 93468 77888
rect 93508 77848 93510 77888
rect 93672 77848 93681 77888
rect 93295 77806 93342 77848
rect 93466 77806 93510 77848
rect 93634 77806 93681 77848
rect 108415 77888 108462 77930
rect 108586 77888 108630 77930
rect 108754 77888 108801 77930
rect 108415 77848 108424 77888
rect 108586 77848 108588 77888
rect 108628 77848 108630 77888
rect 108792 77848 108801 77888
rect 108415 77806 108462 77848
rect 108586 77806 108630 77848
rect 108754 77806 108801 77848
rect 123535 77888 123582 77930
rect 123706 77888 123750 77930
rect 123874 77888 123921 77930
rect 123535 77848 123544 77888
rect 123706 77848 123708 77888
rect 123748 77848 123750 77888
rect 123912 77848 123921 77888
rect 123535 77806 123582 77848
rect 123706 77806 123750 77848
rect 123874 77806 123921 77848
rect 138655 77888 138702 77930
rect 138826 77888 138870 77930
rect 138994 77888 139041 77930
rect 138655 77848 138664 77888
rect 138826 77848 138828 77888
rect 138868 77848 138870 77888
rect 139032 77848 139041 77888
rect 138655 77806 138702 77848
rect 138826 77806 138870 77848
rect 138994 77806 139041 77848
rect 79415 77132 79462 77174
rect 79586 77132 79630 77174
rect 79754 77132 79801 77174
rect 79415 77092 79424 77132
rect 79586 77092 79588 77132
rect 79628 77092 79630 77132
rect 79792 77092 79801 77132
rect 79415 77050 79462 77092
rect 79586 77050 79630 77092
rect 79754 77050 79801 77092
rect 94535 77132 94582 77174
rect 94706 77132 94750 77174
rect 94874 77132 94921 77174
rect 94535 77092 94544 77132
rect 94706 77092 94708 77132
rect 94748 77092 94750 77132
rect 94912 77092 94921 77132
rect 94535 77050 94582 77092
rect 94706 77050 94750 77092
rect 94874 77050 94921 77092
rect 109655 77132 109702 77174
rect 109826 77132 109870 77174
rect 109994 77132 110041 77174
rect 109655 77092 109664 77132
rect 109826 77092 109828 77132
rect 109868 77092 109870 77132
rect 110032 77092 110041 77132
rect 109655 77050 109702 77092
rect 109826 77050 109870 77092
rect 109994 77050 110041 77092
rect 124775 77132 124822 77174
rect 124946 77132 124990 77174
rect 125114 77132 125161 77174
rect 124775 77092 124784 77132
rect 124946 77092 124948 77132
rect 124988 77092 124990 77132
rect 125152 77092 125161 77132
rect 124775 77050 124822 77092
rect 124946 77050 124990 77092
rect 125114 77050 125161 77092
rect 139895 77132 139942 77174
rect 140066 77132 140110 77174
rect 140234 77132 140281 77174
rect 139895 77092 139904 77132
rect 140066 77092 140068 77132
rect 140108 77092 140110 77132
rect 140272 77092 140281 77132
rect 139895 77050 139942 77092
rect 140066 77050 140110 77092
rect 140234 77050 140281 77092
rect 78175 76376 78222 76418
rect 78346 76376 78390 76418
rect 78514 76376 78561 76418
rect 78175 76336 78184 76376
rect 78346 76336 78348 76376
rect 78388 76336 78390 76376
rect 78552 76336 78561 76376
rect 78175 76294 78222 76336
rect 78346 76294 78390 76336
rect 78514 76294 78561 76336
rect 93295 76376 93342 76418
rect 93466 76376 93510 76418
rect 93634 76376 93681 76418
rect 93295 76336 93304 76376
rect 93466 76336 93468 76376
rect 93508 76336 93510 76376
rect 93672 76336 93681 76376
rect 93295 76294 93342 76336
rect 93466 76294 93510 76336
rect 93634 76294 93681 76336
rect 108415 76376 108462 76418
rect 108586 76376 108630 76418
rect 108754 76376 108801 76418
rect 108415 76336 108424 76376
rect 108586 76336 108588 76376
rect 108628 76336 108630 76376
rect 108792 76336 108801 76376
rect 108415 76294 108462 76336
rect 108586 76294 108630 76336
rect 108754 76294 108801 76336
rect 123535 76376 123582 76418
rect 123706 76376 123750 76418
rect 123874 76376 123921 76418
rect 123535 76336 123544 76376
rect 123706 76336 123708 76376
rect 123748 76336 123750 76376
rect 123912 76336 123921 76376
rect 123535 76294 123582 76336
rect 123706 76294 123750 76336
rect 123874 76294 123921 76336
rect 138655 76376 138702 76418
rect 138826 76376 138870 76418
rect 138994 76376 139041 76418
rect 138655 76336 138664 76376
rect 138826 76336 138828 76376
rect 138868 76336 138870 76376
rect 139032 76336 139041 76376
rect 138655 76294 138702 76336
rect 138826 76294 138870 76336
rect 138994 76294 139041 76336
rect 79415 75620 79462 75662
rect 79586 75620 79630 75662
rect 79754 75620 79801 75662
rect 79415 75580 79424 75620
rect 79586 75580 79588 75620
rect 79628 75580 79630 75620
rect 79792 75580 79801 75620
rect 79415 75538 79462 75580
rect 79586 75538 79630 75580
rect 79754 75538 79801 75580
rect 94535 75620 94582 75662
rect 94706 75620 94750 75662
rect 94874 75620 94921 75662
rect 94535 75580 94544 75620
rect 94706 75580 94708 75620
rect 94748 75580 94750 75620
rect 94912 75580 94921 75620
rect 94535 75538 94582 75580
rect 94706 75538 94750 75580
rect 94874 75538 94921 75580
rect 109655 75620 109702 75662
rect 109826 75620 109870 75662
rect 109994 75620 110041 75662
rect 109655 75580 109664 75620
rect 109826 75580 109828 75620
rect 109868 75580 109870 75620
rect 110032 75580 110041 75620
rect 109655 75538 109702 75580
rect 109826 75538 109870 75580
rect 109994 75538 110041 75580
rect 124775 75620 124822 75662
rect 124946 75620 124990 75662
rect 125114 75620 125161 75662
rect 124775 75580 124784 75620
rect 124946 75580 124948 75620
rect 124988 75580 124990 75620
rect 125152 75580 125161 75620
rect 124775 75538 124822 75580
rect 124946 75538 124990 75580
rect 125114 75538 125161 75580
rect 139895 75620 139942 75662
rect 140066 75620 140110 75662
rect 140234 75620 140281 75662
rect 139895 75580 139904 75620
rect 140066 75580 140068 75620
rect 140108 75580 140110 75620
rect 140272 75580 140281 75620
rect 139895 75538 139942 75580
rect 140066 75538 140110 75580
rect 140234 75538 140281 75580
rect 90691 71212 90700 71252
rect 90740 71212 92140 71252
rect 92180 71212 92189 71252
<< via5 >>
rect 79462 148196 79586 148238
rect 79630 148196 79754 148238
rect 79462 148156 79464 148196
rect 79464 148156 79506 148196
rect 79506 148156 79546 148196
rect 79546 148156 79586 148196
rect 79630 148156 79670 148196
rect 79670 148156 79710 148196
rect 79710 148156 79752 148196
rect 79752 148156 79754 148196
rect 79462 148114 79586 148156
rect 79630 148114 79754 148156
rect 94582 148196 94706 148238
rect 94750 148196 94874 148238
rect 94582 148156 94584 148196
rect 94584 148156 94626 148196
rect 94626 148156 94666 148196
rect 94666 148156 94706 148196
rect 94750 148156 94790 148196
rect 94790 148156 94830 148196
rect 94830 148156 94872 148196
rect 94872 148156 94874 148196
rect 94582 148114 94706 148156
rect 94750 148114 94874 148156
rect 109702 148196 109826 148238
rect 109870 148196 109994 148238
rect 109702 148156 109704 148196
rect 109704 148156 109746 148196
rect 109746 148156 109786 148196
rect 109786 148156 109826 148196
rect 109870 148156 109910 148196
rect 109910 148156 109950 148196
rect 109950 148156 109992 148196
rect 109992 148156 109994 148196
rect 109702 148114 109826 148156
rect 109870 148114 109994 148156
rect 124822 148196 124946 148238
rect 124990 148196 125114 148238
rect 124822 148156 124824 148196
rect 124824 148156 124866 148196
rect 124866 148156 124906 148196
rect 124906 148156 124946 148196
rect 124990 148156 125030 148196
rect 125030 148156 125070 148196
rect 125070 148156 125112 148196
rect 125112 148156 125114 148196
rect 124822 148114 124946 148156
rect 124990 148114 125114 148156
rect 139942 148196 140066 148238
rect 140110 148196 140234 148238
rect 139942 148156 139944 148196
rect 139944 148156 139986 148196
rect 139986 148156 140026 148196
rect 140026 148156 140066 148196
rect 140110 148156 140150 148196
rect 140150 148156 140190 148196
rect 140190 148156 140232 148196
rect 140232 148156 140234 148196
rect 139942 148114 140066 148156
rect 140110 148114 140234 148156
rect 78222 147440 78346 147482
rect 78390 147440 78514 147482
rect 78222 147400 78224 147440
rect 78224 147400 78266 147440
rect 78266 147400 78306 147440
rect 78306 147400 78346 147440
rect 78390 147400 78430 147440
rect 78430 147400 78470 147440
rect 78470 147400 78512 147440
rect 78512 147400 78514 147440
rect 78222 147358 78346 147400
rect 78390 147358 78514 147400
rect 93342 147440 93466 147482
rect 93510 147440 93634 147482
rect 93342 147400 93344 147440
rect 93344 147400 93386 147440
rect 93386 147400 93426 147440
rect 93426 147400 93466 147440
rect 93510 147400 93550 147440
rect 93550 147400 93590 147440
rect 93590 147400 93632 147440
rect 93632 147400 93634 147440
rect 93342 147358 93466 147400
rect 93510 147358 93634 147400
rect 108462 147440 108586 147482
rect 108630 147440 108754 147482
rect 108462 147400 108464 147440
rect 108464 147400 108506 147440
rect 108506 147400 108546 147440
rect 108546 147400 108586 147440
rect 108630 147400 108670 147440
rect 108670 147400 108710 147440
rect 108710 147400 108752 147440
rect 108752 147400 108754 147440
rect 108462 147358 108586 147400
rect 108630 147358 108754 147400
rect 123582 147440 123706 147482
rect 123750 147440 123874 147482
rect 123582 147400 123584 147440
rect 123584 147400 123626 147440
rect 123626 147400 123666 147440
rect 123666 147400 123706 147440
rect 123750 147400 123790 147440
rect 123790 147400 123830 147440
rect 123830 147400 123872 147440
rect 123872 147400 123874 147440
rect 123582 147358 123706 147400
rect 123750 147358 123874 147400
rect 138702 147440 138826 147482
rect 138870 147440 138994 147482
rect 138702 147400 138704 147440
rect 138704 147400 138746 147440
rect 138746 147400 138786 147440
rect 138786 147400 138826 147440
rect 138870 147400 138910 147440
rect 138910 147400 138950 147440
rect 138950 147400 138992 147440
rect 138992 147400 138994 147440
rect 138702 147358 138826 147400
rect 138870 147358 138994 147400
rect 79462 146684 79586 146726
rect 79630 146684 79754 146726
rect 79462 146644 79464 146684
rect 79464 146644 79506 146684
rect 79506 146644 79546 146684
rect 79546 146644 79586 146684
rect 79630 146644 79670 146684
rect 79670 146644 79710 146684
rect 79710 146644 79752 146684
rect 79752 146644 79754 146684
rect 79462 146602 79586 146644
rect 79630 146602 79754 146644
rect 94582 146684 94706 146726
rect 94750 146684 94874 146726
rect 94582 146644 94584 146684
rect 94584 146644 94626 146684
rect 94626 146644 94666 146684
rect 94666 146644 94706 146684
rect 94750 146644 94790 146684
rect 94790 146644 94830 146684
rect 94830 146644 94872 146684
rect 94872 146644 94874 146684
rect 94582 146602 94706 146644
rect 94750 146602 94874 146644
rect 109702 146684 109826 146726
rect 109870 146684 109994 146726
rect 109702 146644 109704 146684
rect 109704 146644 109746 146684
rect 109746 146644 109786 146684
rect 109786 146644 109826 146684
rect 109870 146644 109910 146684
rect 109910 146644 109950 146684
rect 109950 146644 109992 146684
rect 109992 146644 109994 146684
rect 109702 146602 109826 146644
rect 109870 146602 109994 146644
rect 124822 146684 124946 146726
rect 124990 146684 125114 146726
rect 124822 146644 124824 146684
rect 124824 146644 124866 146684
rect 124866 146644 124906 146684
rect 124906 146644 124946 146684
rect 124990 146644 125030 146684
rect 125030 146644 125070 146684
rect 125070 146644 125112 146684
rect 125112 146644 125114 146684
rect 124822 146602 124946 146644
rect 124990 146602 125114 146644
rect 139942 146684 140066 146726
rect 140110 146684 140234 146726
rect 139942 146644 139944 146684
rect 139944 146644 139986 146684
rect 139986 146644 140026 146684
rect 140026 146644 140066 146684
rect 140110 146644 140150 146684
rect 140150 146644 140190 146684
rect 140190 146644 140232 146684
rect 140232 146644 140234 146684
rect 139942 146602 140066 146644
rect 140110 146602 140234 146644
rect 78222 145928 78346 145970
rect 78390 145928 78514 145970
rect 78222 145888 78224 145928
rect 78224 145888 78266 145928
rect 78266 145888 78306 145928
rect 78306 145888 78346 145928
rect 78390 145888 78430 145928
rect 78430 145888 78470 145928
rect 78470 145888 78512 145928
rect 78512 145888 78514 145928
rect 78222 145846 78346 145888
rect 78390 145846 78514 145888
rect 93342 145928 93466 145970
rect 93510 145928 93634 145970
rect 93342 145888 93344 145928
rect 93344 145888 93386 145928
rect 93386 145888 93426 145928
rect 93426 145888 93466 145928
rect 93510 145888 93550 145928
rect 93550 145888 93590 145928
rect 93590 145888 93632 145928
rect 93632 145888 93634 145928
rect 93342 145846 93466 145888
rect 93510 145846 93634 145888
rect 108462 145928 108586 145970
rect 108630 145928 108754 145970
rect 108462 145888 108464 145928
rect 108464 145888 108506 145928
rect 108506 145888 108546 145928
rect 108546 145888 108586 145928
rect 108630 145888 108670 145928
rect 108670 145888 108710 145928
rect 108710 145888 108752 145928
rect 108752 145888 108754 145928
rect 108462 145846 108586 145888
rect 108630 145846 108754 145888
rect 123582 145928 123706 145970
rect 123750 145928 123874 145970
rect 123582 145888 123584 145928
rect 123584 145888 123626 145928
rect 123626 145888 123666 145928
rect 123666 145888 123706 145928
rect 123750 145888 123790 145928
rect 123790 145888 123830 145928
rect 123830 145888 123872 145928
rect 123872 145888 123874 145928
rect 123582 145846 123706 145888
rect 123750 145846 123874 145888
rect 138702 145928 138826 145970
rect 138870 145928 138994 145970
rect 138702 145888 138704 145928
rect 138704 145888 138746 145928
rect 138746 145888 138786 145928
rect 138786 145888 138826 145928
rect 138870 145888 138910 145928
rect 138910 145888 138950 145928
rect 138950 145888 138992 145928
rect 138992 145888 138994 145928
rect 138702 145846 138826 145888
rect 138870 145846 138994 145888
rect 79462 145172 79586 145214
rect 79630 145172 79754 145214
rect 79462 145132 79464 145172
rect 79464 145132 79506 145172
rect 79506 145132 79546 145172
rect 79546 145132 79586 145172
rect 79630 145132 79670 145172
rect 79670 145132 79710 145172
rect 79710 145132 79752 145172
rect 79752 145132 79754 145172
rect 79462 145090 79586 145132
rect 79630 145090 79754 145132
rect 94582 145172 94706 145214
rect 94750 145172 94874 145214
rect 94582 145132 94584 145172
rect 94584 145132 94626 145172
rect 94626 145132 94666 145172
rect 94666 145132 94706 145172
rect 94750 145132 94790 145172
rect 94790 145132 94830 145172
rect 94830 145132 94872 145172
rect 94872 145132 94874 145172
rect 94582 145090 94706 145132
rect 94750 145090 94874 145132
rect 109702 145172 109826 145214
rect 109870 145172 109994 145214
rect 109702 145132 109704 145172
rect 109704 145132 109746 145172
rect 109746 145132 109786 145172
rect 109786 145132 109826 145172
rect 109870 145132 109910 145172
rect 109910 145132 109950 145172
rect 109950 145132 109992 145172
rect 109992 145132 109994 145172
rect 109702 145090 109826 145132
rect 109870 145090 109994 145132
rect 124822 145172 124946 145214
rect 124990 145172 125114 145214
rect 124822 145132 124824 145172
rect 124824 145132 124866 145172
rect 124866 145132 124906 145172
rect 124906 145132 124946 145172
rect 124990 145132 125030 145172
rect 125030 145132 125070 145172
rect 125070 145132 125112 145172
rect 125112 145132 125114 145172
rect 124822 145090 124946 145132
rect 124990 145090 125114 145132
rect 139942 145172 140066 145214
rect 140110 145172 140234 145214
rect 139942 145132 139944 145172
rect 139944 145132 139986 145172
rect 139986 145132 140026 145172
rect 140026 145132 140066 145172
rect 140110 145132 140150 145172
rect 140150 145132 140190 145172
rect 140190 145132 140232 145172
rect 140232 145132 140234 145172
rect 139942 145090 140066 145132
rect 140110 145090 140234 145132
rect 78222 144416 78346 144458
rect 78390 144416 78514 144458
rect 78222 144376 78224 144416
rect 78224 144376 78266 144416
rect 78266 144376 78306 144416
rect 78306 144376 78346 144416
rect 78390 144376 78430 144416
rect 78430 144376 78470 144416
rect 78470 144376 78512 144416
rect 78512 144376 78514 144416
rect 78222 144334 78346 144376
rect 78390 144334 78514 144376
rect 93342 144416 93466 144458
rect 93510 144416 93634 144458
rect 93342 144376 93344 144416
rect 93344 144376 93386 144416
rect 93386 144376 93426 144416
rect 93426 144376 93466 144416
rect 93510 144376 93550 144416
rect 93550 144376 93590 144416
rect 93590 144376 93632 144416
rect 93632 144376 93634 144416
rect 93342 144334 93466 144376
rect 93510 144334 93634 144376
rect 108462 144416 108586 144458
rect 108630 144416 108754 144458
rect 108462 144376 108464 144416
rect 108464 144376 108506 144416
rect 108506 144376 108546 144416
rect 108546 144376 108586 144416
rect 108630 144376 108670 144416
rect 108670 144376 108710 144416
rect 108710 144376 108752 144416
rect 108752 144376 108754 144416
rect 108462 144334 108586 144376
rect 108630 144334 108754 144376
rect 123582 144416 123706 144458
rect 123750 144416 123874 144458
rect 123582 144376 123584 144416
rect 123584 144376 123626 144416
rect 123626 144376 123666 144416
rect 123666 144376 123706 144416
rect 123750 144376 123790 144416
rect 123790 144376 123830 144416
rect 123830 144376 123872 144416
rect 123872 144376 123874 144416
rect 123582 144334 123706 144376
rect 123750 144334 123874 144376
rect 138702 144416 138826 144458
rect 138870 144416 138994 144458
rect 138702 144376 138704 144416
rect 138704 144376 138746 144416
rect 138746 144376 138786 144416
rect 138786 144376 138826 144416
rect 138870 144376 138910 144416
rect 138910 144376 138950 144416
rect 138950 144376 138992 144416
rect 138992 144376 138994 144416
rect 138702 144334 138826 144376
rect 138870 144334 138994 144376
rect 79462 143660 79586 143702
rect 79630 143660 79754 143702
rect 79462 143620 79464 143660
rect 79464 143620 79506 143660
rect 79506 143620 79546 143660
rect 79546 143620 79586 143660
rect 79630 143620 79670 143660
rect 79670 143620 79710 143660
rect 79710 143620 79752 143660
rect 79752 143620 79754 143660
rect 79462 143578 79586 143620
rect 79630 143578 79754 143620
rect 94582 143660 94706 143702
rect 94750 143660 94874 143702
rect 94582 143620 94584 143660
rect 94584 143620 94626 143660
rect 94626 143620 94666 143660
rect 94666 143620 94706 143660
rect 94750 143620 94790 143660
rect 94790 143620 94830 143660
rect 94830 143620 94872 143660
rect 94872 143620 94874 143660
rect 94582 143578 94706 143620
rect 94750 143578 94874 143620
rect 109702 143660 109826 143702
rect 109870 143660 109994 143702
rect 109702 143620 109704 143660
rect 109704 143620 109746 143660
rect 109746 143620 109786 143660
rect 109786 143620 109826 143660
rect 109870 143620 109910 143660
rect 109910 143620 109950 143660
rect 109950 143620 109992 143660
rect 109992 143620 109994 143660
rect 109702 143578 109826 143620
rect 109870 143578 109994 143620
rect 124822 143660 124946 143702
rect 124990 143660 125114 143702
rect 124822 143620 124824 143660
rect 124824 143620 124866 143660
rect 124866 143620 124906 143660
rect 124906 143620 124946 143660
rect 124990 143620 125030 143660
rect 125030 143620 125070 143660
rect 125070 143620 125112 143660
rect 125112 143620 125114 143660
rect 124822 143578 124946 143620
rect 124990 143578 125114 143620
rect 139942 143660 140066 143702
rect 140110 143660 140234 143702
rect 139942 143620 139944 143660
rect 139944 143620 139986 143660
rect 139986 143620 140026 143660
rect 140026 143620 140066 143660
rect 140110 143620 140150 143660
rect 140150 143620 140190 143660
rect 140190 143620 140232 143660
rect 140232 143620 140234 143660
rect 139942 143578 140066 143620
rect 140110 143578 140234 143620
rect 78222 142904 78346 142946
rect 78390 142904 78514 142946
rect 78222 142864 78224 142904
rect 78224 142864 78266 142904
rect 78266 142864 78306 142904
rect 78306 142864 78346 142904
rect 78390 142864 78430 142904
rect 78430 142864 78470 142904
rect 78470 142864 78512 142904
rect 78512 142864 78514 142904
rect 78222 142822 78346 142864
rect 78390 142822 78514 142864
rect 93342 142904 93466 142946
rect 93510 142904 93634 142946
rect 93342 142864 93344 142904
rect 93344 142864 93386 142904
rect 93386 142864 93426 142904
rect 93426 142864 93466 142904
rect 93510 142864 93550 142904
rect 93550 142864 93590 142904
rect 93590 142864 93632 142904
rect 93632 142864 93634 142904
rect 93342 142822 93466 142864
rect 93510 142822 93634 142864
rect 108462 142904 108586 142946
rect 108630 142904 108754 142946
rect 108462 142864 108464 142904
rect 108464 142864 108506 142904
rect 108506 142864 108546 142904
rect 108546 142864 108586 142904
rect 108630 142864 108670 142904
rect 108670 142864 108710 142904
rect 108710 142864 108752 142904
rect 108752 142864 108754 142904
rect 108462 142822 108586 142864
rect 108630 142822 108754 142864
rect 123582 142904 123706 142946
rect 123750 142904 123874 142946
rect 123582 142864 123584 142904
rect 123584 142864 123626 142904
rect 123626 142864 123666 142904
rect 123666 142864 123706 142904
rect 123750 142864 123790 142904
rect 123790 142864 123830 142904
rect 123830 142864 123872 142904
rect 123872 142864 123874 142904
rect 123582 142822 123706 142864
rect 123750 142822 123874 142864
rect 138702 142904 138826 142946
rect 138870 142904 138994 142946
rect 138702 142864 138704 142904
rect 138704 142864 138746 142904
rect 138746 142864 138786 142904
rect 138786 142864 138826 142904
rect 138870 142864 138910 142904
rect 138910 142864 138950 142904
rect 138950 142864 138992 142904
rect 138992 142864 138994 142904
rect 138702 142822 138826 142864
rect 138870 142822 138994 142864
rect 79462 142148 79586 142190
rect 79630 142148 79754 142190
rect 79462 142108 79464 142148
rect 79464 142108 79506 142148
rect 79506 142108 79546 142148
rect 79546 142108 79586 142148
rect 79630 142108 79670 142148
rect 79670 142108 79710 142148
rect 79710 142108 79752 142148
rect 79752 142108 79754 142148
rect 79462 142066 79586 142108
rect 79630 142066 79754 142108
rect 94582 142148 94706 142190
rect 94750 142148 94874 142190
rect 94582 142108 94584 142148
rect 94584 142108 94626 142148
rect 94626 142108 94666 142148
rect 94666 142108 94706 142148
rect 94750 142108 94790 142148
rect 94790 142108 94830 142148
rect 94830 142108 94872 142148
rect 94872 142108 94874 142148
rect 94582 142066 94706 142108
rect 94750 142066 94874 142108
rect 109702 142148 109826 142190
rect 109870 142148 109994 142190
rect 109702 142108 109704 142148
rect 109704 142108 109746 142148
rect 109746 142108 109786 142148
rect 109786 142108 109826 142148
rect 109870 142108 109910 142148
rect 109910 142108 109950 142148
rect 109950 142108 109992 142148
rect 109992 142108 109994 142148
rect 109702 142066 109826 142108
rect 109870 142066 109994 142108
rect 124822 142148 124946 142190
rect 124990 142148 125114 142190
rect 124822 142108 124824 142148
rect 124824 142108 124866 142148
rect 124866 142108 124906 142148
rect 124906 142108 124946 142148
rect 124990 142108 125030 142148
rect 125030 142108 125070 142148
rect 125070 142108 125112 142148
rect 125112 142108 125114 142148
rect 124822 142066 124946 142108
rect 124990 142066 125114 142108
rect 139942 142148 140066 142190
rect 140110 142148 140234 142190
rect 139942 142108 139944 142148
rect 139944 142108 139986 142148
rect 139986 142108 140026 142148
rect 140026 142108 140066 142148
rect 140110 142108 140150 142148
rect 140150 142108 140190 142148
rect 140190 142108 140232 142148
rect 140232 142108 140234 142148
rect 139942 142066 140066 142108
rect 140110 142066 140234 142108
rect 78222 141392 78346 141434
rect 78390 141392 78514 141434
rect 78222 141352 78224 141392
rect 78224 141352 78266 141392
rect 78266 141352 78306 141392
rect 78306 141352 78346 141392
rect 78390 141352 78430 141392
rect 78430 141352 78470 141392
rect 78470 141352 78512 141392
rect 78512 141352 78514 141392
rect 78222 141310 78346 141352
rect 78390 141310 78514 141352
rect 93342 141392 93466 141434
rect 93510 141392 93634 141434
rect 93342 141352 93344 141392
rect 93344 141352 93386 141392
rect 93386 141352 93426 141392
rect 93426 141352 93466 141392
rect 93510 141352 93550 141392
rect 93550 141352 93590 141392
rect 93590 141352 93632 141392
rect 93632 141352 93634 141392
rect 93342 141310 93466 141352
rect 93510 141310 93634 141352
rect 108462 141392 108586 141434
rect 108630 141392 108754 141434
rect 108462 141352 108464 141392
rect 108464 141352 108506 141392
rect 108506 141352 108546 141392
rect 108546 141352 108586 141392
rect 108630 141352 108670 141392
rect 108670 141352 108710 141392
rect 108710 141352 108752 141392
rect 108752 141352 108754 141392
rect 108462 141310 108586 141352
rect 108630 141310 108754 141352
rect 123582 141392 123706 141434
rect 123750 141392 123874 141434
rect 123582 141352 123584 141392
rect 123584 141352 123626 141392
rect 123626 141352 123666 141392
rect 123666 141352 123706 141392
rect 123750 141352 123790 141392
rect 123790 141352 123830 141392
rect 123830 141352 123872 141392
rect 123872 141352 123874 141392
rect 123582 141310 123706 141352
rect 123750 141310 123874 141352
rect 138702 141392 138826 141434
rect 138870 141392 138994 141434
rect 138702 141352 138704 141392
rect 138704 141352 138746 141392
rect 138746 141352 138786 141392
rect 138786 141352 138826 141392
rect 138870 141352 138910 141392
rect 138910 141352 138950 141392
rect 138950 141352 138992 141392
rect 138992 141352 138994 141392
rect 138702 141310 138826 141352
rect 138870 141310 138994 141352
rect 79462 140636 79586 140678
rect 79630 140636 79754 140678
rect 79462 140596 79464 140636
rect 79464 140596 79506 140636
rect 79506 140596 79546 140636
rect 79546 140596 79586 140636
rect 79630 140596 79670 140636
rect 79670 140596 79710 140636
rect 79710 140596 79752 140636
rect 79752 140596 79754 140636
rect 79462 140554 79586 140596
rect 79630 140554 79754 140596
rect 94582 140636 94706 140678
rect 94750 140636 94874 140678
rect 94582 140596 94584 140636
rect 94584 140596 94626 140636
rect 94626 140596 94666 140636
rect 94666 140596 94706 140636
rect 94750 140596 94790 140636
rect 94790 140596 94830 140636
rect 94830 140596 94872 140636
rect 94872 140596 94874 140636
rect 94582 140554 94706 140596
rect 94750 140554 94874 140596
rect 109702 140636 109826 140678
rect 109870 140636 109994 140678
rect 109702 140596 109704 140636
rect 109704 140596 109746 140636
rect 109746 140596 109786 140636
rect 109786 140596 109826 140636
rect 109870 140596 109910 140636
rect 109910 140596 109950 140636
rect 109950 140596 109992 140636
rect 109992 140596 109994 140636
rect 109702 140554 109826 140596
rect 109870 140554 109994 140596
rect 124822 140636 124946 140678
rect 124990 140636 125114 140678
rect 124822 140596 124824 140636
rect 124824 140596 124866 140636
rect 124866 140596 124906 140636
rect 124906 140596 124946 140636
rect 124990 140596 125030 140636
rect 125030 140596 125070 140636
rect 125070 140596 125112 140636
rect 125112 140596 125114 140636
rect 124822 140554 124946 140596
rect 124990 140554 125114 140596
rect 139942 140636 140066 140678
rect 140110 140636 140234 140678
rect 139942 140596 139944 140636
rect 139944 140596 139986 140636
rect 139986 140596 140026 140636
rect 140026 140596 140066 140636
rect 140110 140596 140150 140636
rect 140150 140596 140190 140636
rect 140190 140596 140232 140636
rect 140232 140596 140234 140636
rect 139942 140554 140066 140596
rect 140110 140554 140234 140596
rect 78222 139880 78346 139922
rect 78390 139880 78514 139922
rect 78222 139840 78224 139880
rect 78224 139840 78266 139880
rect 78266 139840 78306 139880
rect 78306 139840 78346 139880
rect 78390 139840 78430 139880
rect 78430 139840 78470 139880
rect 78470 139840 78512 139880
rect 78512 139840 78514 139880
rect 78222 139798 78346 139840
rect 78390 139798 78514 139840
rect 93342 139880 93466 139922
rect 93510 139880 93634 139922
rect 93342 139840 93344 139880
rect 93344 139840 93386 139880
rect 93386 139840 93426 139880
rect 93426 139840 93466 139880
rect 93510 139840 93550 139880
rect 93550 139840 93590 139880
rect 93590 139840 93632 139880
rect 93632 139840 93634 139880
rect 93342 139798 93466 139840
rect 93510 139798 93634 139840
rect 108462 139880 108586 139922
rect 108630 139880 108754 139922
rect 108462 139840 108464 139880
rect 108464 139840 108506 139880
rect 108506 139840 108546 139880
rect 108546 139840 108586 139880
rect 108630 139840 108670 139880
rect 108670 139840 108710 139880
rect 108710 139840 108752 139880
rect 108752 139840 108754 139880
rect 108462 139798 108586 139840
rect 108630 139798 108754 139840
rect 123582 139880 123706 139922
rect 123750 139880 123874 139922
rect 123582 139840 123584 139880
rect 123584 139840 123626 139880
rect 123626 139840 123666 139880
rect 123666 139840 123706 139880
rect 123750 139840 123790 139880
rect 123790 139840 123830 139880
rect 123830 139840 123872 139880
rect 123872 139840 123874 139880
rect 123582 139798 123706 139840
rect 123750 139798 123874 139840
rect 138702 139880 138826 139922
rect 138870 139880 138994 139922
rect 138702 139840 138704 139880
rect 138704 139840 138746 139880
rect 138746 139840 138786 139880
rect 138786 139840 138826 139880
rect 138870 139840 138910 139880
rect 138910 139840 138950 139880
rect 138950 139840 138992 139880
rect 138992 139840 138994 139880
rect 138702 139798 138826 139840
rect 138870 139798 138994 139840
rect 79462 139124 79586 139166
rect 79630 139124 79754 139166
rect 79462 139084 79464 139124
rect 79464 139084 79506 139124
rect 79506 139084 79546 139124
rect 79546 139084 79586 139124
rect 79630 139084 79670 139124
rect 79670 139084 79710 139124
rect 79710 139084 79752 139124
rect 79752 139084 79754 139124
rect 79462 139042 79586 139084
rect 79630 139042 79754 139084
rect 94582 139124 94706 139166
rect 94750 139124 94874 139166
rect 94582 139084 94584 139124
rect 94584 139084 94626 139124
rect 94626 139084 94666 139124
rect 94666 139084 94706 139124
rect 94750 139084 94790 139124
rect 94790 139084 94830 139124
rect 94830 139084 94872 139124
rect 94872 139084 94874 139124
rect 94582 139042 94706 139084
rect 94750 139042 94874 139084
rect 109702 139124 109826 139166
rect 109870 139124 109994 139166
rect 109702 139084 109704 139124
rect 109704 139084 109746 139124
rect 109746 139084 109786 139124
rect 109786 139084 109826 139124
rect 109870 139084 109910 139124
rect 109910 139084 109950 139124
rect 109950 139084 109992 139124
rect 109992 139084 109994 139124
rect 109702 139042 109826 139084
rect 109870 139042 109994 139084
rect 124822 139124 124946 139166
rect 124990 139124 125114 139166
rect 124822 139084 124824 139124
rect 124824 139084 124866 139124
rect 124866 139084 124906 139124
rect 124906 139084 124946 139124
rect 124990 139084 125030 139124
rect 125030 139084 125070 139124
rect 125070 139084 125112 139124
rect 125112 139084 125114 139124
rect 124822 139042 124946 139084
rect 124990 139042 125114 139084
rect 139942 139124 140066 139166
rect 140110 139124 140234 139166
rect 139942 139084 139944 139124
rect 139944 139084 139986 139124
rect 139986 139084 140026 139124
rect 140026 139084 140066 139124
rect 140110 139084 140150 139124
rect 140150 139084 140190 139124
rect 140190 139084 140232 139124
rect 140232 139084 140234 139124
rect 139942 139042 140066 139084
rect 140110 139042 140234 139084
rect 78222 138368 78346 138410
rect 78390 138368 78514 138410
rect 78222 138328 78224 138368
rect 78224 138328 78266 138368
rect 78266 138328 78306 138368
rect 78306 138328 78346 138368
rect 78390 138328 78430 138368
rect 78430 138328 78470 138368
rect 78470 138328 78512 138368
rect 78512 138328 78514 138368
rect 78222 138286 78346 138328
rect 78390 138286 78514 138328
rect 93342 138368 93466 138410
rect 93510 138368 93634 138410
rect 93342 138328 93344 138368
rect 93344 138328 93386 138368
rect 93386 138328 93426 138368
rect 93426 138328 93466 138368
rect 93510 138328 93550 138368
rect 93550 138328 93590 138368
rect 93590 138328 93632 138368
rect 93632 138328 93634 138368
rect 93342 138286 93466 138328
rect 93510 138286 93634 138328
rect 108462 138368 108586 138410
rect 108630 138368 108754 138410
rect 108462 138328 108464 138368
rect 108464 138328 108506 138368
rect 108506 138328 108546 138368
rect 108546 138328 108586 138368
rect 108630 138328 108670 138368
rect 108670 138328 108710 138368
rect 108710 138328 108752 138368
rect 108752 138328 108754 138368
rect 108462 138286 108586 138328
rect 108630 138286 108754 138328
rect 123582 138368 123706 138410
rect 123750 138368 123874 138410
rect 123582 138328 123584 138368
rect 123584 138328 123626 138368
rect 123626 138328 123666 138368
rect 123666 138328 123706 138368
rect 123750 138328 123790 138368
rect 123790 138328 123830 138368
rect 123830 138328 123872 138368
rect 123872 138328 123874 138368
rect 123582 138286 123706 138328
rect 123750 138286 123874 138328
rect 138702 138368 138826 138410
rect 138870 138368 138994 138410
rect 138702 138328 138704 138368
rect 138704 138328 138746 138368
rect 138746 138328 138786 138368
rect 138786 138328 138826 138368
rect 138870 138328 138910 138368
rect 138910 138328 138950 138368
rect 138950 138328 138992 138368
rect 138992 138328 138994 138368
rect 138702 138286 138826 138328
rect 138870 138286 138994 138328
rect 79462 137612 79586 137654
rect 79630 137612 79754 137654
rect 79462 137572 79464 137612
rect 79464 137572 79506 137612
rect 79506 137572 79546 137612
rect 79546 137572 79586 137612
rect 79630 137572 79670 137612
rect 79670 137572 79710 137612
rect 79710 137572 79752 137612
rect 79752 137572 79754 137612
rect 79462 137530 79586 137572
rect 79630 137530 79754 137572
rect 94582 137612 94706 137654
rect 94750 137612 94874 137654
rect 94582 137572 94584 137612
rect 94584 137572 94626 137612
rect 94626 137572 94666 137612
rect 94666 137572 94706 137612
rect 94750 137572 94790 137612
rect 94790 137572 94830 137612
rect 94830 137572 94872 137612
rect 94872 137572 94874 137612
rect 94582 137530 94706 137572
rect 94750 137530 94874 137572
rect 109702 137612 109826 137654
rect 109870 137612 109994 137654
rect 109702 137572 109704 137612
rect 109704 137572 109746 137612
rect 109746 137572 109786 137612
rect 109786 137572 109826 137612
rect 109870 137572 109910 137612
rect 109910 137572 109950 137612
rect 109950 137572 109992 137612
rect 109992 137572 109994 137612
rect 109702 137530 109826 137572
rect 109870 137530 109994 137572
rect 124822 137612 124946 137654
rect 124990 137612 125114 137654
rect 124822 137572 124824 137612
rect 124824 137572 124866 137612
rect 124866 137572 124906 137612
rect 124906 137572 124946 137612
rect 124990 137572 125030 137612
rect 125030 137572 125070 137612
rect 125070 137572 125112 137612
rect 125112 137572 125114 137612
rect 124822 137530 124946 137572
rect 124990 137530 125114 137572
rect 139942 137612 140066 137654
rect 140110 137612 140234 137654
rect 139942 137572 139944 137612
rect 139944 137572 139986 137612
rect 139986 137572 140026 137612
rect 140026 137572 140066 137612
rect 140110 137572 140150 137612
rect 140150 137572 140190 137612
rect 140190 137572 140232 137612
rect 140232 137572 140234 137612
rect 139942 137530 140066 137572
rect 140110 137530 140234 137572
rect 78222 136856 78346 136898
rect 78390 136856 78514 136898
rect 78222 136816 78224 136856
rect 78224 136816 78266 136856
rect 78266 136816 78306 136856
rect 78306 136816 78346 136856
rect 78390 136816 78430 136856
rect 78430 136816 78470 136856
rect 78470 136816 78512 136856
rect 78512 136816 78514 136856
rect 78222 136774 78346 136816
rect 78390 136774 78514 136816
rect 93342 136856 93466 136898
rect 93510 136856 93634 136898
rect 93342 136816 93344 136856
rect 93344 136816 93386 136856
rect 93386 136816 93426 136856
rect 93426 136816 93466 136856
rect 93510 136816 93550 136856
rect 93550 136816 93590 136856
rect 93590 136816 93632 136856
rect 93632 136816 93634 136856
rect 93342 136774 93466 136816
rect 93510 136774 93634 136816
rect 108462 136856 108586 136898
rect 108630 136856 108754 136898
rect 108462 136816 108464 136856
rect 108464 136816 108506 136856
rect 108506 136816 108546 136856
rect 108546 136816 108586 136856
rect 108630 136816 108670 136856
rect 108670 136816 108710 136856
rect 108710 136816 108752 136856
rect 108752 136816 108754 136856
rect 108462 136774 108586 136816
rect 108630 136774 108754 136816
rect 123582 136856 123706 136898
rect 123750 136856 123874 136898
rect 123582 136816 123584 136856
rect 123584 136816 123626 136856
rect 123626 136816 123666 136856
rect 123666 136816 123706 136856
rect 123750 136816 123790 136856
rect 123790 136816 123830 136856
rect 123830 136816 123872 136856
rect 123872 136816 123874 136856
rect 123582 136774 123706 136816
rect 123750 136774 123874 136816
rect 138702 136856 138826 136898
rect 138870 136856 138994 136898
rect 138702 136816 138704 136856
rect 138704 136816 138746 136856
rect 138746 136816 138786 136856
rect 138786 136816 138826 136856
rect 138870 136816 138910 136856
rect 138910 136816 138950 136856
rect 138950 136816 138992 136856
rect 138992 136816 138994 136856
rect 138702 136774 138826 136816
rect 138870 136774 138994 136816
rect 79462 136100 79586 136142
rect 79630 136100 79754 136142
rect 79462 136060 79464 136100
rect 79464 136060 79506 136100
rect 79506 136060 79546 136100
rect 79546 136060 79586 136100
rect 79630 136060 79670 136100
rect 79670 136060 79710 136100
rect 79710 136060 79752 136100
rect 79752 136060 79754 136100
rect 79462 136018 79586 136060
rect 79630 136018 79754 136060
rect 94582 136100 94706 136142
rect 94750 136100 94874 136142
rect 94582 136060 94584 136100
rect 94584 136060 94626 136100
rect 94626 136060 94666 136100
rect 94666 136060 94706 136100
rect 94750 136060 94790 136100
rect 94790 136060 94830 136100
rect 94830 136060 94872 136100
rect 94872 136060 94874 136100
rect 94582 136018 94706 136060
rect 94750 136018 94874 136060
rect 109702 136100 109826 136142
rect 109870 136100 109994 136142
rect 109702 136060 109704 136100
rect 109704 136060 109746 136100
rect 109746 136060 109786 136100
rect 109786 136060 109826 136100
rect 109870 136060 109910 136100
rect 109910 136060 109950 136100
rect 109950 136060 109992 136100
rect 109992 136060 109994 136100
rect 109702 136018 109826 136060
rect 109870 136018 109994 136060
rect 124822 136100 124946 136142
rect 124990 136100 125114 136142
rect 124822 136060 124824 136100
rect 124824 136060 124866 136100
rect 124866 136060 124906 136100
rect 124906 136060 124946 136100
rect 124990 136060 125030 136100
rect 125030 136060 125070 136100
rect 125070 136060 125112 136100
rect 125112 136060 125114 136100
rect 124822 136018 124946 136060
rect 124990 136018 125114 136060
rect 139942 136100 140066 136142
rect 140110 136100 140234 136142
rect 139942 136060 139944 136100
rect 139944 136060 139986 136100
rect 139986 136060 140026 136100
rect 140026 136060 140066 136100
rect 140110 136060 140150 136100
rect 140150 136060 140190 136100
rect 140190 136060 140232 136100
rect 140232 136060 140234 136100
rect 139942 136018 140066 136060
rect 140110 136018 140234 136060
rect 78222 135344 78346 135386
rect 78390 135344 78514 135386
rect 78222 135304 78224 135344
rect 78224 135304 78266 135344
rect 78266 135304 78306 135344
rect 78306 135304 78346 135344
rect 78390 135304 78430 135344
rect 78430 135304 78470 135344
rect 78470 135304 78512 135344
rect 78512 135304 78514 135344
rect 78222 135262 78346 135304
rect 78390 135262 78514 135304
rect 93342 135344 93466 135386
rect 93510 135344 93634 135386
rect 93342 135304 93344 135344
rect 93344 135304 93386 135344
rect 93386 135304 93426 135344
rect 93426 135304 93466 135344
rect 93510 135304 93550 135344
rect 93550 135304 93590 135344
rect 93590 135304 93632 135344
rect 93632 135304 93634 135344
rect 93342 135262 93466 135304
rect 93510 135262 93634 135304
rect 108462 135344 108586 135386
rect 108630 135344 108754 135386
rect 108462 135304 108464 135344
rect 108464 135304 108506 135344
rect 108506 135304 108546 135344
rect 108546 135304 108586 135344
rect 108630 135304 108670 135344
rect 108670 135304 108710 135344
rect 108710 135304 108752 135344
rect 108752 135304 108754 135344
rect 108462 135262 108586 135304
rect 108630 135262 108754 135304
rect 123582 135344 123706 135386
rect 123750 135344 123874 135386
rect 123582 135304 123584 135344
rect 123584 135304 123626 135344
rect 123626 135304 123666 135344
rect 123666 135304 123706 135344
rect 123750 135304 123790 135344
rect 123790 135304 123830 135344
rect 123830 135304 123872 135344
rect 123872 135304 123874 135344
rect 123582 135262 123706 135304
rect 123750 135262 123874 135304
rect 138702 135344 138826 135386
rect 138870 135344 138994 135386
rect 138702 135304 138704 135344
rect 138704 135304 138746 135344
rect 138746 135304 138786 135344
rect 138786 135304 138826 135344
rect 138870 135304 138910 135344
rect 138910 135304 138950 135344
rect 138950 135304 138992 135344
rect 138992 135304 138994 135344
rect 138702 135262 138826 135304
rect 138870 135262 138994 135304
rect 79462 134588 79586 134630
rect 79630 134588 79754 134630
rect 79462 134548 79464 134588
rect 79464 134548 79506 134588
rect 79506 134548 79546 134588
rect 79546 134548 79586 134588
rect 79630 134548 79670 134588
rect 79670 134548 79710 134588
rect 79710 134548 79752 134588
rect 79752 134548 79754 134588
rect 79462 134506 79586 134548
rect 79630 134506 79754 134548
rect 94582 134588 94706 134630
rect 94750 134588 94874 134630
rect 94582 134548 94584 134588
rect 94584 134548 94626 134588
rect 94626 134548 94666 134588
rect 94666 134548 94706 134588
rect 94750 134548 94790 134588
rect 94790 134548 94830 134588
rect 94830 134548 94872 134588
rect 94872 134548 94874 134588
rect 94582 134506 94706 134548
rect 94750 134506 94874 134548
rect 109702 134588 109826 134630
rect 109870 134588 109994 134630
rect 109702 134548 109704 134588
rect 109704 134548 109746 134588
rect 109746 134548 109786 134588
rect 109786 134548 109826 134588
rect 109870 134548 109910 134588
rect 109910 134548 109950 134588
rect 109950 134548 109992 134588
rect 109992 134548 109994 134588
rect 109702 134506 109826 134548
rect 109870 134506 109994 134548
rect 124822 134588 124946 134630
rect 124990 134588 125114 134630
rect 124822 134548 124824 134588
rect 124824 134548 124866 134588
rect 124866 134548 124906 134588
rect 124906 134548 124946 134588
rect 124990 134548 125030 134588
rect 125030 134548 125070 134588
rect 125070 134548 125112 134588
rect 125112 134548 125114 134588
rect 124822 134506 124946 134548
rect 124990 134506 125114 134548
rect 139942 134588 140066 134630
rect 140110 134588 140234 134630
rect 139942 134548 139944 134588
rect 139944 134548 139986 134588
rect 139986 134548 140026 134588
rect 140026 134548 140066 134588
rect 140110 134548 140150 134588
rect 140150 134548 140190 134588
rect 140190 134548 140232 134588
rect 140232 134548 140234 134588
rect 139942 134506 140066 134548
rect 140110 134506 140234 134548
rect 78222 133832 78346 133874
rect 78390 133832 78514 133874
rect 78222 133792 78224 133832
rect 78224 133792 78266 133832
rect 78266 133792 78306 133832
rect 78306 133792 78346 133832
rect 78390 133792 78430 133832
rect 78430 133792 78470 133832
rect 78470 133792 78512 133832
rect 78512 133792 78514 133832
rect 78222 133750 78346 133792
rect 78390 133750 78514 133792
rect 93342 133832 93466 133874
rect 93510 133832 93634 133874
rect 93342 133792 93344 133832
rect 93344 133792 93386 133832
rect 93386 133792 93426 133832
rect 93426 133792 93466 133832
rect 93510 133792 93550 133832
rect 93550 133792 93590 133832
rect 93590 133792 93632 133832
rect 93632 133792 93634 133832
rect 93342 133750 93466 133792
rect 93510 133750 93634 133792
rect 108462 133832 108586 133874
rect 108630 133832 108754 133874
rect 108462 133792 108464 133832
rect 108464 133792 108506 133832
rect 108506 133792 108546 133832
rect 108546 133792 108586 133832
rect 108630 133792 108670 133832
rect 108670 133792 108710 133832
rect 108710 133792 108752 133832
rect 108752 133792 108754 133832
rect 108462 133750 108586 133792
rect 108630 133750 108754 133792
rect 123582 133832 123706 133874
rect 123750 133832 123874 133874
rect 123582 133792 123584 133832
rect 123584 133792 123626 133832
rect 123626 133792 123666 133832
rect 123666 133792 123706 133832
rect 123750 133792 123790 133832
rect 123790 133792 123830 133832
rect 123830 133792 123872 133832
rect 123872 133792 123874 133832
rect 123582 133750 123706 133792
rect 123750 133750 123874 133792
rect 138702 133832 138826 133874
rect 138870 133832 138994 133874
rect 138702 133792 138704 133832
rect 138704 133792 138746 133832
rect 138746 133792 138786 133832
rect 138786 133792 138826 133832
rect 138870 133792 138910 133832
rect 138910 133792 138950 133832
rect 138950 133792 138992 133832
rect 138992 133792 138994 133832
rect 138702 133750 138826 133792
rect 138870 133750 138994 133792
rect 79462 133076 79586 133118
rect 79630 133076 79754 133118
rect 79462 133036 79464 133076
rect 79464 133036 79506 133076
rect 79506 133036 79546 133076
rect 79546 133036 79586 133076
rect 79630 133036 79670 133076
rect 79670 133036 79710 133076
rect 79710 133036 79752 133076
rect 79752 133036 79754 133076
rect 79462 132994 79586 133036
rect 79630 132994 79754 133036
rect 94582 133076 94706 133118
rect 94750 133076 94874 133118
rect 94582 133036 94584 133076
rect 94584 133036 94626 133076
rect 94626 133036 94666 133076
rect 94666 133036 94706 133076
rect 94750 133036 94790 133076
rect 94790 133036 94830 133076
rect 94830 133036 94872 133076
rect 94872 133036 94874 133076
rect 94582 132994 94706 133036
rect 94750 132994 94874 133036
rect 109702 133076 109826 133118
rect 109870 133076 109994 133118
rect 109702 133036 109704 133076
rect 109704 133036 109746 133076
rect 109746 133036 109786 133076
rect 109786 133036 109826 133076
rect 109870 133036 109910 133076
rect 109910 133036 109950 133076
rect 109950 133036 109992 133076
rect 109992 133036 109994 133076
rect 109702 132994 109826 133036
rect 109870 132994 109994 133036
rect 124822 133076 124946 133118
rect 124990 133076 125114 133118
rect 124822 133036 124824 133076
rect 124824 133036 124866 133076
rect 124866 133036 124906 133076
rect 124906 133036 124946 133076
rect 124990 133036 125030 133076
rect 125030 133036 125070 133076
rect 125070 133036 125112 133076
rect 125112 133036 125114 133076
rect 124822 132994 124946 133036
rect 124990 132994 125114 133036
rect 139942 133076 140066 133118
rect 140110 133076 140234 133118
rect 139942 133036 139944 133076
rect 139944 133036 139986 133076
rect 139986 133036 140026 133076
rect 140026 133036 140066 133076
rect 140110 133036 140150 133076
rect 140150 133036 140190 133076
rect 140190 133036 140232 133076
rect 140232 133036 140234 133076
rect 139942 132994 140066 133036
rect 140110 132994 140234 133036
rect 78222 132320 78346 132362
rect 78390 132320 78514 132362
rect 78222 132280 78224 132320
rect 78224 132280 78266 132320
rect 78266 132280 78306 132320
rect 78306 132280 78346 132320
rect 78390 132280 78430 132320
rect 78430 132280 78470 132320
rect 78470 132280 78512 132320
rect 78512 132280 78514 132320
rect 78222 132238 78346 132280
rect 78390 132238 78514 132280
rect 93342 132320 93466 132362
rect 93510 132320 93634 132362
rect 93342 132280 93344 132320
rect 93344 132280 93386 132320
rect 93386 132280 93426 132320
rect 93426 132280 93466 132320
rect 93510 132280 93550 132320
rect 93550 132280 93590 132320
rect 93590 132280 93632 132320
rect 93632 132280 93634 132320
rect 93342 132238 93466 132280
rect 93510 132238 93634 132280
rect 108462 132320 108586 132362
rect 108630 132320 108754 132362
rect 108462 132280 108464 132320
rect 108464 132280 108506 132320
rect 108506 132280 108546 132320
rect 108546 132280 108586 132320
rect 108630 132280 108670 132320
rect 108670 132280 108710 132320
rect 108710 132280 108752 132320
rect 108752 132280 108754 132320
rect 108462 132238 108586 132280
rect 108630 132238 108754 132280
rect 123582 132320 123706 132362
rect 123750 132320 123874 132362
rect 123582 132280 123584 132320
rect 123584 132280 123626 132320
rect 123626 132280 123666 132320
rect 123666 132280 123706 132320
rect 123750 132280 123790 132320
rect 123790 132280 123830 132320
rect 123830 132280 123872 132320
rect 123872 132280 123874 132320
rect 123582 132238 123706 132280
rect 123750 132238 123874 132280
rect 138702 132320 138826 132362
rect 138870 132320 138994 132362
rect 138702 132280 138704 132320
rect 138704 132280 138746 132320
rect 138746 132280 138786 132320
rect 138786 132280 138826 132320
rect 138870 132280 138910 132320
rect 138910 132280 138950 132320
rect 138950 132280 138992 132320
rect 138992 132280 138994 132320
rect 138702 132238 138826 132280
rect 138870 132238 138994 132280
rect 79462 131564 79586 131606
rect 79630 131564 79754 131606
rect 79462 131524 79464 131564
rect 79464 131524 79506 131564
rect 79506 131524 79546 131564
rect 79546 131524 79586 131564
rect 79630 131524 79670 131564
rect 79670 131524 79710 131564
rect 79710 131524 79752 131564
rect 79752 131524 79754 131564
rect 79462 131482 79586 131524
rect 79630 131482 79754 131524
rect 94582 131564 94706 131606
rect 94750 131564 94874 131606
rect 94582 131524 94584 131564
rect 94584 131524 94626 131564
rect 94626 131524 94666 131564
rect 94666 131524 94706 131564
rect 94750 131524 94790 131564
rect 94790 131524 94830 131564
rect 94830 131524 94872 131564
rect 94872 131524 94874 131564
rect 94582 131482 94706 131524
rect 94750 131482 94874 131524
rect 109702 131564 109826 131606
rect 109870 131564 109994 131606
rect 109702 131524 109704 131564
rect 109704 131524 109746 131564
rect 109746 131524 109786 131564
rect 109786 131524 109826 131564
rect 109870 131524 109910 131564
rect 109910 131524 109950 131564
rect 109950 131524 109992 131564
rect 109992 131524 109994 131564
rect 109702 131482 109826 131524
rect 109870 131482 109994 131524
rect 124822 131564 124946 131606
rect 124990 131564 125114 131606
rect 124822 131524 124824 131564
rect 124824 131524 124866 131564
rect 124866 131524 124906 131564
rect 124906 131524 124946 131564
rect 124990 131524 125030 131564
rect 125030 131524 125070 131564
rect 125070 131524 125112 131564
rect 125112 131524 125114 131564
rect 124822 131482 124946 131524
rect 124990 131482 125114 131524
rect 139942 131564 140066 131606
rect 140110 131564 140234 131606
rect 139942 131524 139944 131564
rect 139944 131524 139986 131564
rect 139986 131524 140026 131564
rect 140026 131524 140066 131564
rect 140110 131524 140150 131564
rect 140150 131524 140190 131564
rect 140190 131524 140232 131564
rect 140232 131524 140234 131564
rect 139942 131482 140066 131524
rect 140110 131482 140234 131524
rect 78222 130808 78346 130850
rect 78390 130808 78514 130850
rect 78222 130768 78224 130808
rect 78224 130768 78266 130808
rect 78266 130768 78306 130808
rect 78306 130768 78346 130808
rect 78390 130768 78430 130808
rect 78430 130768 78470 130808
rect 78470 130768 78512 130808
rect 78512 130768 78514 130808
rect 78222 130726 78346 130768
rect 78390 130726 78514 130768
rect 93342 130808 93466 130850
rect 93510 130808 93634 130850
rect 93342 130768 93344 130808
rect 93344 130768 93386 130808
rect 93386 130768 93426 130808
rect 93426 130768 93466 130808
rect 93510 130768 93550 130808
rect 93550 130768 93590 130808
rect 93590 130768 93632 130808
rect 93632 130768 93634 130808
rect 93342 130726 93466 130768
rect 93510 130726 93634 130768
rect 108462 130808 108586 130850
rect 108630 130808 108754 130850
rect 108462 130768 108464 130808
rect 108464 130768 108506 130808
rect 108506 130768 108546 130808
rect 108546 130768 108586 130808
rect 108630 130768 108670 130808
rect 108670 130768 108710 130808
rect 108710 130768 108752 130808
rect 108752 130768 108754 130808
rect 108462 130726 108586 130768
rect 108630 130726 108754 130768
rect 123582 130808 123706 130850
rect 123750 130808 123874 130850
rect 123582 130768 123584 130808
rect 123584 130768 123626 130808
rect 123626 130768 123666 130808
rect 123666 130768 123706 130808
rect 123750 130768 123790 130808
rect 123790 130768 123830 130808
rect 123830 130768 123872 130808
rect 123872 130768 123874 130808
rect 123582 130726 123706 130768
rect 123750 130726 123874 130768
rect 138702 130808 138826 130850
rect 138870 130808 138994 130850
rect 138702 130768 138704 130808
rect 138704 130768 138746 130808
rect 138746 130768 138786 130808
rect 138786 130768 138826 130808
rect 138870 130768 138910 130808
rect 138910 130768 138950 130808
rect 138950 130768 138992 130808
rect 138992 130768 138994 130808
rect 138702 130726 138826 130768
rect 138870 130726 138994 130768
rect 79462 130052 79586 130094
rect 79630 130052 79754 130094
rect 79462 130012 79464 130052
rect 79464 130012 79506 130052
rect 79506 130012 79546 130052
rect 79546 130012 79586 130052
rect 79630 130012 79670 130052
rect 79670 130012 79710 130052
rect 79710 130012 79752 130052
rect 79752 130012 79754 130052
rect 79462 129970 79586 130012
rect 79630 129970 79754 130012
rect 94582 130052 94706 130094
rect 94750 130052 94874 130094
rect 94582 130012 94584 130052
rect 94584 130012 94626 130052
rect 94626 130012 94666 130052
rect 94666 130012 94706 130052
rect 94750 130012 94790 130052
rect 94790 130012 94830 130052
rect 94830 130012 94872 130052
rect 94872 130012 94874 130052
rect 94582 129970 94706 130012
rect 94750 129970 94874 130012
rect 109702 130052 109826 130094
rect 109870 130052 109994 130094
rect 109702 130012 109704 130052
rect 109704 130012 109746 130052
rect 109746 130012 109786 130052
rect 109786 130012 109826 130052
rect 109870 130012 109910 130052
rect 109910 130012 109950 130052
rect 109950 130012 109992 130052
rect 109992 130012 109994 130052
rect 109702 129970 109826 130012
rect 109870 129970 109994 130012
rect 124822 130052 124946 130094
rect 124990 130052 125114 130094
rect 124822 130012 124824 130052
rect 124824 130012 124866 130052
rect 124866 130012 124906 130052
rect 124906 130012 124946 130052
rect 124990 130012 125030 130052
rect 125030 130012 125070 130052
rect 125070 130012 125112 130052
rect 125112 130012 125114 130052
rect 124822 129970 124946 130012
rect 124990 129970 125114 130012
rect 139942 130052 140066 130094
rect 140110 130052 140234 130094
rect 139942 130012 139944 130052
rect 139944 130012 139986 130052
rect 139986 130012 140026 130052
rect 140026 130012 140066 130052
rect 140110 130012 140150 130052
rect 140150 130012 140190 130052
rect 140190 130012 140232 130052
rect 140232 130012 140234 130052
rect 139942 129970 140066 130012
rect 140110 129970 140234 130012
rect 78222 129296 78346 129338
rect 78390 129296 78514 129338
rect 78222 129256 78224 129296
rect 78224 129256 78266 129296
rect 78266 129256 78306 129296
rect 78306 129256 78346 129296
rect 78390 129256 78430 129296
rect 78430 129256 78470 129296
rect 78470 129256 78512 129296
rect 78512 129256 78514 129296
rect 78222 129214 78346 129256
rect 78390 129214 78514 129256
rect 93342 129296 93466 129338
rect 93510 129296 93634 129338
rect 93342 129256 93344 129296
rect 93344 129256 93386 129296
rect 93386 129256 93426 129296
rect 93426 129256 93466 129296
rect 93510 129256 93550 129296
rect 93550 129256 93590 129296
rect 93590 129256 93632 129296
rect 93632 129256 93634 129296
rect 93342 129214 93466 129256
rect 93510 129214 93634 129256
rect 108462 129296 108586 129338
rect 108630 129296 108754 129338
rect 108462 129256 108464 129296
rect 108464 129256 108506 129296
rect 108506 129256 108546 129296
rect 108546 129256 108586 129296
rect 108630 129256 108670 129296
rect 108670 129256 108710 129296
rect 108710 129256 108752 129296
rect 108752 129256 108754 129296
rect 108462 129214 108586 129256
rect 108630 129214 108754 129256
rect 123582 129296 123706 129338
rect 123750 129296 123874 129338
rect 123582 129256 123584 129296
rect 123584 129256 123626 129296
rect 123626 129256 123666 129296
rect 123666 129256 123706 129296
rect 123750 129256 123790 129296
rect 123790 129256 123830 129296
rect 123830 129256 123872 129296
rect 123872 129256 123874 129296
rect 123582 129214 123706 129256
rect 123750 129214 123874 129256
rect 138702 129296 138826 129338
rect 138870 129296 138994 129338
rect 138702 129256 138704 129296
rect 138704 129256 138746 129296
rect 138746 129256 138786 129296
rect 138786 129256 138826 129296
rect 138870 129256 138910 129296
rect 138910 129256 138950 129296
rect 138950 129256 138992 129296
rect 138992 129256 138994 129296
rect 138702 129214 138826 129256
rect 138870 129214 138994 129256
rect 79462 128540 79586 128582
rect 79630 128540 79754 128582
rect 79462 128500 79464 128540
rect 79464 128500 79506 128540
rect 79506 128500 79546 128540
rect 79546 128500 79586 128540
rect 79630 128500 79670 128540
rect 79670 128500 79710 128540
rect 79710 128500 79752 128540
rect 79752 128500 79754 128540
rect 79462 128458 79586 128500
rect 79630 128458 79754 128500
rect 94582 128540 94706 128582
rect 94750 128540 94874 128582
rect 94582 128500 94584 128540
rect 94584 128500 94626 128540
rect 94626 128500 94666 128540
rect 94666 128500 94706 128540
rect 94750 128500 94790 128540
rect 94790 128500 94830 128540
rect 94830 128500 94872 128540
rect 94872 128500 94874 128540
rect 94582 128458 94706 128500
rect 94750 128458 94874 128500
rect 109702 128540 109826 128582
rect 109870 128540 109994 128582
rect 109702 128500 109704 128540
rect 109704 128500 109746 128540
rect 109746 128500 109786 128540
rect 109786 128500 109826 128540
rect 109870 128500 109910 128540
rect 109910 128500 109950 128540
rect 109950 128500 109992 128540
rect 109992 128500 109994 128540
rect 109702 128458 109826 128500
rect 109870 128458 109994 128500
rect 124822 128540 124946 128582
rect 124990 128540 125114 128582
rect 124822 128500 124824 128540
rect 124824 128500 124866 128540
rect 124866 128500 124906 128540
rect 124906 128500 124946 128540
rect 124990 128500 125030 128540
rect 125030 128500 125070 128540
rect 125070 128500 125112 128540
rect 125112 128500 125114 128540
rect 124822 128458 124946 128500
rect 124990 128458 125114 128500
rect 139942 128540 140066 128582
rect 140110 128540 140234 128582
rect 139942 128500 139944 128540
rect 139944 128500 139986 128540
rect 139986 128500 140026 128540
rect 140026 128500 140066 128540
rect 140110 128500 140150 128540
rect 140150 128500 140190 128540
rect 140190 128500 140232 128540
rect 140232 128500 140234 128540
rect 139942 128458 140066 128500
rect 140110 128458 140234 128500
rect 78222 127784 78346 127826
rect 78390 127784 78514 127826
rect 78222 127744 78224 127784
rect 78224 127744 78266 127784
rect 78266 127744 78306 127784
rect 78306 127744 78346 127784
rect 78390 127744 78430 127784
rect 78430 127744 78470 127784
rect 78470 127744 78512 127784
rect 78512 127744 78514 127784
rect 78222 127702 78346 127744
rect 78390 127702 78514 127744
rect 93342 127784 93466 127826
rect 93510 127784 93634 127826
rect 93342 127744 93344 127784
rect 93344 127744 93386 127784
rect 93386 127744 93426 127784
rect 93426 127744 93466 127784
rect 93510 127744 93550 127784
rect 93550 127744 93590 127784
rect 93590 127744 93632 127784
rect 93632 127744 93634 127784
rect 93342 127702 93466 127744
rect 93510 127702 93634 127744
rect 108462 127784 108586 127826
rect 108630 127784 108754 127826
rect 108462 127744 108464 127784
rect 108464 127744 108506 127784
rect 108506 127744 108546 127784
rect 108546 127744 108586 127784
rect 108630 127744 108670 127784
rect 108670 127744 108710 127784
rect 108710 127744 108752 127784
rect 108752 127744 108754 127784
rect 108462 127702 108586 127744
rect 108630 127702 108754 127744
rect 123582 127784 123706 127826
rect 123750 127784 123874 127826
rect 123582 127744 123584 127784
rect 123584 127744 123626 127784
rect 123626 127744 123666 127784
rect 123666 127744 123706 127784
rect 123750 127744 123790 127784
rect 123790 127744 123830 127784
rect 123830 127744 123872 127784
rect 123872 127744 123874 127784
rect 123582 127702 123706 127744
rect 123750 127702 123874 127744
rect 138702 127784 138826 127826
rect 138870 127784 138994 127826
rect 138702 127744 138704 127784
rect 138704 127744 138746 127784
rect 138746 127744 138786 127784
rect 138786 127744 138826 127784
rect 138870 127744 138910 127784
rect 138910 127744 138950 127784
rect 138950 127744 138992 127784
rect 138992 127744 138994 127784
rect 138702 127702 138826 127744
rect 138870 127702 138994 127744
rect 79462 127028 79586 127070
rect 79630 127028 79754 127070
rect 79462 126988 79464 127028
rect 79464 126988 79506 127028
rect 79506 126988 79546 127028
rect 79546 126988 79586 127028
rect 79630 126988 79670 127028
rect 79670 126988 79710 127028
rect 79710 126988 79752 127028
rect 79752 126988 79754 127028
rect 79462 126946 79586 126988
rect 79630 126946 79754 126988
rect 94582 127028 94706 127070
rect 94750 127028 94874 127070
rect 94582 126988 94584 127028
rect 94584 126988 94626 127028
rect 94626 126988 94666 127028
rect 94666 126988 94706 127028
rect 94750 126988 94790 127028
rect 94790 126988 94830 127028
rect 94830 126988 94872 127028
rect 94872 126988 94874 127028
rect 94582 126946 94706 126988
rect 94750 126946 94874 126988
rect 109702 127028 109826 127070
rect 109870 127028 109994 127070
rect 109702 126988 109704 127028
rect 109704 126988 109746 127028
rect 109746 126988 109786 127028
rect 109786 126988 109826 127028
rect 109870 126988 109910 127028
rect 109910 126988 109950 127028
rect 109950 126988 109992 127028
rect 109992 126988 109994 127028
rect 109702 126946 109826 126988
rect 109870 126946 109994 126988
rect 124822 127028 124946 127070
rect 124990 127028 125114 127070
rect 124822 126988 124824 127028
rect 124824 126988 124866 127028
rect 124866 126988 124906 127028
rect 124906 126988 124946 127028
rect 124990 126988 125030 127028
rect 125030 126988 125070 127028
rect 125070 126988 125112 127028
rect 125112 126988 125114 127028
rect 124822 126946 124946 126988
rect 124990 126946 125114 126988
rect 139942 127028 140066 127070
rect 140110 127028 140234 127070
rect 139942 126988 139944 127028
rect 139944 126988 139986 127028
rect 139986 126988 140026 127028
rect 140026 126988 140066 127028
rect 140110 126988 140150 127028
rect 140150 126988 140190 127028
rect 140190 126988 140232 127028
rect 140232 126988 140234 127028
rect 139942 126946 140066 126988
rect 140110 126946 140234 126988
rect 78222 126272 78346 126314
rect 78390 126272 78514 126314
rect 78222 126232 78224 126272
rect 78224 126232 78266 126272
rect 78266 126232 78306 126272
rect 78306 126232 78346 126272
rect 78390 126232 78430 126272
rect 78430 126232 78470 126272
rect 78470 126232 78512 126272
rect 78512 126232 78514 126272
rect 78222 126190 78346 126232
rect 78390 126190 78514 126232
rect 93342 126272 93466 126314
rect 93510 126272 93634 126314
rect 93342 126232 93344 126272
rect 93344 126232 93386 126272
rect 93386 126232 93426 126272
rect 93426 126232 93466 126272
rect 93510 126232 93550 126272
rect 93550 126232 93590 126272
rect 93590 126232 93632 126272
rect 93632 126232 93634 126272
rect 93342 126190 93466 126232
rect 93510 126190 93634 126232
rect 108462 126272 108586 126314
rect 108630 126272 108754 126314
rect 108462 126232 108464 126272
rect 108464 126232 108506 126272
rect 108506 126232 108546 126272
rect 108546 126232 108586 126272
rect 108630 126232 108670 126272
rect 108670 126232 108710 126272
rect 108710 126232 108752 126272
rect 108752 126232 108754 126272
rect 108462 126190 108586 126232
rect 108630 126190 108754 126232
rect 123582 126272 123706 126314
rect 123750 126272 123874 126314
rect 123582 126232 123584 126272
rect 123584 126232 123626 126272
rect 123626 126232 123666 126272
rect 123666 126232 123706 126272
rect 123750 126232 123790 126272
rect 123790 126232 123830 126272
rect 123830 126232 123872 126272
rect 123872 126232 123874 126272
rect 123582 126190 123706 126232
rect 123750 126190 123874 126232
rect 138702 126272 138826 126314
rect 138870 126272 138994 126314
rect 138702 126232 138704 126272
rect 138704 126232 138746 126272
rect 138746 126232 138786 126272
rect 138786 126232 138826 126272
rect 138870 126232 138910 126272
rect 138910 126232 138950 126272
rect 138950 126232 138992 126272
rect 138992 126232 138994 126272
rect 138702 126190 138826 126232
rect 138870 126190 138994 126232
rect 79462 125516 79586 125558
rect 79630 125516 79754 125558
rect 79462 125476 79464 125516
rect 79464 125476 79506 125516
rect 79506 125476 79546 125516
rect 79546 125476 79586 125516
rect 79630 125476 79670 125516
rect 79670 125476 79710 125516
rect 79710 125476 79752 125516
rect 79752 125476 79754 125516
rect 79462 125434 79586 125476
rect 79630 125434 79754 125476
rect 94582 125516 94706 125558
rect 94750 125516 94874 125558
rect 94582 125476 94584 125516
rect 94584 125476 94626 125516
rect 94626 125476 94666 125516
rect 94666 125476 94706 125516
rect 94750 125476 94790 125516
rect 94790 125476 94830 125516
rect 94830 125476 94872 125516
rect 94872 125476 94874 125516
rect 94582 125434 94706 125476
rect 94750 125434 94874 125476
rect 109702 125516 109826 125558
rect 109870 125516 109994 125558
rect 109702 125476 109704 125516
rect 109704 125476 109746 125516
rect 109746 125476 109786 125516
rect 109786 125476 109826 125516
rect 109870 125476 109910 125516
rect 109910 125476 109950 125516
rect 109950 125476 109992 125516
rect 109992 125476 109994 125516
rect 109702 125434 109826 125476
rect 109870 125434 109994 125476
rect 124822 125516 124946 125558
rect 124990 125516 125114 125558
rect 124822 125476 124824 125516
rect 124824 125476 124866 125516
rect 124866 125476 124906 125516
rect 124906 125476 124946 125516
rect 124990 125476 125030 125516
rect 125030 125476 125070 125516
rect 125070 125476 125112 125516
rect 125112 125476 125114 125516
rect 124822 125434 124946 125476
rect 124990 125434 125114 125476
rect 139942 125516 140066 125558
rect 140110 125516 140234 125558
rect 139942 125476 139944 125516
rect 139944 125476 139986 125516
rect 139986 125476 140026 125516
rect 140026 125476 140066 125516
rect 140110 125476 140150 125516
rect 140150 125476 140190 125516
rect 140190 125476 140232 125516
rect 140232 125476 140234 125516
rect 139942 125434 140066 125476
rect 140110 125434 140234 125476
rect 78222 124760 78346 124802
rect 78390 124760 78514 124802
rect 78222 124720 78224 124760
rect 78224 124720 78266 124760
rect 78266 124720 78306 124760
rect 78306 124720 78346 124760
rect 78390 124720 78430 124760
rect 78430 124720 78470 124760
rect 78470 124720 78512 124760
rect 78512 124720 78514 124760
rect 78222 124678 78346 124720
rect 78390 124678 78514 124720
rect 93342 124760 93466 124802
rect 93510 124760 93634 124802
rect 93342 124720 93344 124760
rect 93344 124720 93386 124760
rect 93386 124720 93426 124760
rect 93426 124720 93466 124760
rect 93510 124720 93550 124760
rect 93550 124720 93590 124760
rect 93590 124720 93632 124760
rect 93632 124720 93634 124760
rect 93342 124678 93466 124720
rect 93510 124678 93634 124720
rect 108462 124760 108586 124802
rect 108630 124760 108754 124802
rect 108462 124720 108464 124760
rect 108464 124720 108506 124760
rect 108506 124720 108546 124760
rect 108546 124720 108586 124760
rect 108630 124720 108670 124760
rect 108670 124720 108710 124760
rect 108710 124720 108752 124760
rect 108752 124720 108754 124760
rect 108462 124678 108586 124720
rect 108630 124678 108754 124720
rect 123582 124760 123706 124802
rect 123750 124760 123874 124802
rect 123582 124720 123584 124760
rect 123584 124720 123626 124760
rect 123626 124720 123666 124760
rect 123666 124720 123706 124760
rect 123750 124720 123790 124760
rect 123790 124720 123830 124760
rect 123830 124720 123872 124760
rect 123872 124720 123874 124760
rect 123582 124678 123706 124720
rect 123750 124678 123874 124720
rect 138702 124760 138826 124802
rect 138870 124760 138994 124802
rect 138702 124720 138704 124760
rect 138704 124720 138746 124760
rect 138746 124720 138786 124760
rect 138786 124720 138826 124760
rect 138870 124720 138910 124760
rect 138910 124720 138950 124760
rect 138950 124720 138992 124760
rect 138992 124720 138994 124760
rect 138702 124678 138826 124720
rect 138870 124678 138994 124720
rect 79462 124004 79586 124046
rect 79630 124004 79754 124046
rect 79462 123964 79464 124004
rect 79464 123964 79506 124004
rect 79506 123964 79546 124004
rect 79546 123964 79586 124004
rect 79630 123964 79670 124004
rect 79670 123964 79710 124004
rect 79710 123964 79752 124004
rect 79752 123964 79754 124004
rect 79462 123922 79586 123964
rect 79630 123922 79754 123964
rect 94582 124004 94706 124046
rect 94750 124004 94874 124046
rect 94582 123964 94584 124004
rect 94584 123964 94626 124004
rect 94626 123964 94666 124004
rect 94666 123964 94706 124004
rect 94750 123964 94790 124004
rect 94790 123964 94830 124004
rect 94830 123964 94872 124004
rect 94872 123964 94874 124004
rect 94582 123922 94706 123964
rect 94750 123922 94874 123964
rect 109702 124004 109826 124046
rect 109870 124004 109994 124046
rect 109702 123964 109704 124004
rect 109704 123964 109746 124004
rect 109746 123964 109786 124004
rect 109786 123964 109826 124004
rect 109870 123964 109910 124004
rect 109910 123964 109950 124004
rect 109950 123964 109992 124004
rect 109992 123964 109994 124004
rect 109702 123922 109826 123964
rect 109870 123922 109994 123964
rect 124822 124004 124946 124046
rect 124990 124004 125114 124046
rect 124822 123964 124824 124004
rect 124824 123964 124866 124004
rect 124866 123964 124906 124004
rect 124906 123964 124946 124004
rect 124990 123964 125030 124004
rect 125030 123964 125070 124004
rect 125070 123964 125112 124004
rect 125112 123964 125114 124004
rect 124822 123922 124946 123964
rect 124990 123922 125114 123964
rect 139942 124004 140066 124046
rect 140110 124004 140234 124046
rect 139942 123964 139944 124004
rect 139944 123964 139986 124004
rect 139986 123964 140026 124004
rect 140026 123964 140066 124004
rect 140110 123964 140150 124004
rect 140150 123964 140190 124004
rect 140190 123964 140232 124004
rect 140232 123964 140234 124004
rect 139942 123922 140066 123964
rect 140110 123922 140234 123964
rect 78222 123248 78346 123290
rect 78390 123248 78514 123290
rect 78222 123208 78224 123248
rect 78224 123208 78266 123248
rect 78266 123208 78306 123248
rect 78306 123208 78346 123248
rect 78390 123208 78430 123248
rect 78430 123208 78470 123248
rect 78470 123208 78512 123248
rect 78512 123208 78514 123248
rect 78222 123166 78346 123208
rect 78390 123166 78514 123208
rect 93342 123248 93466 123290
rect 93510 123248 93634 123290
rect 93342 123208 93344 123248
rect 93344 123208 93386 123248
rect 93386 123208 93426 123248
rect 93426 123208 93466 123248
rect 93510 123208 93550 123248
rect 93550 123208 93590 123248
rect 93590 123208 93632 123248
rect 93632 123208 93634 123248
rect 93342 123166 93466 123208
rect 93510 123166 93634 123208
rect 108462 123248 108586 123290
rect 108630 123248 108754 123290
rect 108462 123208 108464 123248
rect 108464 123208 108506 123248
rect 108506 123208 108546 123248
rect 108546 123208 108586 123248
rect 108630 123208 108670 123248
rect 108670 123208 108710 123248
rect 108710 123208 108752 123248
rect 108752 123208 108754 123248
rect 108462 123166 108586 123208
rect 108630 123166 108754 123208
rect 123582 123248 123706 123290
rect 123750 123248 123874 123290
rect 123582 123208 123584 123248
rect 123584 123208 123626 123248
rect 123626 123208 123666 123248
rect 123666 123208 123706 123248
rect 123750 123208 123790 123248
rect 123790 123208 123830 123248
rect 123830 123208 123872 123248
rect 123872 123208 123874 123248
rect 123582 123166 123706 123208
rect 123750 123166 123874 123208
rect 138702 123248 138826 123290
rect 138870 123248 138994 123290
rect 138702 123208 138704 123248
rect 138704 123208 138746 123248
rect 138746 123208 138786 123248
rect 138786 123208 138826 123248
rect 138870 123208 138910 123248
rect 138910 123208 138950 123248
rect 138950 123208 138992 123248
rect 138992 123208 138994 123248
rect 138702 123166 138826 123208
rect 138870 123166 138994 123208
rect 79462 122492 79586 122534
rect 79630 122492 79754 122534
rect 79462 122452 79464 122492
rect 79464 122452 79506 122492
rect 79506 122452 79546 122492
rect 79546 122452 79586 122492
rect 79630 122452 79670 122492
rect 79670 122452 79710 122492
rect 79710 122452 79752 122492
rect 79752 122452 79754 122492
rect 79462 122410 79586 122452
rect 79630 122410 79754 122452
rect 94582 122492 94706 122534
rect 94750 122492 94874 122534
rect 94582 122452 94584 122492
rect 94584 122452 94626 122492
rect 94626 122452 94666 122492
rect 94666 122452 94706 122492
rect 94750 122452 94790 122492
rect 94790 122452 94830 122492
rect 94830 122452 94872 122492
rect 94872 122452 94874 122492
rect 94582 122410 94706 122452
rect 94750 122410 94874 122452
rect 109702 122492 109826 122534
rect 109870 122492 109994 122534
rect 109702 122452 109704 122492
rect 109704 122452 109746 122492
rect 109746 122452 109786 122492
rect 109786 122452 109826 122492
rect 109870 122452 109910 122492
rect 109910 122452 109950 122492
rect 109950 122452 109992 122492
rect 109992 122452 109994 122492
rect 109702 122410 109826 122452
rect 109870 122410 109994 122452
rect 124822 122492 124946 122534
rect 124990 122492 125114 122534
rect 124822 122452 124824 122492
rect 124824 122452 124866 122492
rect 124866 122452 124906 122492
rect 124906 122452 124946 122492
rect 124990 122452 125030 122492
rect 125030 122452 125070 122492
rect 125070 122452 125112 122492
rect 125112 122452 125114 122492
rect 124822 122410 124946 122452
rect 124990 122410 125114 122452
rect 139942 122492 140066 122534
rect 140110 122492 140234 122534
rect 139942 122452 139944 122492
rect 139944 122452 139986 122492
rect 139986 122452 140026 122492
rect 140026 122452 140066 122492
rect 140110 122452 140150 122492
rect 140150 122452 140190 122492
rect 140190 122452 140232 122492
rect 140232 122452 140234 122492
rect 139942 122410 140066 122452
rect 140110 122410 140234 122452
rect 78222 121736 78346 121778
rect 78390 121736 78514 121778
rect 78222 121696 78224 121736
rect 78224 121696 78266 121736
rect 78266 121696 78306 121736
rect 78306 121696 78346 121736
rect 78390 121696 78430 121736
rect 78430 121696 78470 121736
rect 78470 121696 78512 121736
rect 78512 121696 78514 121736
rect 78222 121654 78346 121696
rect 78390 121654 78514 121696
rect 93342 121736 93466 121778
rect 93510 121736 93634 121778
rect 93342 121696 93344 121736
rect 93344 121696 93386 121736
rect 93386 121696 93426 121736
rect 93426 121696 93466 121736
rect 93510 121696 93550 121736
rect 93550 121696 93590 121736
rect 93590 121696 93632 121736
rect 93632 121696 93634 121736
rect 93342 121654 93466 121696
rect 93510 121654 93634 121696
rect 108462 121736 108586 121778
rect 108630 121736 108754 121778
rect 108462 121696 108464 121736
rect 108464 121696 108506 121736
rect 108506 121696 108546 121736
rect 108546 121696 108586 121736
rect 108630 121696 108670 121736
rect 108670 121696 108710 121736
rect 108710 121696 108752 121736
rect 108752 121696 108754 121736
rect 108462 121654 108586 121696
rect 108630 121654 108754 121696
rect 123582 121736 123706 121778
rect 123750 121736 123874 121778
rect 123582 121696 123584 121736
rect 123584 121696 123626 121736
rect 123626 121696 123666 121736
rect 123666 121696 123706 121736
rect 123750 121696 123790 121736
rect 123790 121696 123830 121736
rect 123830 121696 123872 121736
rect 123872 121696 123874 121736
rect 123582 121654 123706 121696
rect 123750 121654 123874 121696
rect 138702 121736 138826 121778
rect 138870 121736 138994 121778
rect 138702 121696 138704 121736
rect 138704 121696 138746 121736
rect 138746 121696 138786 121736
rect 138786 121696 138826 121736
rect 138870 121696 138910 121736
rect 138910 121696 138950 121736
rect 138950 121696 138992 121736
rect 138992 121696 138994 121736
rect 138702 121654 138826 121696
rect 138870 121654 138994 121696
rect 79462 120980 79586 121022
rect 79630 120980 79754 121022
rect 79462 120940 79464 120980
rect 79464 120940 79506 120980
rect 79506 120940 79546 120980
rect 79546 120940 79586 120980
rect 79630 120940 79670 120980
rect 79670 120940 79710 120980
rect 79710 120940 79752 120980
rect 79752 120940 79754 120980
rect 79462 120898 79586 120940
rect 79630 120898 79754 120940
rect 94582 120980 94706 121022
rect 94750 120980 94874 121022
rect 94582 120940 94584 120980
rect 94584 120940 94626 120980
rect 94626 120940 94666 120980
rect 94666 120940 94706 120980
rect 94750 120940 94790 120980
rect 94790 120940 94830 120980
rect 94830 120940 94872 120980
rect 94872 120940 94874 120980
rect 94582 120898 94706 120940
rect 94750 120898 94874 120940
rect 109702 120980 109826 121022
rect 109870 120980 109994 121022
rect 109702 120940 109704 120980
rect 109704 120940 109746 120980
rect 109746 120940 109786 120980
rect 109786 120940 109826 120980
rect 109870 120940 109910 120980
rect 109910 120940 109950 120980
rect 109950 120940 109992 120980
rect 109992 120940 109994 120980
rect 109702 120898 109826 120940
rect 109870 120898 109994 120940
rect 124822 120980 124946 121022
rect 124990 120980 125114 121022
rect 124822 120940 124824 120980
rect 124824 120940 124866 120980
rect 124866 120940 124906 120980
rect 124906 120940 124946 120980
rect 124990 120940 125030 120980
rect 125030 120940 125070 120980
rect 125070 120940 125112 120980
rect 125112 120940 125114 120980
rect 124822 120898 124946 120940
rect 124990 120898 125114 120940
rect 139942 120980 140066 121022
rect 140110 120980 140234 121022
rect 139942 120940 139944 120980
rect 139944 120940 139986 120980
rect 139986 120940 140026 120980
rect 140026 120940 140066 120980
rect 140110 120940 140150 120980
rect 140150 120940 140190 120980
rect 140190 120940 140232 120980
rect 140232 120940 140234 120980
rect 139942 120898 140066 120940
rect 140110 120898 140234 120940
rect 78222 120224 78346 120266
rect 78390 120224 78514 120266
rect 78222 120184 78224 120224
rect 78224 120184 78266 120224
rect 78266 120184 78306 120224
rect 78306 120184 78346 120224
rect 78390 120184 78430 120224
rect 78430 120184 78470 120224
rect 78470 120184 78512 120224
rect 78512 120184 78514 120224
rect 78222 120142 78346 120184
rect 78390 120142 78514 120184
rect 93342 120224 93466 120266
rect 93510 120224 93634 120266
rect 93342 120184 93344 120224
rect 93344 120184 93386 120224
rect 93386 120184 93426 120224
rect 93426 120184 93466 120224
rect 93510 120184 93550 120224
rect 93550 120184 93590 120224
rect 93590 120184 93632 120224
rect 93632 120184 93634 120224
rect 93342 120142 93466 120184
rect 93510 120142 93634 120184
rect 108462 120224 108586 120266
rect 108630 120224 108754 120266
rect 108462 120184 108464 120224
rect 108464 120184 108506 120224
rect 108506 120184 108546 120224
rect 108546 120184 108586 120224
rect 108630 120184 108670 120224
rect 108670 120184 108710 120224
rect 108710 120184 108752 120224
rect 108752 120184 108754 120224
rect 108462 120142 108586 120184
rect 108630 120142 108754 120184
rect 123582 120224 123706 120266
rect 123750 120224 123874 120266
rect 123582 120184 123584 120224
rect 123584 120184 123626 120224
rect 123626 120184 123666 120224
rect 123666 120184 123706 120224
rect 123750 120184 123790 120224
rect 123790 120184 123830 120224
rect 123830 120184 123872 120224
rect 123872 120184 123874 120224
rect 123582 120142 123706 120184
rect 123750 120142 123874 120184
rect 138702 120224 138826 120266
rect 138870 120224 138994 120266
rect 138702 120184 138704 120224
rect 138704 120184 138746 120224
rect 138746 120184 138786 120224
rect 138786 120184 138826 120224
rect 138870 120184 138910 120224
rect 138910 120184 138950 120224
rect 138950 120184 138992 120224
rect 138992 120184 138994 120224
rect 138702 120142 138826 120184
rect 138870 120142 138994 120184
rect 79462 119468 79586 119510
rect 79630 119468 79754 119510
rect 79462 119428 79464 119468
rect 79464 119428 79506 119468
rect 79506 119428 79546 119468
rect 79546 119428 79586 119468
rect 79630 119428 79670 119468
rect 79670 119428 79710 119468
rect 79710 119428 79752 119468
rect 79752 119428 79754 119468
rect 79462 119386 79586 119428
rect 79630 119386 79754 119428
rect 94582 119468 94706 119510
rect 94750 119468 94874 119510
rect 94582 119428 94584 119468
rect 94584 119428 94626 119468
rect 94626 119428 94666 119468
rect 94666 119428 94706 119468
rect 94750 119428 94790 119468
rect 94790 119428 94830 119468
rect 94830 119428 94872 119468
rect 94872 119428 94874 119468
rect 94582 119386 94706 119428
rect 94750 119386 94874 119428
rect 109702 119468 109826 119510
rect 109870 119468 109994 119510
rect 109702 119428 109704 119468
rect 109704 119428 109746 119468
rect 109746 119428 109786 119468
rect 109786 119428 109826 119468
rect 109870 119428 109910 119468
rect 109910 119428 109950 119468
rect 109950 119428 109992 119468
rect 109992 119428 109994 119468
rect 109702 119386 109826 119428
rect 109870 119386 109994 119428
rect 124822 119468 124946 119510
rect 124990 119468 125114 119510
rect 124822 119428 124824 119468
rect 124824 119428 124866 119468
rect 124866 119428 124906 119468
rect 124906 119428 124946 119468
rect 124990 119428 125030 119468
rect 125030 119428 125070 119468
rect 125070 119428 125112 119468
rect 125112 119428 125114 119468
rect 124822 119386 124946 119428
rect 124990 119386 125114 119428
rect 139942 119468 140066 119510
rect 140110 119468 140234 119510
rect 139942 119428 139944 119468
rect 139944 119428 139986 119468
rect 139986 119428 140026 119468
rect 140026 119428 140066 119468
rect 140110 119428 140150 119468
rect 140150 119428 140190 119468
rect 140190 119428 140232 119468
rect 140232 119428 140234 119468
rect 139942 119386 140066 119428
rect 140110 119386 140234 119428
rect 78222 118712 78346 118754
rect 78390 118712 78514 118754
rect 78222 118672 78224 118712
rect 78224 118672 78266 118712
rect 78266 118672 78306 118712
rect 78306 118672 78346 118712
rect 78390 118672 78430 118712
rect 78430 118672 78470 118712
rect 78470 118672 78512 118712
rect 78512 118672 78514 118712
rect 78222 118630 78346 118672
rect 78390 118630 78514 118672
rect 93342 118712 93466 118754
rect 93510 118712 93634 118754
rect 93342 118672 93344 118712
rect 93344 118672 93386 118712
rect 93386 118672 93426 118712
rect 93426 118672 93466 118712
rect 93510 118672 93550 118712
rect 93550 118672 93590 118712
rect 93590 118672 93632 118712
rect 93632 118672 93634 118712
rect 93342 118630 93466 118672
rect 93510 118630 93634 118672
rect 108462 118712 108586 118754
rect 108630 118712 108754 118754
rect 108462 118672 108464 118712
rect 108464 118672 108506 118712
rect 108506 118672 108546 118712
rect 108546 118672 108586 118712
rect 108630 118672 108670 118712
rect 108670 118672 108710 118712
rect 108710 118672 108752 118712
rect 108752 118672 108754 118712
rect 108462 118630 108586 118672
rect 108630 118630 108754 118672
rect 123582 118712 123706 118754
rect 123750 118712 123874 118754
rect 123582 118672 123584 118712
rect 123584 118672 123626 118712
rect 123626 118672 123666 118712
rect 123666 118672 123706 118712
rect 123750 118672 123790 118712
rect 123790 118672 123830 118712
rect 123830 118672 123872 118712
rect 123872 118672 123874 118712
rect 123582 118630 123706 118672
rect 123750 118630 123874 118672
rect 138702 118712 138826 118754
rect 138870 118712 138994 118754
rect 138702 118672 138704 118712
rect 138704 118672 138746 118712
rect 138746 118672 138786 118712
rect 138786 118672 138826 118712
rect 138870 118672 138910 118712
rect 138910 118672 138950 118712
rect 138950 118672 138992 118712
rect 138992 118672 138994 118712
rect 138702 118630 138826 118672
rect 138870 118630 138994 118672
rect 79462 117956 79586 117998
rect 79630 117956 79754 117998
rect 79462 117916 79464 117956
rect 79464 117916 79506 117956
rect 79506 117916 79546 117956
rect 79546 117916 79586 117956
rect 79630 117916 79670 117956
rect 79670 117916 79710 117956
rect 79710 117916 79752 117956
rect 79752 117916 79754 117956
rect 79462 117874 79586 117916
rect 79630 117874 79754 117916
rect 94582 117956 94706 117998
rect 94750 117956 94874 117998
rect 94582 117916 94584 117956
rect 94584 117916 94626 117956
rect 94626 117916 94666 117956
rect 94666 117916 94706 117956
rect 94750 117916 94790 117956
rect 94790 117916 94830 117956
rect 94830 117916 94872 117956
rect 94872 117916 94874 117956
rect 94582 117874 94706 117916
rect 94750 117874 94874 117916
rect 109702 117956 109826 117998
rect 109870 117956 109994 117998
rect 109702 117916 109704 117956
rect 109704 117916 109746 117956
rect 109746 117916 109786 117956
rect 109786 117916 109826 117956
rect 109870 117916 109910 117956
rect 109910 117916 109950 117956
rect 109950 117916 109992 117956
rect 109992 117916 109994 117956
rect 109702 117874 109826 117916
rect 109870 117874 109994 117916
rect 124822 117956 124946 117998
rect 124990 117956 125114 117998
rect 124822 117916 124824 117956
rect 124824 117916 124866 117956
rect 124866 117916 124906 117956
rect 124906 117916 124946 117956
rect 124990 117916 125030 117956
rect 125030 117916 125070 117956
rect 125070 117916 125112 117956
rect 125112 117916 125114 117956
rect 124822 117874 124946 117916
rect 124990 117874 125114 117916
rect 139942 117956 140066 117998
rect 140110 117956 140234 117998
rect 139942 117916 139944 117956
rect 139944 117916 139986 117956
rect 139986 117916 140026 117956
rect 140026 117916 140066 117956
rect 140110 117916 140150 117956
rect 140150 117916 140190 117956
rect 140190 117916 140232 117956
rect 140232 117916 140234 117956
rect 139942 117874 140066 117916
rect 140110 117874 140234 117916
rect 78222 117200 78346 117242
rect 78390 117200 78514 117242
rect 78222 117160 78224 117200
rect 78224 117160 78266 117200
rect 78266 117160 78306 117200
rect 78306 117160 78346 117200
rect 78390 117160 78430 117200
rect 78430 117160 78470 117200
rect 78470 117160 78512 117200
rect 78512 117160 78514 117200
rect 78222 117118 78346 117160
rect 78390 117118 78514 117160
rect 93342 117200 93466 117242
rect 93510 117200 93634 117242
rect 93342 117160 93344 117200
rect 93344 117160 93386 117200
rect 93386 117160 93426 117200
rect 93426 117160 93466 117200
rect 93510 117160 93550 117200
rect 93550 117160 93590 117200
rect 93590 117160 93632 117200
rect 93632 117160 93634 117200
rect 93342 117118 93466 117160
rect 93510 117118 93634 117160
rect 108462 117200 108586 117242
rect 108630 117200 108754 117242
rect 108462 117160 108464 117200
rect 108464 117160 108506 117200
rect 108506 117160 108546 117200
rect 108546 117160 108586 117200
rect 108630 117160 108670 117200
rect 108670 117160 108710 117200
rect 108710 117160 108752 117200
rect 108752 117160 108754 117200
rect 108462 117118 108586 117160
rect 108630 117118 108754 117160
rect 123582 117200 123706 117242
rect 123750 117200 123874 117242
rect 123582 117160 123584 117200
rect 123584 117160 123626 117200
rect 123626 117160 123666 117200
rect 123666 117160 123706 117200
rect 123750 117160 123790 117200
rect 123790 117160 123830 117200
rect 123830 117160 123872 117200
rect 123872 117160 123874 117200
rect 123582 117118 123706 117160
rect 123750 117118 123874 117160
rect 138702 117200 138826 117242
rect 138870 117200 138994 117242
rect 138702 117160 138704 117200
rect 138704 117160 138746 117200
rect 138746 117160 138786 117200
rect 138786 117160 138826 117200
rect 138870 117160 138910 117200
rect 138910 117160 138950 117200
rect 138950 117160 138992 117200
rect 138992 117160 138994 117200
rect 138702 117118 138826 117160
rect 138870 117118 138994 117160
rect 79462 116444 79586 116486
rect 79630 116444 79754 116486
rect 79462 116404 79464 116444
rect 79464 116404 79506 116444
rect 79506 116404 79546 116444
rect 79546 116404 79586 116444
rect 79630 116404 79670 116444
rect 79670 116404 79710 116444
rect 79710 116404 79752 116444
rect 79752 116404 79754 116444
rect 79462 116362 79586 116404
rect 79630 116362 79754 116404
rect 94582 116444 94706 116486
rect 94750 116444 94874 116486
rect 94582 116404 94584 116444
rect 94584 116404 94626 116444
rect 94626 116404 94666 116444
rect 94666 116404 94706 116444
rect 94750 116404 94790 116444
rect 94790 116404 94830 116444
rect 94830 116404 94872 116444
rect 94872 116404 94874 116444
rect 94582 116362 94706 116404
rect 94750 116362 94874 116404
rect 109702 116444 109826 116486
rect 109870 116444 109994 116486
rect 109702 116404 109704 116444
rect 109704 116404 109746 116444
rect 109746 116404 109786 116444
rect 109786 116404 109826 116444
rect 109870 116404 109910 116444
rect 109910 116404 109950 116444
rect 109950 116404 109992 116444
rect 109992 116404 109994 116444
rect 109702 116362 109826 116404
rect 109870 116362 109994 116404
rect 124822 116444 124946 116486
rect 124990 116444 125114 116486
rect 124822 116404 124824 116444
rect 124824 116404 124866 116444
rect 124866 116404 124906 116444
rect 124906 116404 124946 116444
rect 124990 116404 125030 116444
rect 125030 116404 125070 116444
rect 125070 116404 125112 116444
rect 125112 116404 125114 116444
rect 124822 116362 124946 116404
rect 124990 116362 125114 116404
rect 139942 116444 140066 116486
rect 140110 116444 140234 116486
rect 139942 116404 139944 116444
rect 139944 116404 139986 116444
rect 139986 116404 140026 116444
rect 140026 116404 140066 116444
rect 140110 116404 140150 116444
rect 140150 116404 140190 116444
rect 140190 116404 140232 116444
rect 140232 116404 140234 116444
rect 139942 116362 140066 116404
rect 140110 116362 140234 116404
rect 78222 115688 78346 115730
rect 78390 115688 78514 115730
rect 78222 115648 78224 115688
rect 78224 115648 78266 115688
rect 78266 115648 78306 115688
rect 78306 115648 78346 115688
rect 78390 115648 78430 115688
rect 78430 115648 78470 115688
rect 78470 115648 78512 115688
rect 78512 115648 78514 115688
rect 78222 115606 78346 115648
rect 78390 115606 78514 115648
rect 93342 115688 93466 115730
rect 93510 115688 93634 115730
rect 93342 115648 93344 115688
rect 93344 115648 93386 115688
rect 93386 115648 93426 115688
rect 93426 115648 93466 115688
rect 93510 115648 93550 115688
rect 93550 115648 93590 115688
rect 93590 115648 93632 115688
rect 93632 115648 93634 115688
rect 93342 115606 93466 115648
rect 93510 115606 93634 115648
rect 108462 115688 108586 115730
rect 108630 115688 108754 115730
rect 108462 115648 108464 115688
rect 108464 115648 108506 115688
rect 108506 115648 108546 115688
rect 108546 115648 108586 115688
rect 108630 115648 108670 115688
rect 108670 115648 108710 115688
rect 108710 115648 108752 115688
rect 108752 115648 108754 115688
rect 108462 115606 108586 115648
rect 108630 115606 108754 115648
rect 123582 115688 123706 115730
rect 123750 115688 123874 115730
rect 123582 115648 123584 115688
rect 123584 115648 123626 115688
rect 123626 115648 123666 115688
rect 123666 115648 123706 115688
rect 123750 115648 123790 115688
rect 123790 115648 123830 115688
rect 123830 115648 123872 115688
rect 123872 115648 123874 115688
rect 123582 115606 123706 115648
rect 123750 115606 123874 115648
rect 138702 115688 138826 115730
rect 138870 115688 138994 115730
rect 138702 115648 138704 115688
rect 138704 115648 138746 115688
rect 138746 115648 138786 115688
rect 138786 115648 138826 115688
rect 138870 115648 138910 115688
rect 138910 115648 138950 115688
rect 138950 115648 138992 115688
rect 138992 115648 138994 115688
rect 138702 115606 138826 115648
rect 138870 115606 138994 115648
rect 79462 114932 79586 114974
rect 79630 114932 79754 114974
rect 79462 114892 79464 114932
rect 79464 114892 79506 114932
rect 79506 114892 79546 114932
rect 79546 114892 79586 114932
rect 79630 114892 79670 114932
rect 79670 114892 79710 114932
rect 79710 114892 79752 114932
rect 79752 114892 79754 114932
rect 79462 114850 79586 114892
rect 79630 114850 79754 114892
rect 94582 114932 94706 114974
rect 94750 114932 94874 114974
rect 94582 114892 94584 114932
rect 94584 114892 94626 114932
rect 94626 114892 94666 114932
rect 94666 114892 94706 114932
rect 94750 114892 94790 114932
rect 94790 114892 94830 114932
rect 94830 114892 94872 114932
rect 94872 114892 94874 114932
rect 94582 114850 94706 114892
rect 94750 114850 94874 114892
rect 109702 114932 109826 114974
rect 109870 114932 109994 114974
rect 109702 114892 109704 114932
rect 109704 114892 109746 114932
rect 109746 114892 109786 114932
rect 109786 114892 109826 114932
rect 109870 114892 109910 114932
rect 109910 114892 109950 114932
rect 109950 114892 109992 114932
rect 109992 114892 109994 114932
rect 109702 114850 109826 114892
rect 109870 114850 109994 114892
rect 124822 114932 124946 114974
rect 124990 114932 125114 114974
rect 124822 114892 124824 114932
rect 124824 114892 124866 114932
rect 124866 114892 124906 114932
rect 124906 114892 124946 114932
rect 124990 114892 125030 114932
rect 125030 114892 125070 114932
rect 125070 114892 125112 114932
rect 125112 114892 125114 114932
rect 124822 114850 124946 114892
rect 124990 114850 125114 114892
rect 139942 114932 140066 114974
rect 140110 114932 140234 114974
rect 139942 114892 139944 114932
rect 139944 114892 139986 114932
rect 139986 114892 140026 114932
rect 140026 114892 140066 114932
rect 140110 114892 140150 114932
rect 140150 114892 140190 114932
rect 140190 114892 140232 114932
rect 140232 114892 140234 114932
rect 139942 114850 140066 114892
rect 140110 114850 140234 114892
rect 78222 114176 78346 114218
rect 78390 114176 78514 114218
rect 78222 114136 78224 114176
rect 78224 114136 78266 114176
rect 78266 114136 78306 114176
rect 78306 114136 78346 114176
rect 78390 114136 78430 114176
rect 78430 114136 78470 114176
rect 78470 114136 78512 114176
rect 78512 114136 78514 114176
rect 78222 114094 78346 114136
rect 78390 114094 78514 114136
rect 93342 114176 93466 114218
rect 93510 114176 93634 114218
rect 93342 114136 93344 114176
rect 93344 114136 93386 114176
rect 93386 114136 93426 114176
rect 93426 114136 93466 114176
rect 93510 114136 93550 114176
rect 93550 114136 93590 114176
rect 93590 114136 93632 114176
rect 93632 114136 93634 114176
rect 93342 114094 93466 114136
rect 93510 114094 93634 114136
rect 108462 114176 108586 114218
rect 108630 114176 108754 114218
rect 108462 114136 108464 114176
rect 108464 114136 108506 114176
rect 108506 114136 108546 114176
rect 108546 114136 108586 114176
rect 108630 114136 108670 114176
rect 108670 114136 108710 114176
rect 108710 114136 108752 114176
rect 108752 114136 108754 114176
rect 108462 114094 108586 114136
rect 108630 114094 108754 114136
rect 123582 114176 123706 114218
rect 123750 114176 123874 114218
rect 123582 114136 123584 114176
rect 123584 114136 123626 114176
rect 123626 114136 123666 114176
rect 123666 114136 123706 114176
rect 123750 114136 123790 114176
rect 123790 114136 123830 114176
rect 123830 114136 123872 114176
rect 123872 114136 123874 114176
rect 123582 114094 123706 114136
rect 123750 114094 123874 114136
rect 138702 114176 138826 114218
rect 138870 114176 138994 114218
rect 138702 114136 138704 114176
rect 138704 114136 138746 114176
rect 138746 114136 138786 114176
rect 138786 114136 138826 114176
rect 138870 114136 138910 114176
rect 138910 114136 138950 114176
rect 138950 114136 138992 114176
rect 138992 114136 138994 114176
rect 138702 114094 138826 114136
rect 138870 114094 138994 114136
rect 79462 113420 79586 113462
rect 79630 113420 79754 113462
rect 79462 113380 79464 113420
rect 79464 113380 79506 113420
rect 79506 113380 79546 113420
rect 79546 113380 79586 113420
rect 79630 113380 79670 113420
rect 79670 113380 79710 113420
rect 79710 113380 79752 113420
rect 79752 113380 79754 113420
rect 79462 113338 79586 113380
rect 79630 113338 79754 113380
rect 94582 113420 94706 113462
rect 94750 113420 94874 113462
rect 94582 113380 94584 113420
rect 94584 113380 94626 113420
rect 94626 113380 94666 113420
rect 94666 113380 94706 113420
rect 94750 113380 94790 113420
rect 94790 113380 94830 113420
rect 94830 113380 94872 113420
rect 94872 113380 94874 113420
rect 94582 113338 94706 113380
rect 94750 113338 94874 113380
rect 109702 113420 109826 113462
rect 109870 113420 109994 113462
rect 109702 113380 109704 113420
rect 109704 113380 109746 113420
rect 109746 113380 109786 113420
rect 109786 113380 109826 113420
rect 109870 113380 109910 113420
rect 109910 113380 109950 113420
rect 109950 113380 109992 113420
rect 109992 113380 109994 113420
rect 109702 113338 109826 113380
rect 109870 113338 109994 113380
rect 124822 113420 124946 113462
rect 124990 113420 125114 113462
rect 124822 113380 124824 113420
rect 124824 113380 124866 113420
rect 124866 113380 124906 113420
rect 124906 113380 124946 113420
rect 124990 113380 125030 113420
rect 125030 113380 125070 113420
rect 125070 113380 125112 113420
rect 125112 113380 125114 113420
rect 124822 113338 124946 113380
rect 124990 113338 125114 113380
rect 139942 113420 140066 113462
rect 140110 113420 140234 113462
rect 139942 113380 139944 113420
rect 139944 113380 139986 113420
rect 139986 113380 140026 113420
rect 140026 113380 140066 113420
rect 140110 113380 140150 113420
rect 140150 113380 140190 113420
rect 140190 113380 140232 113420
rect 140232 113380 140234 113420
rect 139942 113338 140066 113380
rect 140110 113338 140234 113380
rect 78222 112664 78346 112706
rect 78390 112664 78514 112706
rect 78222 112624 78224 112664
rect 78224 112624 78266 112664
rect 78266 112624 78306 112664
rect 78306 112624 78346 112664
rect 78390 112624 78430 112664
rect 78430 112624 78470 112664
rect 78470 112624 78512 112664
rect 78512 112624 78514 112664
rect 78222 112582 78346 112624
rect 78390 112582 78514 112624
rect 93342 112664 93466 112706
rect 93510 112664 93634 112706
rect 93342 112624 93344 112664
rect 93344 112624 93386 112664
rect 93386 112624 93426 112664
rect 93426 112624 93466 112664
rect 93510 112624 93550 112664
rect 93550 112624 93590 112664
rect 93590 112624 93632 112664
rect 93632 112624 93634 112664
rect 93342 112582 93466 112624
rect 93510 112582 93634 112624
rect 108462 112664 108586 112706
rect 108630 112664 108754 112706
rect 108462 112624 108464 112664
rect 108464 112624 108506 112664
rect 108506 112624 108546 112664
rect 108546 112624 108586 112664
rect 108630 112624 108670 112664
rect 108670 112624 108710 112664
rect 108710 112624 108752 112664
rect 108752 112624 108754 112664
rect 108462 112582 108586 112624
rect 108630 112582 108754 112624
rect 123582 112664 123706 112706
rect 123750 112664 123874 112706
rect 123582 112624 123584 112664
rect 123584 112624 123626 112664
rect 123626 112624 123666 112664
rect 123666 112624 123706 112664
rect 123750 112624 123790 112664
rect 123790 112624 123830 112664
rect 123830 112624 123872 112664
rect 123872 112624 123874 112664
rect 123582 112582 123706 112624
rect 123750 112582 123874 112624
rect 138702 112664 138826 112706
rect 138870 112664 138994 112706
rect 138702 112624 138704 112664
rect 138704 112624 138746 112664
rect 138746 112624 138786 112664
rect 138786 112624 138826 112664
rect 138870 112624 138910 112664
rect 138910 112624 138950 112664
rect 138950 112624 138992 112664
rect 138992 112624 138994 112664
rect 138702 112582 138826 112624
rect 138870 112582 138994 112624
rect 79462 111908 79586 111950
rect 79630 111908 79754 111950
rect 79462 111868 79464 111908
rect 79464 111868 79506 111908
rect 79506 111868 79546 111908
rect 79546 111868 79586 111908
rect 79630 111868 79670 111908
rect 79670 111868 79710 111908
rect 79710 111868 79752 111908
rect 79752 111868 79754 111908
rect 79462 111826 79586 111868
rect 79630 111826 79754 111868
rect 94582 111908 94706 111950
rect 94750 111908 94874 111950
rect 94582 111868 94584 111908
rect 94584 111868 94626 111908
rect 94626 111868 94666 111908
rect 94666 111868 94706 111908
rect 94750 111868 94790 111908
rect 94790 111868 94830 111908
rect 94830 111868 94872 111908
rect 94872 111868 94874 111908
rect 94582 111826 94706 111868
rect 94750 111826 94874 111868
rect 109702 111908 109826 111950
rect 109870 111908 109994 111950
rect 109702 111868 109704 111908
rect 109704 111868 109746 111908
rect 109746 111868 109786 111908
rect 109786 111868 109826 111908
rect 109870 111868 109910 111908
rect 109910 111868 109950 111908
rect 109950 111868 109992 111908
rect 109992 111868 109994 111908
rect 109702 111826 109826 111868
rect 109870 111826 109994 111868
rect 124822 111908 124946 111950
rect 124990 111908 125114 111950
rect 124822 111868 124824 111908
rect 124824 111868 124866 111908
rect 124866 111868 124906 111908
rect 124906 111868 124946 111908
rect 124990 111868 125030 111908
rect 125030 111868 125070 111908
rect 125070 111868 125112 111908
rect 125112 111868 125114 111908
rect 124822 111826 124946 111868
rect 124990 111826 125114 111868
rect 139942 111908 140066 111950
rect 140110 111908 140234 111950
rect 139942 111868 139944 111908
rect 139944 111868 139986 111908
rect 139986 111868 140026 111908
rect 140026 111868 140066 111908
rect 140110 111868 140150 111908
rect 140150 111868 140190 111908
rect 140190 111868 140232 111908
rect 140232 111868 140234 111908
rect 139942 111826 140066 111868
rect 140110 111826 140234 111868
rect 78222 111152 78346 111194
rect 78390 111152 78514 111194
rect 78222 111112 78224 111152
rect 78224 111112 78266 111152
rect 78266 111112 78306 111152
rect 78306 111112 78346 111152
rect 78390 111112 78430 111152
rect 78430 111112 78470 111152
rect 78470 111112 78512 111152
rect 78512 111112 78514 111152
rect 78222 111070 78346 111112
rect 78390 111070 78514 111112
rect 93342 111152 93466 111194
rect 93510 111152 93634 111194
rect 93342 111112 93344 111152
rect 93344 111112 93386 111152
rect 93386 111112 93426 111152
rect 93426 111112 93466 111152
rect 93510 111112 93550 111152
rect 93550 111112 93590 111152
rect 93590 111112 93632 111152
rect 93632 111112 93634 111152
rect 93342 111070 93466 111112
rect 93510 111070 93634 111112
rect 108462 111152 108586 111194
rect 108630 111152 108754 111194
rect 108462 111112 108464 111152
rect 108464 111112 108506 111152
rect 108506 111112 108546 111152
rect 108546 111112 108586 111152
rect 108630 111112 108670 111152
rect 108670 111112 108710 111152
rect 108710 111112 108752 111152
rect 108752 111112 108754 111152
rect 108462 111070 108586 111112
rect 108630 111070 108754 111112
rect 123582 111152 123706 111194
rect 123750 111152 123874 111194
rect 123582 111112 123584 111152
rect 123584 111112 123626 111152
rect 123626 111112 123666 111152
rect 123666 111112 123706 111152
rect 123750 111112 123790 111152
rect 123790 111112 123830 111152
rect 123830 111112 123872 111152
rect 123872 111112 123874 111152
rect 123582 111070 123706 111112
rect 123750 111070 123874 111112
rect 138702 111152 138826 111194
rect 138870 111152 138994 111194
rect 138702 111112 138704 111152
rect 138704 111112 138746 111152
rect 138746 111112 138786 111152
rect 138786 111112 138826 111152
rect 138870 111112 138910 111152
rect 138910 111112 138950 111152
rect 138950 111112 138992 111152
rect 138992 111112 138994 111152
rect 138702 111070 138826 111112
rect 138870 111070 138994 111112
rect 79462 110396 79586 110438
rect 79630 110396 79754 110438
rect 79462 110356 79464 110396
rect 79464 110356 79506 110396
rect 79506 110356 79546 110396
rect 79546 110356 79586 110396
rect 79630 110356 79670 110396
rect 79670 110356 79710 110396
rect 79710 110356 79752 110396
rect 79752 110356 79754 110396
rect 79462 110314 79586 110356
rect 79630 110314 79754 110356
rect 94582 110396 94706 110438
rect 94750 110396 94874 110438
rect 94582 110356 94584 110396
rect 94584 110356 94626 110396
rect 94626 110356 94666 110396
rect 94666 110356 94706 110396
rect 94750 110356 94790 110396
rect 94790 110356 94830 110396
rect 94830 110356 94872 110396
rect 94872 110356 94874 110396
rect 94582 110314 94706 110356
rect 94750 110314 94874 110356
rect 109702 110396 109826 110438
rect 109870 110396 109994 110438
rect 109702 110356 109704 110396
rect 109704 110356 109746 110396
rect 109746 110356 109786 110396
rect 109786 110356 109826 110396
rect 109870 110356 109910 110396
rect 109910 110356 109950 110396
rect 109950 110356 109992 110396
rect 109992 110356 109994 110396
rect 109702 110314 109826 110356
rect 109870 110314 109994 110356
rect 124822 110396 124946 110438
rect 124990 110396 125114 110438
rect 124822 110356 124824 110396
rect 124824 110356 124866 110396
rect 124866 110356 124906 110396
rect 124906 110356 124946 110396
rect 124990 110356 125030 110396
rect 125030 110356 125070 110396
rect 125070 110356 125112 110396
rect 125112 110356 125114 110396
rect 124822 110314 124946 110356
rect 124990 110314 125114 110356
rect 139942 110396 140066 110438
rect 140110 110396 140234 110438
rect 139942 110356 139944 110396
rect 139944 110356 139986 110396
rect 139986 110356 140026 110396
rect 140026 110356 140066 110396
rect 140110 110356 140150 110396
rect 140150 110356 140190 110396
rect 140190 110356 140232 110396
rect 140232 110356 140234 110396
rect 139942 110314 140066 110356
rect 140110 110314 140234 110356
rect 78222 109640 78346 109682
rect 78390 109640 78514 109682
rect 78222 109600 78224 109640
rect 78224 109600 78266 109640
rect 78266 109600 78306 109640
rect 78306 109600 78346 109640
rect 78390 109600 78430 109640
rect 78430 109600 78470 109640
rect 78470 109600 78512 109640
rect 78512 109600 78514 109640
rect 78222 109558 78346 109600
rect 78390 109558 78514 109600
rect 93342 109640 93466 109682
rect 93510 109640 93634 109682
rect 93342 109600 93344 109640
rect 93344 109600 93386 109640
rect 93386 109600 93426 109640
rect 93426 109600 93466 109640
rect 93510 109600 93550 109640
rect 93550 109600 93590 109640
rect 93590 109600 93632 109640
rect 93632 109600 93634 109640
rect 93342 109558 93466 109600
rect 93510 109558 93634 109600
rect 108462 109640 108586 109682
rect 108630 109640 108754 109682
rect 108462 109600 108464 109640
rect 108464 109600 108506 109640
rect 108506 109600 108546 109640
rect 108546 109600 108586 109640
rect 108630 109600 108670 109640
rect 108670 109600 108710 109640
rect 108710 109600 108752 109640
rect 108752 109600 108754 109640
rect 108462 109558 108586 109600
rect 108630 109558 108754 109600
rect 123582 109640 123706 109682
rect 123750 109640 123874 109682
rect 123582 109600 123584 109640
rect 123584 109600 123626 109640
rect 123626 109600 123666 109640
rect 123666 109600 123706 109640
rect 123750 109600 123790 109640
rect 123790 109600 123830 109640
rect 123830 109600 123872 109640
rect 123872 109600 123874 109640
rect 123582 109558 123706 109600
rect 123750 109558 123874 109600
rect 138702 109640 138826 109682
rect 138870 109640 138994 109682
rect 138702 109600 138704 109640
rect 138704 109600 138746 109640
rect 138746 109600 138786 109640
rect 138786 109600 138826 109640
rect 138870 109600 138910 109640
rect 138910 109600 138950 109640
rect 138950 109600 138992 109640
rect 138992 109600 138994 109640
rect 138702 109558 138826 109600
rect 138870 109558 138994 109600
rect 79462 108884 79586 108926
rect 79630 108884 79754 108926
rect 79462 108844 79464 108884
rect 79464 108844 79506 108884
rect 79506 108844 79546 108884
rect 79546 108844 79586 108884
rect 79630 108844 79670 108884
rect 79670 108844 79710 108884
rect 79710 108844 79752 108884
rect 79752 108844 79754 108884
rect 79462 108802 79586 108844
rect 79630 108802 79754 108844
rect 94582 108884 94706 108926
rect 94750 108884 94874 108926
rect 94582 108844 94584 108884
rect 94584 108844 94626 108884
rect 94626 108844 94666 108884
rect 94666 108844 94706 108884
rect 94750 108844 94790 108884
rect 94790 108844 94830 108884
rect 94830 108844 94872 108884
rect 94872 108844 94874 108884
rect 94582 108802 94706 108844
rect 94750 108802 94874 108844
rect 109702 108884 109826 108926
rect 109870 108884 109994 108926
rect 109702 108844 109704 108884
rect 109704 108844 109746 108884
rect 109746 108844 109786 108884
rect 109786 108844 109826 108884
rect 109870 108844 109910 108884
rect 109910 108844 109950 108884
rect 109950 108844 109992 108884
rect 109992 108844 109994 108884
rect 109702 108802 109826 108844
rect 109870 108802 109994 108844
rect 124822 108884 124946 108926
rect 124990 108884 125114 108926
rect 124822 108844 124824 108884
rect 124824 108844 124866 108884
rect 124866 108844 124906 108884
rect 124906 108844 124946 108884
rect 124990 108844 125030 108884
rect 125030 108844 125070 108884
rect 125070 108844 125112 108884
rect 125112 108844 125114 108884
rect 124822 108802 124946 108844
rect 124990 108802 125114 108844
rect 139942 108884 140066 108926
rect 140110 108884 140234 108926
rect 139942 108844 139944 108884
rect 139944 108844 139986 108884
rect 139986 108844 140026 108884
rect 140026 108844 140066 108884
rect 140110 108844 140150 108884
rect 140150 108844 140190 108884
rect 140190 108844 140232 108884
rect 140232 108844 140234 108884
rect 139942 108802 140066 108844
rect 140110 108802 140234 108844
rect 78222 108128 78346 108170
rect 78390 108128 78514 108170
rect 78222 108088 78224 108128
rect 78224 108088 78266 108128
rect 78266 108088 78306 108128
rect 78306 108088 78346 108128
rect 78390 108088 78430 108128
rect 78430 108088 78470 108128
rect 78470 108088 78512 108128
rect 78512 108088 78514 108128
rect 78222 108046 78346 108088
rect 78390 108046 78514 108088
rect 93342 108128 93466 108170
rect 93510 108128 93634 108170
rect 93342 108088 93344 108128
rect 93344 108088 93386 108128
rect 93386 108088 93426 108128
rect 93426 108088 93466 108128
rect 93510 108088 93550 108128
rect 93550 108088 93590 108128
rect 93590 108088 93632 108128
rect 93632 108088 93634 108128
rect 93342 108046 93466 108088
rect 93510 108046 93634 108088
rect 108462 108128 108586 108170
rect 108630 108128 108754 108170
rect 108462 108088 108464 108128
rect 108464 108088 108506 108128
rect 108506 108088 108546 108128
rect 108546 108088 108586 108128
rect 108630 108088 108670 108128
rect 108670 108088 108710 108128
rect 108710 108088 108752 108128
rect 108752 108088 108754 108128
rect 108462 108046 108586 108088
rect 108630 108046 108754 108088
rect 123582 108128 123706 108170
rect 123750 108128 123874 108170
rect 123582 108088 123584 108128
rect 123584 108088 123626 108128
rect 123626 108088 123666 108128
rect 123666 108088 123706 108128
rect 123750 108088 123790 108128
rect 123790 108088 123830 108128
rect 123830 108088 123872 108128
rect 123872 108088 123874 108128
rect 123582 108046 123706 108088
rect 123750 108046 123874 108088
rect 138702 108128 138826 108170
rect 138870 108128 138994 108170
rect 138702 108088 138704 108128
rect 138704 108088 138746 108128
rect 138746 108088 138786 108128
rect 138786 108088 138826 108128
rect 138870 108088 138910 108128
rect 138910 108088 138950 108128
rect 138950 108088 138992 108128
rect 138992 108088 138994 108128
rect 138702 108046 138826 108088
rect 138870 108046 138994 108088
rect 79462 107372 79586 107414
rect 79630 107372 79754 107414
rect 79462 107332 79464 107372
rect 79464 107332 79506 107372
rect 79506 107332 79546 107372
rect 79546 107332 79586 107372
rect 79630 107332 79670 107372
rect 79670 107332 79710 107372
rect 79710 107332 79752 107372
rect 79752 107332 79754 107372
rect 79462 107290 79586 107332
rect 79630 107290 79754 107332
rect 94582 107372 94706 107414
rect 94750 107372 94874 107414
rect 94582 107332 94584 107372
rect 94584 107332 94626 107372
rect 94626 107332 94666 107372
rect 94666 107332 94706 107372
rect 94750 107332 94790 107372
rect 94790 107332 94830 107372
rect 94830 107332 94872 107372
rect 94872 107332 94874 107372
rect 94582 107290 94706 107332
rect 94750 107290 94874 107332
rect 109702 107372 109826 107414
rect 109870 107372 109994 107414
rect 109702 107332 109704 107372
rect 109704 107332 109746 107372
rect 109746 107332 109786 107372
rect 109786 107332 109826 107372
rect 109870 107332 109910 107372
rect 109910 107332 109950 107372
rect 109950 107332 109992 107372
rect 109992 107332 109994 107372
rect 109702 107290 109826 107332
rect 109870 107290 109994 107332
rect 124822 107372 124946 107414
rect 124990 107372 125114 107414
rect 124822 107332 124824 107372
rect 124824 107332 124866 107372
rect 124866 107332 124906 107372
rect 124906 107332 124946 107372
rect 124990 107332 125030 107372
rect 125030 107332 125070 107372
rect 125070 107332 125112 107372
rect 125112 107332 125114 107372
rect 124822 107290 124946 107332
rect 124990 107290 125114 107332
rect 139942 107372 140066 107414
rect 140110 107372 140234 107414
rect 139942 107332 139944 107372
rect 139944 107332 139986 107372
rect 139986 107332 140026 107372
rect 140026 107332 140066 107372
rect 140110 107332 140150 107372
rect 140150 107332 140190 107372
rect 140190 107332 140232 107372
rect 140232 107332 140234 107372
rect 139942 107290 140066 107332
rect 140110 107290 140234 107332
rect 78222 106616 78346 106658
rect 78390 106616 78514 106658
rect 78222 106576 78224 106616
rect 78224 106576 78266 106616
rect 78266 106576 78306 106616
rect 78306 106576 78346 106616
rect 78390 106576 78430 106616
rect 78430 106576 78470 106616
rect 78470 106576 78512 106616
rect 78512 106576 78514 106616
rect 78222 106534 78346 106576
rect 78390 106534 78514 106576
rect 93342 106616 93466 106658
rect 93510 106616 93634 106658
rect 93342 106576 93344 106616
rect 93344 106576 93386 106616
rect 93386 106576 93426 106616
rect 93426 106576 93466 106616
rect 93510 106576 93550 106616
rect 93550 106576 93590 106616
rect 93590 106576 93632 106616
rect 93632 106576 93634 106616
rect 93342 106534 93466 106576
rect 93510 106534 93634 106576
rect 108462 106616 108586 106658
rect 108630 106616 108754 106658
rect 108462 106576 108464 106616
rect 108464 106576 108506 106616
rect 108506 106576 108546 106616
rect 108546 106576 108586 106616
rect 108630 106576 108670 106616
rect 108670 106576 108710 106616
rect 108710 106576 108752 106616
rect 108752 106576 108754 106616
rect 108462 106534 108586 106576
rect 108630 106534 108754 106576
rect 123582 106616 123706 106658
rect 123750 106616 123874 106658
rect 123582 106576 123584 106616
rect 123584 106576 123626 106616
rect 123626 106576 123666 106616
rect 123666 106576 123706 106616
rect 123750 106576 123790 106616
rect 123790 106576 123830 106616
rect 123830 106576 123872 106616
rect 123872 106576 123874 106616
rect 123582 106534 123706 106576
rect 123750 106534 123874 106576
rect 138702 106616 138826 106658
rect 138870 106616 138994 106658
rect 138702 106576 138704 106616
rect 138704 106576 138746 106616
rect 138746 106576 138786 106616
rect 138786 106576 138826 106616
rect 138870 106576 138910 106616
rect 138910 106576 138950 106616
rect 138950 106576 138992 106616
rect 138992 106576 138994 106616
rect 138702 106534 138826 106576
rect 138870 106534 138994 106576
rect 79462 105860 79586 105902
rect 79630 105860 79754 105902
rect 79462 105820 79464 105860
rect 79464 105820 79506 105860
rect 79506 105820 79546 105860
rect 79546 105820 79586 105860
rect 79630 105820 79670 105860
rect 79670 105820 79710 105860
rect 79710 105820 79752 105860
rect 79752 105820 79754 105860
rect 79462 105778 79586 105820
rect 79630 105778 79754 105820
rect 94582 105860 94706 105902
rect 94750 105860 94874 105902
rect 94582 105820 94584 105860
rect 94584 105820 94626 105860
rect 94626 105820 94666 105860
rect 94666 105820 94706 105860
rect 94750 105820 94790 105860
rect 94790 105820 94830 105860
rect 94830 105820 94872 105860
rect 94872 105820 94874 105860
rect 94582 105778 94706 105820
rect 94750 105778 94874 105820
rect 109702 105860 109826 105902
rect 109870 105860 109994 105902
rect 109702 105820 109704 105860
rect 109704 105820 109746 105860
rect 109746 105820 109786 105860
rect 109786 105820 109826 105860
rect 109870 105820 109910 105860
rect 109910 105820 109950 105860
rect 109950 105820 109992 105860
rect 109992 105820 109994 105860
rect 109702 105778 109826 105820
rect 109870 105778 109994 105820
rect 124822 105860 124946 105902
rect 124990 105860 125114 105902
rect 124822 105820 124824 105860
rect 124824 105820 124866 105860
rect 124866 105820 124906 105860
rect 124906 105820 124946 105860
rect 124990 105820 125030 105860
rect 125030 105820 125070 105860
rect 125070 105820 125112 105860
rect 125112 105820 125114 105860
rect 124822 105778 124946 105820
rect 124990 105778 125114 105820
rect 139942 105860 140066 105902
rect 140110 105860 140234 105902
rect 139942 105820 139944 105860
rect 139944 105820 139986 105860
rect 139986 105820 140026 105860
rect 140026 105820 140066 105860
rect 140110 105820 140150 105860
rect 140150 105820 140190 105860
rect 140190 105820 140232 105860
rect 140232 105820 140234 105860
rect 139942 105778 140066 105820
rect 140110 105778 140234 105820
rect 78222 105104 78346 105146
rect 78390 105104 78514 105146
rect 78222 105064 78224 105104
rect 78224 105064 78266 105104
rect 78266 105064 78306 105104
rect 78306 105064 78346 105104
rect 78390 105064 78430 105104
rect 78430 105064 78470 105104
rect 78470 105064 78512 105104
rect 78512 105064 78514 105104
rect 78222 105022 78346 105064
rect 78390 105022 78514 105064
rect 93342 105104 93466 105146
rect 93510 105104 93634 105146
rect 93342 105064 93344 105104
rect 93344 105064 93386 105104
rect 93386 105064 93426 105104
rect 93426 105064 93466 105104
rect 93510 105064 93550 105104
rect 93550 105064 93590 105104
rect 93590 105064 93632 105104
rect 93632 105064 93634 105104
rect 93342 105022 93466 105064
rect 93510 105022 93634 105064
rect 108462 105104 108586 105146
rect 108630 105104 108754 105146
rect 108462 105064 108464 105104
rect 108464 105064 108506 105104
rect 108506 105064 108546 105104
rect 108546 105064 108586 105104
rect 108630 105064 108670 105104
rect 108670 105064 108710 105104
rect 108710 105064 108752 105104
rect 108752 105064 108754 105104
rect 108462 105022 108586 105064
rect 108630 105022 108754 105064
rect 123582 105104 123706 105146
rect 123750 105104 123874 105146
rect 123582 105064 123584 105104
rect 123584 105064 123626 105104
rect 123626 105064 123666 105104
rect 123666 105064 123706 105104
rect 123750 105064 123790 105104
rect 123790 105064 123830 105104
rect 123830 105064 123872 105104
rect 123872 105064 123874 105104
rect 123582 105022 123706 105064
rect 123750 105022 123874 105064
rect 138702 105104 138826 105146
rect 138870 105104 138994 105146
rect 138702 105064 138704 105104
rect 138704 105064 138746 105104
rect 138746 105064 138786 105104
rect 138786 105064 138826 105104
rect 138870 105064 138910 105104
rect 138910 105064 138950 105104
rect 138950 105064 138992 105104
rect 138992 105064 138994 105104
rect 138702 105022 138826 105064
rect 138870 105022 138994 105064
rect 79462 104348 79586 104390
rect 79630 104348 79754 104390
rect 79462 104308 79464 104348
rect 79464 104308 79506 104348
rect 79506 104308 79546 104348
rect 79546 104308 79586 104348
rect 79630 104308 79670 104348
rect 79670 104308 79710 104348
rect 79710 104308 79752 104348
rect 79752 104308 79754 104348
rect 79462 104266 79586 104308
rect 79630 104266 79754 104308
rect 94582 104348 94706 104390
rect 94750 104348 94874 104390
rect 94582 104308 94584 104348
rect 94584 104308 94626 104348
rect 94626 104308 94666 104348
rect 94666 104308 94706 104348
rect 94750 104308 94790 104348
rect 94790 104308 94830 104348
rect 94830 104308 94872 104348
rect 94872 104308 94874 104348
rect 94582 104266 94706 104308
rect 94750 104266 94874 104308
rect 109702 104348 109826 104390
rect 109870 104348 109994 104390
rect 109702 104308 109704 104348
rect 109704 104308 109746 104348
rect 109746 104308 109786 104348
rect 109786 104308 109826 104348
rect 109870 104308 109910 104348
rect 109910 104308 109950 104348
rect 109950 104308 109992 104348
rect 109992 104308 109994 104348
rect 109702 104266 109826 104308
rect 109870 104266 109994 104308
rect 124822 104348 124946 104390
rect 124990 104348 125114 104390
rect 124822 104308 124824 104348
rect 124824 104308 124866 104348
rect 124866 104308 124906 104348
rect 124906 104308 124946 104348
rect 124990 104308 125030 104348
rect 125030 104308 125070 104348
rect 125070 104308 125112 104348
rect 125112 104308 125114 104348
rect 124822 104266 124946 104308
rect 124990 104266 125114 104308
rect 139942 104348 140066 104390
rect 140110 104348 140234 104390
rect 139942 104308 139944 104348
rect 139944 104308 139986 104348
rect 139986 104308 140026 104348
rect 140026 104308 140066 104348
rect 140110 104308 140150 104348
rect 140150 104308 140190 104348
rect 140190 104308 140232 104348
rect 140232 104308 140234 104348
rect 139942 104266 140066 104308
rect 140110 104266 140234 104308
rect 78222 103592 78346 103634
rect 78390 103592 78514 103634
rect 78222 103552 78224 103592
rect 78224 103552 78266 103592
rect 78266 103552 78306 103592
rect 78306 103552 78346 103592
rect 78390 103552 78430 103592
rect 78430 103552 78470 103592
rect 78470 103552 78512 103592
rect 78512 103552 78514 103592
rect 78222 103510 78346 103552
rect 78390 103510 78514 103552
rect 93342 103592 93466 103634
rect 93510 103592 93634 103634
rect 93342 103552 93344 103592
rect 93344 103552 93386 103592
rect 93386 103552 93426 103592
rect 93426 103552 93466 103592
rect 93510 103552 93550 103592
rect 93550 103552 93590 103592
rect 93590 103552 93632 103592
rect 93632 103552 93634 103592
rect 93342 103510 93466 103552
rect 93510 103510 93634 103552
rect 108462 103592 108586 103634
rect 108630 103592 108754 103634
rect 108462 103552 108464 103592
rect 108464 103552 108506 103592
rect 108506 103552 108546 103592
rect 108546 103552 108586 103592
rect 108630 103552 108670 103592
rect 108670 103552 108710 103592
rect 108710 103552 108752 103592
rect 108752 103552 108754 103592
rect 108462 103510 108586 103552
rect 108630 103510 108754 103552
rect 123582 103592 123706 103634
rect 123750 103592 123874 103634
rect 123582 103552 123584 103592
rect 123584 103552 123626 103592
rect 123626 103552 123666 103592
rect 123666 103552 123706 103592
rect 123750 103552 123790 103592
rect 123790 103552 123830 103592
rect 123830 103552 123872 103592
rect 123872 103552 123874 103592
rect 123582 103510 123706 103552
rect 123750 103510 123874 103552
rect 138702 103592 138826 103634
rect 138870 103592 138994 103634
rect 138702 103552 138704 103592
rect 138704 103552 138746 103592
rect 138746 103552 138786 103592
rect 138786 103552 138826 103592
rect 138870 103552 138910 103592
rect 138910 103552 138950 103592
rect 138950 103552 138992 103592
rect 138992 103552 138994 103592
rect 138702 103510 138826 103552
rect 138870 103510 138994 103552
rect 79462 102836 79586 102878
rect 79630 102836 79754 102878
rect 79462 102796 79464 102836
rect 79464 102796 79506 102836
rect 79506 102796 79546 102836
rect 79546 102796 79586 102836
rect 79630 102796 79670 102836
rect 79670 102796 79710 102836
rect 79710 102796 79752 102836
rect 79752 102796 79754 102836
rect 79462 102754 79586 102796
rect 79630 102754 79754 102796
rect 94582 102836 94706 102878
rect 94750 102836 94874 102878
rect 94582 102796 94584 102836
rect 94584 102796 94626 102836
rect 94626 102796 94666 102836
rect 94666 102796 94706 102836
rect 94750 102796 94790 102836
rect 94790 102796 94830 102836
rect 94830 102796 94872 102836
rect 94872 102796 94874 102836
rect 94582 102754 94706 102796
rect 94750 102754 94874 102796
rect 109702 102836 109826 102878
rect 109870 102836 109994 102878
rect 109702 102796 109704 102836
rect 109704 102796 109746 102836
rect 109746 102796 109786 102836
rect 109786 102796 109826 102836
rect 109870 102796 109910 102836
rect 109910 102796 109950 102836
rect 109950 102796 109992 102836
rect 109992 102796 109994 102836
rect 109702 102754 109826 102796
rect 109870 102754 109994 102796
rect 124822 102836 124946 102878
rect 124990 102836 125114 102878
rect 124822 102796 124824 102836
rect 124824 102796 124866 102836
rect 124866 102796 124906 102836
rect 124906 102796 124946 102836
rect 124990 102796 125030 102836
rect 125030 102796 125070 102836
rect 125070 102796 125112 102836
rect 125112 102796 125114 102836
rect 124822 102754 124946 102796
rect 124990 102754 125114 102796
rect 139942 102836 140066 102878
rect 140110 102836 140234 102878
rect 139942 102796 139944 102836
rect 139944 102796 139986 102836
rect 139986 102796 140026 102836
rect 140026 102796 140066 102836
rect 140110 102796 140150 102836
rect 140150 102796 140190 102836
rect 140190 102796 140232 102836
rect 140232 102796 140234 102836
rect 139942 102754 140066 102796
rect 140110 102754 140234 102796
rect 78222 102080 78346 102122
rect 78390 102080 78514 102122
rect 78222 102040 78224 102080
rect 78224 102040 78266 102080
rect 78266 102040 78306 102080
rect 78306 102040 78346 102080
rect 78390 102040 78430 102080
rect 78430 102040 78470 102080
rect 78470 102040 78512 102080
rect 78512 102040 78514 102080
rect 78222 101998 78346 102040
rect 78390 101998 78514 102040
rect 93342 102080 93466 102122
rect 93510 102080 93634 102122
rect 93342 102040 93344 102080
rect 93344 102040 93386 102080
rect 93386 102040 93426 102080
rect 93426 102040 93466 102080
rect 93510 102040 93550 102080
rect 93550 102040 93590 102080
rect 93590 102040 93632 102080
rect 93632 102040 93634 102080
rect 93342 101998 93466 102040
rect 93510 101998 93634 102040
rect 108462 102080 108586 102122
rect 108630 102080 108754 102122
rect 108462 102040 108464 102080
rect 108464 102040 108506 102080
rect 108506 102040 108546 102080
rect 108546 102040 108586 102080
rect 108630 102040 108670 102080
rect 108670 102040 108710 102080
rect 108710 102040 108752 102080
rect 108752 102040 108754 102080
rect 108462 101998 108586 102040
rect 108630 101998 108754 102040
rect 123582 102080 123706 102122
rect 123750 102080 123874 102122
rect 123582 102040 123584 102080
rect 123584 102040 123626 102080
rect 123626 102040 123666 102080
rect 123666 102040 123706 102080
rect 123750 102040 123790 102080
rect 123790 102040 123830 102080
rect 123830 102040 123872 102080
rect 123872 102040 123874 102080
rect 123582 101998 123706 102040
rect 123750 101998 123874 102040
rect 138702 102080 138826 102122
rect 138870 102080 138994 102122
rect 138702 102040 138704 102080
rect 138704 102040 138746 102080
rect 138746 102040 138786 102080
rect 138786 102040 138826 102080
rect 138870 102040 138910 102080
rect 138910 102040 138950 102080
rect 138950 102040 138992 102080
rect 138992 102040 138994 102080
rect 138702 101998 138826 102040
rect 138870 101998 138994 102040
rect 79462 101324 79586 101366
rect 79630 101324 79754 101366
rect 79462 101284 79464 101324
rect 79464 101284 79506 101324
rect 79506 101284 79546 101324
rect 79546 101284 79586 101324
rect 79630 101284 79670 101324
rect 79670 101284 79710 101324
rect 79710 101284 79752 101324
rect 79752 101284 79754 101324
rect 79462 101242 79586 101284
rect 79630 101242 79754 101284
rect 94582 101324 94706 101366
rect 94750 101324 94874 101366
rect 94582 101284 94584 101324
rect 94584 101284 94626 101324
rect 94626 101284 94666 101324
rect 94666 101284 94706 101324
rect 94750 101284 94790 101324
rect 94790 101284 94830 101324
rect 94830 101284 94872 101324
rect 94872 101284 94874 101324
rect 94582 101242 94706 101284
rect 94750 101242 94874 101284
rect 109702 101324 109826 101366
rect 109870 101324 109994 101366
rect 109702 101284 109704 101324
rect 109704 101284 109746 101324
rect 109746 101284 109786 101324
rect 109786 101284 109826 101324
rect 109870 101284 109910 101324
rect 109910 101284 109950 101324
rect 109950 101284 109992 101324
rect 109992 101284 109994 101324
rect 109702 101242 109826 101284
rect 109870 101242 109994 101284
rect 124822 101324 124946 101366
rect 124990 101324 125114 101366
rect 124822 101284 124824 101324
rect 124824 101284 124866 101324
rect 124866 101284 124906 101324
rect 124906 101284 124946 101324
rect 124990 101284 125030 101324
rect 125030 101284 125070 101324
rect 125070 101284 125112 101324
rect 125112 101284 125114 101324
rect 124822 101242 124946 101284
rect 124990 101242 125114 101284
rect 139942 101324 140066 101366
rect 140110 101324 140234 101366
rect 139942 101284 139944 101324
rect 139944 101284 139986 101324
rect 139986 101284 140026 101324
rect 140026 101284 140066 101324
rect 140110 101284 140150 101324
rect 140150 101284 140190 101324
rect 140190 101284 140232 101324
rect 140232 101284 140234 101324
rect 139942 101242 140066 101284
rect 140110 101242 140234 101284
rect 78222 100568 78346 100610
rect 78390 100568 78514 100610
rect 78222 100528 78224 100568
rect 78224 100528 78266 100568
rect 78266 100528 78306 100568
rect 78306 100528 78346 100568
rect 78390 100528 78430 100568
rect 78430 100528 78470 100568
rect 78470 100528 78512 100568
rect 78512 100528 78514 100568
rect 78222 100486 78346 100528
rect 78390 100486 78514 100528
rect 93342 100568 93466 100610
rect 93510 100568 93634 100610
rect 93342 100528 93344 100568
rect 93344 100528 93386 100568
rect 93386 100528 93426 100568
rect 93426 100528 93466 100568
rect 93510 100528 93550 100568
rect 93550 100528 93590 100568
rect 93590 100528 93632 100568
rect 93632 100528 93634 100568
rect 93342 100486 93466 100528
rect 93510 100486 93634 100528
rect 108462 100568 108586 100610
rect 108630 100568 108754 100610
rect 108462 100528 108464 100568
rect 108464 100528 108506 100568
rect 108506 100528 108546 100568
rect 108546 100528 108586 100568
rect 108630 100528 108670 100568
rect 108670 100528 108710 100568
rect 108710 100528 108752 100568
rect 108752 100528 108754 100568
rect 108462 100486 108586 100528
rect 108630 100486 108754 100528
rect 123582 100568 123706 100610
rect 123750 100568 123874 100610
rect 123582 100528 123584 100568
rect 123584 100528 123626 100568
rect 123626 100528 123666 100568
rect 123666 100528 123706 100568
rect 123750 100528 123790 100568
rect 123790 100528 123830 100568
rect 123830 100528 123872 100568
rect 123872 100528 123874 100568
rect 123582 100486 123706 100528
rect 123750 100486 123874 100528
rect 138702 100568 138826 100610
rect 138870 100568 138994 100610
rect 138702 100528 138704 100568
rect 138704 100528 138746 100568
rect 138746 100528 138786 100568
rect 138786 100528 138826 100568
rect 138870 100528 138910 100568
rect 138910 100528 138950 100568
rect 138950 100528 138992 100568
rect 138992 100528 138994 100568
rect 138702 100486 138826 100528
rect 138870 100486 138994 100528
rect 79462 99812 79586 99854
rect 79630 99812 79754 99854
rect 79462 99772 79464 99812
rect 79464 99772 79506 99812
rect 79506 99772 79546 99812
rect 79546 99772 79586 99812
rect 79630 99772 79670 99812
rect 79670 99772 79710 99812
rect 79710 99772 79752 99812
rect 79752 99772 79754 99812
rect 79462 99730 79586 99772
rect 79630 99730 79754 99772
rect 94582 99812 94706 99854
rect 94750 99812 94874 99854
rect 94582 99772 94584 99812
rect 94584 99772 94626 99812
rect 94626 99772 94666 99812
rect 94666 99772 94706 99812
rect 94750 99772 94790 99812
rect 94790 99772 94830 99812
rect 94830 99772 94872 99812
rect 94872 99772 94874 99812
rect 94582 99730 94706 99772
rect 94750 99730 94874 99772
rect 109702 99812 109826 99854
rect 109870 99812 109994 99854
rect 109702 99772 109704 99812
rect 109704 99772 109746 99812
rect 109746 99772 109786 99812
rect 109786 99772 109826 99812
rect 109870 99772 109910 99812
rect 109910 99772 109950 99812
rect 109950 99772 109992 99812
rect 109992 99772 109994 99812
rect 109702 99730 109826 99772
rect 109870 99730 109994 99772
rect 124822 99812 124946 99854
rect 124990 99812 125114 99854
rect 124822 99772 124824 99812
rect 124824 99772 124866 99812
rect 124866 99772 124906 99812
rect 124906 99772 124946 99812
rect 124990 99772 125030 99812
rect 125030 99772 125070 99812
rect 125070 99772 125112 99812
rect 125112 99772 125114 99812
rect 124822 99730 124946 99772
rect 124990 99730 125114 99772
rect 139942 99812 140066 99854
rect 140110 99812 140234 99854
rect 139942 99772 139944 99812
rect 139944 99772 139986 99812
rect 139986 99772 140026 99812
rect 140026 99772 140066 99812
rect 140110 99772 140150 99812
rect 140150 99772 140190 99812
rect 140190 99772 140232 99812
rect 140232 99772 140234 99812
rect 139942 99730 140066 99772
rect 140110 99730 140234 99772
rect 78222 99056 78346 99098
rect 78390 99056 78514 99098
rect 78222 99016 78224 99056
rect 78224 99016 78266 99056
rect 78266 99016 78306 99056
rect 78306 99016 78346 99056
rect 78390 99016 78430 99056
rect 78430 99016 78470 99056
rect 78470 99016 78512 99056
rect 78512 99016 78514 99056
rect 78222 98974 78346 99016
rect 78390 98974 78514 99016
rect 93342 99056 93466 99098
rect 93510 99056 93634 99098
rect 93342 99016 93344 99056
rect 93344 99016 93386 99056
rect 93386 99016 93426 99056
rect 93426 99016 93466 99056
rect 93510 99016 93550 99056
rect 93550 99016 93590 99056
rect 93590 99016 93632 99056
rect 93632 99016 93634 99056
rect 93342 98974 93466 99016
rect 93510 98974 93634 99016
rect 108462 99056 108586 99098
rect 108630 99056 108754 99098
rect 108462 99016 108464 99056
rect 108464 99016 108506 99056
rect 108506 99016 108546 99056
rect 108546 99016 108586 99056
rect 108630 99016 108670 99056
rect 108670 99016 108710 99056
rect 108710 99016 108752 99056
rect 108752 99016 108754 99056
rect 108462 98974 108586 99016
rect 108630 98974 108754 99016
rect 123582 99056 123706 99098
rect 123750 99056 123874 99098
rect 123582 99016 123584 99056
rect 123584 99016 123626 99056
rect 123626 99016 123666 99056
rect 123666 99016 123706 99056
rect 123750 99016 123790 99056
rect 123790 99016 123830 99056
rect 123830 99016 123872 99056
rect 123872 99016 123874 99056
rect 123582 98974 123706 99016
rect 123750 98974 123874 99016
rect 138702 99056 138826 99098
rect 138870 99056 138994 99098
rect 138702 99016 138704 99056
rect 138704 99016 138746 99056
rect 138746 99016 138786 99056
rect 138786 99016 138826 99056
rect 138870 99016 138910 99056
rect 138910 99016 138950 99056
rect 138950 99016 138992 99056
rect 138992 99016 138994 99056
rect 138702 98974 138826 99016
rect 138870 98974 138994 99016
rect 79462 98300 79586 98342
rect 79630 98300 79754 98342
rect 79462 98260 79464 98300
rect 79464 98260 79506 98300
rect 79506 98260 79546 98300
rect 79546 98260 79586 98300
rect 79630 98260 79670 98300
rect 79670 98260 79710 98300
rect 79710 98260 79752 98300
rect 79752 98260 79754 98300
rect 79462 98218 79586 98260
rect 79630 98218 79754 98260
rect 94582 98300 94706 98342
rect 94750 98300 94874 98342
rect 94582 98260 94584 98300
rect 94584 98260 94626 98300
rect 94626 98260 94666 98300
rect 94666 98260 94706 98300
rect 94750 98260 94790 98300
rect 94790 98260 94830 98300
rect 94830 98260 94872 98300
rect 94872 98260 94874 98300
rect 94582 98218 94706 98260
rect 94750 98218 94874 98260
rect 109702 98300 109826 98342
rect 109870 98300 109994 98342
rect 109702 98260 109704 98300
rect 109704 98260 109746 98300
rect 109746 98260 109786 98300
rect 109786 98260 109826 98300
rect 109870 98260 109910 98300
rect 109910 98260 109950 98300
rect 109950 98260 109992 98300
rect 109992 98260 109994 98300
rect 109702 98218 109826 98260
rect 109870 98218 109994 98260
rect 124822 98300 124946 98342
rect 124990 98300 125114 98342
rect 124822 98260 124824 98300
rect 124824 98260 124866 98300
rect 124866 98260 124906 98300
rect 124906 98260 124946 98300
rect 124990 98260 125030 98300
rect 125030 98260 125070 98300
rect 125070 98260 125112 98300
rect 125112 98260 125114 98300
rect 124822 98218 124946 98260
rect 124990 98218 125114 98260
rect 139942 98300 140066 98342
rect 140110 98300 140234 98342
rect 139942 98260 139944 98300
rect 139944 98260 139986 98300
rect 139986 98260 140026 98300
rect 140026 98260 140066 98300
rect 140110 98260 140150 98300
rect 140150 98260 140190 98300
rect 140190 98260 140232 98300
rect 140232 98260 140234 98300
rect 139942 98218 140066 98260
rect 140110 98218 140234 98260
rect 78222 97544 78346 97586
rect 78390 97544 78514 97586
rect 78222 97504 78224 97544
rect 78224 97504 78266 97544
rect 78266 97504 78306 97544
rect 78306 97504 78346 97544
rect 78390 97504 78430 97544
rect 78430 97504 78470 97544
rect 78470 97504 78512 97544
rect 78512 97504 78514 97544
rect 78222 97462 78346 97504
rect 78390 97462 78514 97504
rect 93342 97544 93466 97586
rect 93510 97544 93634 97586
rect 93342 97504 93344 97544
rect 93344 97504 93386 97544
rect 93386 97504 93426 97544
rect 93426 97504 93466 97544
rect 93510 97504 93550 97544
rect 93550 97504 93590 97544
rect 93590 97504 93632 97544
rect 93632 97504 93634 97544
rect 93342 97462 93466 97504
rect 93510 97462 93634 97504
rect 108462 97544 108586 97586
rect 108630 97544 108754 97586
rect 108462 97504 108464 97544
rect 108464 97504 108506 97544
rect 108506 97504 108546 97544
rect 108546 97504 108586 97544
rect 108630 97504 108670 97544
rect 108670 97504 108710 97544
rect 108710 97504 108752 97544
rect 108752 97504 108754 97544
rect 108462 97462 108586 97504
rect 108630 97462 108754 97504
rect 123582 97544 123706 97586
rect 123750 97544 123874 97586
rect 123582 97504 123584 97544
rect 123584 97504 123626 97544
rect 123626 97504 123666 97544
rect 123666 97504 123706 97544
rect 123750 97504 123790 97544
rect 123790 97504 123830 97544
rect 123830 97504 123872 97544
rect 123872 97504 123874 97544
rect 123582 97462 123706 97504
rect 123750 97462 123874 97504
rect 138702 97544 138826 97586
rect 138870 97544 138994 97586
rect 138702 97504 138704 97544
rect 138704 97504 138746 97544
rect 138746 97504 138786 97544
rect 138786 97504 138826 97544
rect 138870 97504 138910 97544
rect 138910 97504 138950 97544
rect 138950 97504 138992 97544
rect 138992 97504 138994 97544
rect 138702 97462 138826 97504
rect 138870 97462 138994 97504
rect 79462 96788 79586 96830
rect 79630 96788 79754 96830
rect 79462 96748 79464 96788
rect 79464 96748 79506 96788
rect 79506 96748 79546 96788
rect 79546 96748 79586 96788
rect 79630 96748 79670 96788
rect 79670 96748 79710 96788
rect 79710 96748 79752 96788
rect 79752 96748 79754 96788
rect 79462 96706 79586 96748
rect 79630 96706 79754 96748
rect 94582 96788 94706 96830
rect 94750 96788 94874 96830
rect 94582 96748 94584 96788
rect 94584 96748 94626 96788
rect 94626 96748 94666 96788
rect 94666 96748 94706 96788
rect 94750 96748 94790 96788
rect 94790 96748 94830 96788
rect 94830 96748 94872 96788
rect 94872 96748 94874 96788
rect 94582 96706 94706 96748
rect 94750 96706 94874 96748
rect 109702 96788 109826 96830
rect 109870 96788 109994 96830
rect 109702 96748 109704 96788
rect 109704 96748 109746 96788
rect 109746 96748 109786 96788
rect 109786 96748 109826 96788
rect 109870 96748 109910 96788
rect 109910 96748 109950 96788
rect 109950 96748 109992 96788
rect 109992 96748 109994 96788
rect 109702 96706 109826 96748
rect 109870 96706 109994 96748
rect 124822 96788 124946 96830
rect 124990 96788 125114 96830
rect 124822 96748 124824 96788
rect 124824 96748 124866 96788
rect 124866 96748 124906 96788
rect 124906 96748 124946 96788
rect 124990 96748 125030 96788
rect 125030 96748 125070 96788
rect 125070 96748 125112 96788
rect 125112 96748 125114 96788
rect 124822 96706 124946 96748
rect 124990 96706 125114 96748
rect 139942 96788 140066 96830
rect 140110 96788 140234 96830
rect 139942 96748 139944 96788
rect 139944 96748 139986 96788
rect 139986 96748 140026 96788
rect 140026 96748 140066 96788
rect 140110 96748 140150 96788
rect 140150 96748 140190 96788
rect 140190 96748 140232 96788
rect 140232 96748 140234 96788
rect 139942 96706 140066 96748
rect 140110 96706 140234 96748
rect 78222 96032 78346 96074
rect 78390 96032 78514 96074
rect 78222 95992 78224 96032
rect 78224 95992 78266 96032
rect 78266 95992 78306 96032
rect 78306 95992 78346 96032
rect 78390 95992 78430 96032
rect 78430 95992 78470 96032
rect 78470 95992 78512 96032
rect 78512 95992 78514 96032
rect 78222 95950 78346 95992
rect 78390 95950 78514 95992
rect 93342 96032 93466 96074
rect 93510 96032 93634 96074
rect 93342 95992 93344 96032
rect 93344 95992 93386 96032
rect 93386 95992 93426 96032
rect 93426 95992 93466 96032
rect 93510 95992 93550 96032
rect 93550 95992 93590 96032
rect 93590 95992 93632 96032
rect 93632 95992 93634 96032
rect 93342 95950 93466 95992
rect 93510 95950 93634 95992
rect 108462 96032 108586 96074
rect 108630 96032 108754 96074
rect 108462 95992 108464 96032
rect 108464 95992 108506 96032
rect 108506 95992 108546 96032
rect 108546 95992 108586 96032
rect 108630 95992 108670 96032
rect 108670 95992 108710 96032
rect 108710 95992 108752 96032
rect 108752 95992 108754 96032
rect 108462 95950 108586 95992
rect 108630 95950 108754 95992
rect 123582 96032 123706 96074
rect 123750 96032 123874 96074
rect 123582 95992 123584 96032
rect 123584 95992 123626 96032
rect 123626 95992 123666 96032
rect 123666 95992 123706 96032
rect 123750 95992 123790 96032
rect 123790 95992 123830 96032
rect 123830 95992 123872 96032
rect 123872 95992 123874 96032
rect 123582 95950 123706 95992
rect 123750 95950 123874 95992
rect 138702 96032 138826 96074
rect 138870 96032 138994 96074
rect 138702 95992 138704 96032
rect 138704 95992 138746 96032
rect 138746 95992 138786 96032
rect 138786 95992 138826 96032
rect 138870 95992 138910 96032
rect 138910 95992 138950 96032
rect 138950 95992 138992 96032
rect 138992 95992 138994 96032
rect 138702 95950 138826 95992
rect 138870 95950 138994 95992
rect 79462 95276 79586 95318
rect 79630 95276 79754 95318
rect 79462 95236 79464 95276
rect 79464 95236 79506 95276
rect 79506 95236 79546 95276
rect 79546 95236 79586 95276
rect 79630 95236 79670 95276
rect 79670 95236 79710 95276
rect 79710 95236 79752 95276
rect 79752 95236 79754 95276
rect 79462 95194 79586 95236
rect 79630 95194 79754 95236
rect 94582 95276 94706 95318
rect 94750 95276 94874 95318
rect 94582 95236 94584 95276
rect 94584 95236 94626 95276
rect 94626 95236 94666 95276
rect 94666 95236 94706 95276
rect 94750 95236 94790 95276
rect 94790 95236 94830 95276
rect 94830 95236 94872 95276
rect 94872 95236 94874 95276
rect 94582 95194 94706 95236
rect 94750 95194 94874 95236
rect 109702 95276 109826 95318
rect 109870 95276 109994 95318
rect 109702 95236 109704 95276
rect 109704 95236 109746 95276
rect 109746 95236 109786 95276
rect 109786 95236 109826 95276
rect 109870 95236 109910 95276
rect 109910 95236 109950 95276
rect 109950 95236 109992 95276
rect 109992 95236 109994 95276
rect 109702 95194 109826 95236
rect 109870 95194 109994 95236
rect 124822 95276 124946 95318
rect 124990 95276 125114 95318
rect 124822 95236 124824 95276
rect 124824 95236 124866 95276
rect 124866 95236 124906 95276
rect 124906 95236 124946 95276
rect 124990 95236 125030 95276
rect 125030 95236 125070 95276
rect 125070 95236 125112 95276
rect 125112 95236 125114 95276
rect 124822 95194 124946 95236
rect 124990 95194 125114 95236
rect 139942 95276 140066 95318
rect 140110 95276 140234 95318
rect 139942 95236 139944 95276
rect 139944 95236 139986 95276
rect 139986 95236 140026 95276
rect 140026 95236 140066 95276
rect 140110 95236 140150 95276
rect 140150 95236 140190 95276
rect 140190 95236 140232 95276
rect 140232 95236 140234 95276
rect 139942 95194 140066 95236
rect 140110 95194 140234 95236
rect 78222 94520 78346 94562
rect 78390 94520 78514 94562
rect 78222 94480 78224 94520
rect 78224 94480 78266 94520
rect 78266 94480 78306 94520
rect 78306 94480 78346 94520
rect 78390 94480 78430 94520
rect 78430 94480 78470 94520
rect 78470 94480 78512 94520
rect 78512 94480 78514 94520
rect 78222 94438 78346 94480
rect 78390 94438 78514 94480
rect 93342 94520 93466 94562
rect 93510 94520 93634 94562
rect 93342 94480 93344 94520
rect 93344 94480 93386 94520
rect 93386 94480 93426 94520
rect 93426 94480 93466 94520
rect 93510 94480 93550 94520
rect 93550 94480 93590 94520
rect 93590 94480 93632 94520
rect 93632 94480 93634 94520
rect 93342 94438 93466 94480
rect 93510 94438 93634 94480
rect 108462 94520 108586 94562
rect 108630 94520 108754 94562
rect 108462 94480 108464 94520
rect 108464 94480 108506 94520
rect 108506 94480 108546 94520
rect 108546 94480 108586 94520
rect 108630 94480 108670 94520
rect 108670 94480 108710 94520
rect 108710 94480 108752 94520
rect 108752 94480 108754 94520
rect 108462 94438 108586 94480
rect 108630 94438 108754 94480
rect 123582 94520 123706 94562
rect 123750 94520 123874 94562
rect 123582 94480 123584 94520
rect 123584 94480 123626 94520
rect 123626 94480 123666 94520
rect 123666 94480 123706 94520
rect 123750 94480 123790 94520
rect 123790 94480 123830 94520
rect 123830 94480 123872 94520
rect 123872 94480 123874 94520
rect 123582 94438 123706 94480
rect 123750 94438 123874 94480
rect 138702 94520 138826 94562
rect 138870 94520 138994 94562
rect 138702 94480 138704 94520
rect 138704 94480 138746 94520
rect 138746 94480 138786 94520
rect 138786 94480 138826 94520
rect 138870 94480 138910 94520
rect 138910 94480 138950 94520
rect 138950 94480 138992 94520
rect 138992 94480 138994 94520
rect 138702 94438 138826 94480
rect 138870 94438 138994 94480
rect 79462 93764 79586 93806
rect 79630 93764 79754 93806
rect 79462 93724 79464 93764
rect 79464 93724 79506 93764
rect 79506 93724 79546 93764
rect 79546 93724 79586 93764
rect 79630 93724 79670 93764
rect 79670 93724 79710 93764
rect 79710 93724 79752 93764
rect 79752 93724 79754 93764
rect 79462 93682 79586 93724
rect 79630 93682 79754 93724
rect 94582 93764 94706 93806
rect 94750 93764 94874 93806
rect 94582 93724 94584 93764
rect 94584 93724 94626 93764
rect 94626 93724 94666 93764
rect 94666 93724 94706 93764
rect 94750 93724 94790 93764
rect 94790 93724 94830 93764
rect 94830 93724 94872 93764
rect 94872 93724 94874 93764
rect 94582 93682 94706 93724
rect 94750 93682 94874 93724
rect 109702 93764 109826 93806
rect 109870 93764 109994 93806
rect 109702 93724 109704 93764
rect 109704 93724 109746 93764
rect 109746 93724 109786 93764
rect 109786 93724 109826 93764
rect 109870 93724 109910 93764
rect 109910 93724 109950 93764
rect 109950 93724 109992 93764
rect 109992 93724 109994 93764
rect 109702 93682 109826 93724
rect 109870 93682 109994 93724
rect 124822 93764 124946 93806
rect 124990 93764 125114 93806
rect 124822 93724 124824 93764
rect 124824 93724 124866 93764
rect 124866 93724 124906 93764
rect 124906 93724 124946 93764
rect 124990 93724 125030 93764
rect 125030 93724 125070 93764
rect 125070 93724 125112 93764
rect 125112 93724 125114 93764
rect 124822 93682 124946 93724
rect 124990 93682 125114 93724
rect 139942 93764 140066 93806
rect 140110 93764 140234 93806
rect 139942 93724 139944 93764
rect 139944 93724 139986 93764
rect 139986 93724 140026 93764
rect 140026 93724 140066 93764
rect 140110 93724 140150 93764
rect 140150 93724 140190 93764
rect 140190 93724 140232 93764
rect 140232 93724 140234 93764
rect 139942 93682 140066 93724
rect 140110 93682 140234 93724
rect 78222 93008 78346 93050
rect 78390 93008 78514 93050
rect 78222 92968 78224 93008
rect 78224 92968 78266 93008
rect 78266 92968 78306 93008
rect 78306 92968 78346 93008
rect 78390 92968 78430 93008
rect 78430 92968 78470 93008
rect 78470 92968 78512 93008
rect 78512 92968 78514 93008
rect 78222 92926 78346 92968
rect 78390 92926 78514 92968
rect 93342 93008 93466 93050
rect 93510 93008 93634 93050
rect 93342 92968 93344 93008
rect 93344 92968 93386 93008
rect 93386 92968 93426 93008
rect 93426 92968 93466 93008
rect 93510 92968 93550 93008
rect 93550 92968 93590 93008
rect 93590 92968 93632 93008
rect 93632 92968 93634 93008
rect 93342 92926 93466 92968
rect 93510 92926 93634 92968
rect 108462 93008 108586 93050
rect 108630 93008 108754 93050
rect 108462 92968 108464 93008
rect 108464 92968 108506 93008
rect 108506 92968 108546 93008
rect 108546 92968 108586 93008
rect 108630 92968 108670 93008
rect 108670 92968 108710 93008
rect 108710 92968 108752 93008
rect 108752 92968 108754 93008
rect 108462 92926 108586 92968
rect 108630 92926 108754 92968
rect 123582 93008 123706 93050
rect 123750 93008 123874 93050
rect 123582 92968 123584 93008
rect 123584 92968 123626 93008
rect 123626 92968 123666 93008
rect 123666 92968 123706 93008
rect 123750 92968 123790 93008
rect 123790 92968 123830 93008
rect 123830 92968 123872 93008
rect 123872 92968 123874 93008
rect 123582 92926 123706 92968
rect 123750 92926 123874 92968
rect 138702 93008 138826 93050
rect 138870 93008 138994 93050
rect 138702 92968 138704 93008
rect 138704 92968 138746 93008
rect 138746 92968 138786 93008
rect 138786 92968 138826 93008
rect 138870 92968 138910 93008
rect 138910 92968 138950 93008
rect 138950 92968 138992 93008
rect 138992 92968 138994 93008
rect 138702 92926 138826 92968
rect 138870 92926 138994 92968
rect 79462 92252 79586 92294
rect 79630 92252 79754 92294
rect 79462 92212 79464 92252
rect 79464 92212 79506 92252
rect 79506 92212 79546 92252
rect 79546 92212 79586 92252
rect 79630 92212 79670 92252
rect 79670 92212 79710 92252
rect 79710 92212 79752 92252
rect 79752 92212 79754 92252
rect 79462 92170 79586 92212
rect 79630 92170 79754 92212
rect 94582 92252 94706 92294
rect 94750 92252 94874 92294
rect 94582 92212 94584 92252
rect 94584 92212 94626 92252
rect 94626 92212 94666 92252
rect 94666 92212 94706 92252
rect 94750 92212 94790 92252
rect 94790 92212 94830 92252
rect 94830 92212 94872 92252
rect 94872 92212 94874 92252
rect 94582 92170 94706 92212
rect 94750 92170 94874 92212
rect 109702 92252 109826 92294
rect 109870 92252 109994 92294
rect 109702 92212 109704 92252
rect 109704 92212 109746 92252
rect 109746 92212 109786 92252
rect 109786 92212 109826 92252
rect 109870 92212 109910 92252
rect 109910 92212 109950 92252
rect 109950 92212 109992 92252
rect 109992 92212 109994 92252
rect 109702 92170 109826 92212
rect 109870 92170 109994 92212
rect 124822 92252 124946 92294
rect 124990 92252 125114 92294
rect 124822 92212 124824 92252
rect 124824 92212 124866 92252
rect 124866 92212 124906 92252
rect 124906 92212 124946 92252
rect 124990 92212 125030 92252
rect 125030 92212 125070 92252
rect 125070 92212 125112 92252
rect 125112 92212 125114 92252
rect 124822 92170 124946 92212
rect 124990 92170 125114 92212
rect 139942 92252 140066 92294
rect 140110 92252 140234 92294
rect 139942 92212 139944 92252
rect 139944 92212 139986 92252
rect 139986 92212 140026 92252
rect 140026 92212 140066 92252
rect 140110 92212 140150 92252
rect 140150 92212 140190 92252
rect 140190 92212 140232 92252
rect 140232 92212 140234 92252
rect 139942 92170 140066 92212
rect 140110 92170 140234 92212
rect 78222 91496 78346 91538
rect 78390 91496 78514 91538
rect 78222 91456 78224 91496
rect 78224 91456 78266 91496
rect 78266 91456 78306 91496
rect 78306 91456 78346 91496
rect 78390 91456 78430 91496
rect 78430 91456 78470 91496
rect 78470 91456 78512 91496
rect 78512 91456 78514 91496
rect 78222 91414 78346 91456
rect 78390 91414 78514 91456
rect 93342 91496 93466 91538
rect 93510 91496 93634 91538
rect 93342 91456 93344 91496
rect 93344 91456 93386 91496
rect 93386 91456 93426 91496
rect 93426 91456 93466 91496
rect 93510 91456 93550 91496
rect 93550 91456 93590 91496
rect 93590 91456 93632 91496
rect 93632 91456 93634 91496
rect 93342 91414 93466 91456
rect 93510 91414 93634 91456
rect 108462 91496 108586 91538
rect 108630 91496 108754 91538
rect 108462 91456 108464 91496
rect 108464 91456 108506 91496
rect 108506 91456 108546 91496
rect 108546 91456 108586 91496
rect 108630 91456 108670 91496
rect 108670 91456 108710 91496
rect 108710 91456 108752 91496
rect 108752 91456 108754 91496
rect 108462 91414 108586 91456
rect 108630 91414 108754 91456
rect 123582 91496 123706 91538
rect 123750 91496 123874 91538
rect 123582 91456 123584 91496
rect 123584 91456 123626 91496
rect 123626 91456 123666 91496
rect 123666 91456 123706 91496
rect 123750 91456 123790 91496
rect 123790 91456 123830 91496
rect 123830 91456 123872 91496
rect 123872 91456 123874 91496
rect 123582 91414 123706 91456
rect 123750 91414 123874 91456
rect 138702 91496 138826 91538
rect 138870 91496 138994 91538
rect 138702 91456 138704 91496
rect 138704 91456 138746 91496
rect 138746 91456 138786 91496
rect 138786 91456 138826 91496
rect 138870 91456 138910 91496
rect 138910 91456 138950 91496
rect 138950 91456 138992 91496
rect 138992 91456 138994 91496
rect 138702 91414 138826 91456
rect 138870 91414 138994 91456
rect 79462 90740 79586 90782
rect 79630 90740 79754 90782
rect 79462 90700 79464 90740
rect 79464 90700 79506 90740
rect 79506 90700 79546 90740
rect 79546 90700 79586 90740
rect 79630 90700 79670 90740
rect 79670 90700 79710 90740
rect 79710 90700 79752 90740
rect 79752 90700 79754 90740
rect 79462 90658 79586 90700
rect 79630 90658 79754 90700
rect 94582 90740 94706 90782
rect 94750 90740 94874 90782
rect 94582 90700 94584 90740
rect 94584 90700 94626 90740
rect 94626 90700 94666 90740
rect 94666 90700 94706 90740
rect 94750 90700 94790 90740
rect 94790 90700 94830 90740
rect 94830 90700 94872 90740
rect 94872 90700 94874 90740
rect 94582 90658 94706 90700
rect 94750 90658 94874 90700
rect 109702 90740 109826 90782
rect 109870 90740 109994 90782
rect 109702 90700 109704 90740
rect 109704 90700 109746 90740
rect 109746 90700 109786 90740
rect 109786 90700 109826 90740
rect 109870 90700 109910 90740
rect 109910 90700 109950 90740
rect 109950 90700 109992 90740
rect 109992 90700 109994 90740
rect 109702 90658 109826 90700
rect 109870 90658 109994 90700
rect 124822 90740 124946 90782
rect 124990 90740 125114 90782
rect 124822 90700 124824 90740
rect 124824 90700 124866 90740
rect 124866 90700 124906 90740
rect 124906 90700 124946 90740
rect 124990 90700 125030 90740
rect 125030 90700 125070 90740
rect 125070 90700 125112 90740
rect 125112 90700 125114 90740
rect 124822 90658 124946 90700
rect 124990 90658 125114 90700
rect 139942 90740 140066 90782
rect 140110 90740 140234 90782
rect 139942 90700 139944 90740
rect 139944 90700 139986 90740
rect 139986 90700 140026 90740
rect 140026 90700 140066 90740
rect 140110 90700 140150 90740
rect 140150 90700 140190 90740
rect 140190 90700 140232 90740
rect 140232 90700 140234 90740
rect 139942 90658 140066 90700
rect 140110 90658 140234 90700
rect 78222 89984 78346 90026
rect 78390 89984 78514 90026
rect 78222 89944 78224 89984
rect 78224 89944 78266 89984
rect 78266 89944 78306 89984
rect 78306 89944 78346 89984
rect 78390 89944 78430 89984
rect 78430 89944 78470 89984
rect 78470 89944 78512 89984
rect 78512 89944 78514 89984
rect 78222 89902 78346 89944
rect 78390 89902 78514 89944
rect 93342 89984 93466 90026
rect 93510 89984 93634 90026
rect 93342 89944 93344 89984
rect 93344 89944 93386 89984
rect 93386 89944 93426 89984
rect 93426 89944 93466 89984
rect 93510 89944 93550 89984
rect 93550 89944 93590 89984
rect 93590 89944 93632 89984
rect 93632 89944 93634 89984
rect 93342 89902 93466 89944
rect 93510 89902 93634 89944
rect 108462 89984 108586 90026
rect 108630 89984 108754 90026
rect 108462 89944 108464 89984
rect 108464 89944 108506 89984
rect 108506 89944 108546 89984
rect 108546 89944 108586 89984
rect 108630 89944 108670 89984
rect 108670 89944 108710 89984
rect 108710 89944 108752 89984
rect 108752 89944 108754 89984
rect 108462 89902 108586 89944
rect 108630 89902 108754 89944
rect 123582 89984 123706 90026
rect 123750 89984 123874 90026
rect 123582 89944 123584 89984
rect 123584 89944 123626 89984
rect 123626 89944 123666 89984
rect 123666 89944 123706 89984
rect 123750 89944 123790 89984
rect 123790 89944 123830 89984
rect 123830 89944 123872 89984
rect 123872 89944 123874 89984
rect 123582 89902 123706 89944
rect 123750 89902 123874 89944
rect 138702 89984 138826 90026
rect 138870 89984 138994 90026
rect 138702 89944 138704 89984
rect 138704 89944 138746 89984
rect 138746 89944 138786 89984
rect 138786 89944 138826 89984
rect 138870 89944 138910 89984
rect 138910 89944 138950 89984
rect 138950 89944 138992 89984
rect 138992 89944 138994 89984
rect 138702 89902 138826 89944
rect 138870 89902 138994 89944
rect 79462 89228 79586 89270
rect 79630 89228 79754 89270
rect 79462 89188 79464 89228
rect 79464 89188 79506 89228
rect 79506 89188 79546 89228
rect 79546 89188 79586 89228
rect 79630 89188 79670 89228
rect 79670 89188 79710 89228
rect 79710 89188 79752 89228
rect 79752 89188 79754 89228
rect 79462 89146 79586 89188
rect 79630 89146 79754 89188
rect 94582 89228 94706 89270
rect 94750 89228 94874 89270
rect 94582 89188 94584 89228
rect 94584 89188 94626 89228
rect 94626 89188 94666 89228
rect 94666 89188 94706 89228
rect 94750 89188 94790 89228
rect 94790 89188 94830 89228
rect 94830 89188 94872 89228
rect 94872 89188 94874 89228
rect 94582 89146 94706 89188
rect 94750 89146 94874 89188
rect 109702 89228 109826 89270
rect 109870 89228 109994 89270
rect 109702 89188 109704 89228
rect 109704 89188 109746 89228
rect 109746 89188 109786 89228
rect 109786 89188 109826 89228
rect 109870 89188 109910 89228
rect 109910 89188 109950 89228
rect 109950 89188 109992 89228
rect 109992 89188 109994 89228
rect 109702 89146 109826 89188
rect 109870 89146 109994 89188
rect 124822 89228 124946 89270
rect 124990 89228 125114 89270
rect 124822 89188 124824 89228
rect 124824 89188 124866 89228
rect 124866 89188 124906 89228
rect 124906 89188 124946 89228
rect 124990 89188 125030 89228
rect 125030 89188 125070 89228
rect 125070 89188 125112 89228
rect 125112 89188 125114 89228
rect 124822 89146 124946 89188
rect 124990 89146 125114 89188
rect 139942 89228 140066 89270
rect 140110 89228 140234 89270
rect 139942 89188 139944 89228
rect 139944 89188 139986 89228
rect 139986 89188 140026 89228
rect 140026 89188 140066 89228
rect 140110 89188 140150 89228
rect 140150 89188 140190 89228
rect 140190 89188 140232 89228
rect 140232 89188 140234 89228
rect 139942 89146 140066 89188
rect 140110 89146 140234 89188
rect 78222 88472 78346 88514
rect 78390 88472 78514 88514
rect 78222 88432 78224 88472
rect 78224 88432 78266 88472
rect 78266 88432 78306 88472
rect 78306 88432 78346 88472
rect 78390 88432 78430 88472
rect 78430 88432 78470 88472
rect 78470 88432 78512 88472
rect 78512 88432 78514 88472
rect 78222 88390 78346 88432
rect 78390 88390 78514 88432
rect 93342 88472 93466 88514
rect 93510 88472 93634 88514
rect 93342 88432 93344 88472
rect 93344 88432 93386 88472
rect 93386 88432 93426 88472
rect 93426 88432 93466 88472
rect 93510 88432 93550 88472
rect 93550 88432 93590 88472
rect 93590 88432 93632 88472
rect 93632 88432 93634 88472
rect 93342 88390 93466 88432
rect 93510 88390 93634 88432
rect 108462 88472 108586 88514
rect 108630 88472 108754 88514
rect 108462 88432 108464 88472
rect 108464 88432 108506 88472
rect 108506 88432 108546 88472
rect 108546 88432 108586 88472
rect 108630 88432 108670 88472
rect 108670 88432 108710 88472
rect 108710 88432 108752 88472
rect 108752 88432 108754 88472
rect 108462 88390 108586 88432
rect 108630 88390 108754 88432
rect 123582 88472 123706 88514
rect 123750 88472 123874 88514
rect 123582 88432 123584 88472
rect 123584 88432 123626 88472
rect 123626 88432 123666 88472
rect 123666 88432 123706 88472
rect 123750 88432 123790 88472
rect 123790 88432 123830 88472
rect 123830 88432 123872 88472
rect 123872 88432 123874 88472
rect 123582 88390 123706 88432
rect 123750 88390 123874 88432
rect 138702 88472 138826 88514
rect 138870 88472 138994 88514
rect 138702 88432 138704 88472
rect 138704 88432 138746 88472
rect 138746 88432 138786 88472
rect 138786 88432 138826 88472
rect 138870 88432 138910 88472
rect 138910 88432 138950 88472
rect 138950 88432 138992 88472
rect 138992 88432 138994 88472
rect 138702 88390 138826 88432
rect 138870 88390 138994 88432
rect 79462 87716 79586 87758
rect 79630 87716 79754 87758
rect 79462 87676 79464 87716
rect 79464 87676 79506 87716
rect 79506 87676 79546 87716
rect 79546 87676 79586 87716
rect 79630 87676 79670 87716
rect 79670 87676 79710 87716
rect 79710 87676 79752 87716
rect 79752 87676 79754 87716
rect 79462 87634 79586 87676
rect 79630 87634 79754 87676
rect 94582 87716 94706 87758
rect 94750 87716 94874 87758
rect 94582 87676 94584 87716
rect 94584 87676 94626 87716
rect 94626 87676 94666 87716
rect 94666 87676 94706 87716
rect 94750 87676 94790 87716
rect 94790 87676 94830 87716
rect 94830 87676 94872 87716
rect 94872 87676 94874 87716
rect 94582 87634 94706 87676
rect 94750 87634 94874 87676
rect 109702 87716 109826 87758
rect 109870 87716 109994 87758
rect 109702 87676 109704 87716
rect 109704 87676 109746 87716
rect 109746 87676 109786 87716
rect 109786 87676 109826 87716
rect 109870 87676 109910 87716
rect 109910 87676 109950 87716
rect 109950 87676 109992 87716
rect 109992 87676 109994 87716
rect 109702 87634 109826 87676
rect 109870 87634 109994 87676
rect 124822 87716 124946 87758
rect 124990 87716 125114 87758
rect 124822 87676 124824 87716
rect 124824 87676 124866 87716
rect 124866 87676 124906 87716
rect 124906 87676 124946 87716
rect 124990 87676 125030 87716
rect 125030 87676 125070 87716
rect 125070 87676 125112 87716
rect 125112 87676 125114 87716
rect 124822 87634 124946 87676
rect 124990 87634 125114 87676
rect 139942 87716 140066 87758
rect 140110 87716 140234 87758
rect 139942 87676 139944 87716
rect 139944 87676 139986 87716
rect 139986 87676 140026 87716
rect 140026 87676 140066 87716
rect 140110 87676 140150 87716
rect 140150 87676 140190 87716
rect 140190 87676 140232 87716
rect 140232 87676 140234 87716
rect 139942 87634 140066 87676
rect 140110 87634 140234 87676
rect 78222 86960 78346 87002
rect 78390 86960 78514 87002
rect 78222 86920 78224 86960
rect 78224 86920 78266 86960
rect 78266 86920 78306 86960
rect 78306 86920 78346 86960
rect 78390 86920 78430 86960
rect 78430 86920 78470 86960
rect 78470 86920 78512 86960
rect 78512 86920 78514 86960
rect 78222 86878 78346 86920
rect 78390 86878 78514 86920
rect 93342 86960 93466 87002
rect 93510 86960 93634 87002
rect 93342 86920 93344 86960
rect 93344 86920 93386 86960
rect 93386 86920 93426 86960
rect 93426 86920 93466 86960
rect 93510 86920 93550 86960
rect 93550 86920 93590 86960
rect 93590 86920 93632 86960
rect 93632 86920 93634 86960
rect 93342 86878 93466 86920
rect 93510 86878 93634 86920
rect 108462 86960 108586 87002
rect 108630 86960 108754 87002
rect 108462 86920 108464 86960
rect 108464 86920 108506 86960
rect 108506 86920 108546 86960
rect 108546 86920 108586 86960
rect 108630 86920 108670 86960
rect 108670 86920 108710 86960
rect 108710 86920 108752 86960
rect 108752 86920 108754 86960
rect 108462 86878 108586 86920
rect 108630 86878 108754 86920
rect 123582 86960 123706 87002
rect 123750 86960 123874 87002
rect 123582 86920 123584 86960
rect 123584 86920 123626 86960
rect 123626 86920 123666 86960
rect 123666 86920 123706 86960
rect 123750 86920 123790 86960
rect 123790 86920 123830 86960
rect 123830 86920 123872 86960
rect 123872 86920 123874 86960
rect 123582 86878 123706 86920
rect 123750 86878 123874 86920
rect 138702 86960 138826 87002
rect 138870 86960 138994 87002
rect 138702 86920 138704 86960
rect 138704 86920 138746 86960
rect 138746 86920 138786 86960
rect 138786 86920 138826 86960
rect 138870 86920 138910 86960
rect 138910 86920 138950 86960
rect 138950 86920 138992 86960
rect 138992 86920 138994 86960
rect 138702 86878 138826 86920
rect 138870 86878 138994 86920
rect 79462 86204 79586 86246
rect 79630 86204 79754 86246
rect 79462 86164 79464 86204
rect 79464 86164 79506 86204
rect 79506 86164 79546 86204
rect 79546 86164 79586 86204
rect 79630 86164 79670 86204
rect 79670 86164 79710 86204
rect 79710 86164 79752 86204
rect 79752 86164 79754 86204
rect 79462 86122 79586 86164
rect 79630 86122 79754 86164
rect 94582 86204 94706 86246
rect 94750 86204 94874 86246
rect 94582 86164 94584 86204
rect 94584 86164 94626 86204
rect 94626 86164 94666 86204
rect 94666 86164 94706 86204
rect 94750 86164 94790 86204
rect 94790 86164 94830 86204
rect 94830 86164 94872 86204
rect 94872 86164 94874 86204
rect 94582 86122 94706 86164
rect 94750 86122 94874 86164
rect 109702 86204 109826 86246
rect 109870 86204 109994 86246
rect 109702 86164 109704 86204
rect 109704 86164 109746 86204
rect 109746 86164 109786 86204
rect 109786 86164 109826 86204
rect 109870 86164 109910 86204
rect 109910 86164 109950 86204
rect 109950 86164 109992 86204
rect 109992 86164 109994 86204
rect 109702 86122 109826 86164
rect 109870 86122 109994 86164
rect 124822 86204 124946 86246
rect 124990 86204 125114 86246
rect 124822 86164 124824 86204
rect 124824 86164 124866 86204
rect 124866 86164 124906 86204
rect 124906 86164 124946 86204
rect 124990 86164 125030 86204
rect 125030 86164 125070 86204
rect 125070 86164 125112 86204
rect 125112 86164 125114 86204
rect 124822 86122 124946 86164
rect 124990 86122 125114 86164
rect 139942 86204 140066 86246
rect 140110 86204 140234 86246
rect 139942 86164 139944 86204
rect 139944 86164 139986 86204
rect 139986 86164 140026 86204
rect 140026 86164 140066 86204
rect 140110 86164 140150 86204
rect 140150 86164 140190 86204
rect 140190 86164 140232 86204
rect 140232 86164 140234 86204
rect 139942 86122 140066 86164
rect 140110 86122 140234 86164
rect 78222 85448 78346 85490
rect 78390 85448 78514 85490
rect 78222 85408 78224 85448
rect 78224 85408 78266 85448
rect 78266 85408 78306 85448
rect 78306 85408 78346 85448
rect 78390 85408 78430 85448
rect 78430 85408 78470 85448
rect 78470 85408 78512 85448
rect 78512 85408 78514 85448
rect 78222 85366 78346 85408
rect 78390 85366 78514 85408
rect 93342 85448 93466 85490
rect 93510 85448 93634 85490
rect 93342 85408 93344 85448
rect 93344 85408 93386 85448
rect 93386 85408 93426 85448
rect 93426 85408 93466 85448
rect 93510 85408 93550 85448
rect 93550 85408 93590 85448
rect 93590 85408 93632 85448
rect 93632 85408 93634 85448
rect 93342 85366 93466 85408
rect 93510 85366 93634 85408
rect 108462 85448 108586 85490
rect 108630 85448 108754 85490
rect 108462 85408 108464 85448
rect 108464 85408 108506 85448
rect 108506 85408 108546 85448
rect 108546 85408 108586 85448
rect 108630 85408 108670 85448
rect 108670 85408 108710 85448
rect 108710 85408 108752 85448
rect 108752 85408 108754 85448
rect 108462 85366 108586 85408
rect 108630 85366 108754 85408
rect 123582 85448 123706 85490
rect 123750 85448 123874 85490
rect 123582 85408 123584 85448
rect 123584 85408 123626 85448
rect 123626 85408 123666 85448
rect 123666 85408 123706 85448
rect 123750 85408 123790 85448
rect 123790 85408 123830 85448
rect 123830 85408 123872 85448
rect 123872 85408 123874 85448
rect 123582 85366 123706 85408
rect 123750 85366 123874 85408
rect 138702 85448 138826 85490
rect 138870 85448 138994 85490
rect 138702 85408 138704 85448
rect 138704 85408 138746 85448
rect 138746 85408 138786 85448
rect 138786 85408 138826 85448
rect 138870 85408 138910 85448
rect 138910 85408 138950 85448
rect 138950 85408 138992 85448
rect 138992 85408 138994 85448
rect 138702 85366 138826 85408
rect 138870 85366 138994 85408
rect 79462 84692 79586 84734
rect 79630 84692 79754 84734
rect 79462 84652 79464 84692
rect 79464 84652 79506 84692
rect 79506 84652 79546 84692
rect 79546 84652 79586 84692
rect 79630 84652 79670 84692
rect 79670 84652 79710 84692
rect 79710 84652 79752 84692
rect 79752 84652 79754 84692
rect 79462 84610 79586 84652
rect 79630 84610 79754 84652
rect 94582 84692 94706 84734
rect 94750 84692 94874 84734
rect 94582 84652 94584 84692
rect 94584 84652 94626 84692
rect 94626 84652 94666 84692
rect 94666 84652 94706 84692
rect 94750 84652 94790 84692
rect 94790 84652 94830 84692
rect 94830 84652 94872 84692
rect 94872 84652 94874 84692
rect 94582 84610 94706 84652
rect 94750 84610 94874 84652
rect 109702 84692 109826 84734
rect 109870 84692 109994 84734
rect 109702 84652 109704 84692
rect 109704 84652 109746 84692
rect 109746 84652 109786 84692
rect 109786 84652 109826 84692
rect 109870 84652 109910 84692
rect 109910 84652 109950 84692
rect 109950 84652 109992 84692
rect 109992 84652 109994 84692
rect 109702 84610 109826 84652
rect 109870 84610 109994 84652
rect 124822 84692 124946 84734
rect 124990 84692 125114 84734
rect 124822 84652 124824 84692
rect 124824 84652 124866 84692
rect 124866 84652 124906 84692
rect 124906 84652 124946 84692
rect 124990 84652 125030 84692
rect 125030 84652 125070 84692
rect 125070 84652 125112 84692
rect 125112 84652 125114 84692
rect 124822 84610 124946 84652
rect 124990 84610 125114 84652
rect 139942 84692 140066 84734
rect 140110 84692 140234 84734
rect 139942 84652 139944 84692
rect 139944 84652 139986 84692
rect 139986 84652 140026 84692
rect 140026 84652 140066 84692
rect 140110 84652 140150 84692
rect 140150 84652 140190 84692
rect 140190 84652 140232 84692
rect 140232 84652 140234 84692
rect 139942 84610 140066 84652
rect 140110 84610 140234 84652
rect 78222 83936 78346 83978
rect 78390 83936 78514 83978
rect 78222 83896 78224 83936
rect 78224 83896 78266 83936
rect 78266 83896 78306 83936
rect 78306 83896 78346 83936
rect 78390 83896 78430 83936
rect 78430 83896 78470 83936
rect 78470 83896 78512 83936
rect 78512 83896 78514 83936
rect 78222 83854 78346 83896
rect 78390 83854 78514 83896
rect 93342 83936 93466 83978
rect 93510 83936 93634 83978
rect 93342 83896 93344 83936
rect 93344 83896 93386 83936
rect 93386 83896 93426 83936
rect 93426 83896 93466 83936
rect 93510 83896 93550 83936
rect 93550 83896 93590 83936
rect 93590 83896 93632 83936
rect 93632 83896 93634 83936
rect 93342 83854 93466 83896
rect 93510 83854 93634 83896
rect 108462 83936 108586 83978
rect 108630 83936 108754 83978
rect 108462 83896 108464 83936
rect 108464 83896 108506 83936
rect 108506 83896 108546 83936
rect 108546 83896 108586 83936
rect 108630 83896 108670 83936
rect 108670 83896 108710 83936
rect 108710 83896 108752 83936
rect 108752 83896 108754 83936
rect 108462 83854 108586 83896
rect 108630 83854 108754 83896
rect 123582 83936 123706 83978
rect 123750 83936 123874 83978
rect 123582 83896 123584 83936
rect 123584 83896 123626 83936
rect 123626 83896 123666 83936
rect 123666 83896 123706 83936
rect 123750 83896 123790 83936
rect 123790 83896 123830 83936
rect 123830 83896 123872 83936
rect 123872 83896 123874 83936
rect 123582 83854 123706 83896
rect 123750 83854 123874 83896
rect 138702 83936 138826 83978
rect 138870 83936 138994 83978
rect 138702 83896 138704 83936
rect 138704 83896 138746 83936
rect 138746 83896 138786 83936
rect 138786 83896 138826 83936
rect 138870 83896 138910 83936
rect 138910 83896 138950 83936
rect 138950 83896 138992 83936
rect 138992 83896 138994 83936
rect 138702 83854 138826 83896
rect 138870 83854 138994 83896
rect 79462 83180 79586 83222
rect 79630 83180 79754 83222
rect 79462 83140 79464 83180
rect 79464 83140 79506 83180
rect 79506 83140 79546 83180
rect 79546 83140 79586 83180
rect 79630 83140 79670 83180
rect 79670 83140 79710 83180
rect 79710 83140 79752 83180
rect 79752 83140 79754 83180
rect 79462 83098 79586 83140
rect 79630 83098 79754 83140
rect 94582 83180 94706 83222
rect 94750 83180 94874 83222
rect 94582 83140 94584 83180
rect 94584 83140 94626 83180
rect 94626 83140 94666 83180
rect 94666 83140 94706 83180
rect 94750 83140 94790 83180
rect 94790 83140 94830 83180
rect 94830 83140 94872 83180
rect 94872 83140 94874 83180
rect 94582 83098 94706 83140
rect 94750 83098 94874 83140
rect 109702 83180 109826 83222
rect 109870 83180 109994 83222
rect 109702 83140 109704 83180
rect 109704 83140 109746 83180
rect 109746 83140 109786 83180
rect 109786 83140 109826 83180
rect 109870 83140 109910 83180
rect 109910 83140 109950 83180
rect 109950 83140 109992 83180
rect 109992 83140 109994 83180
rect 109702 83098 109826 83140
rect 109870 83098 109994 83140
rect 124822 83180 124946 83222
rect 124990 83180 125114 83222
rect 124822 83140 124824 83180
rect 124824 83140 124866 83180
rect 124866 83140 124906 83180
rect 124906 83140 124946 83180
rect 124990 83140 125030 83180
rect 125030 83140 125070 83180
rect 125070 83140 125112 83180
rect 125112 83140 125114 83180
rect 124822 83098 124946 83140
rect 124990 83098 125114 83140
rect 139942 83180 140066 83222
rect 140110 83180 140234 83222
rect 139942 83140 139944 83180
rect 139944 83140 139986 83180
rect 139986 83140 140026 83180
rect 140026 83140 140066 83180
rect 140110 83140 140150 83180
rect 140150 83140 140190 83180
rect 140190 83140 140232 83180
rect 140232 83140 140234 83180
rect 139942 83098 140066 83140
rect 140110 83098 140234 83140
rect 78222 82424 78346 82466
rect 78390 82424 78514 82466
rect 78222 82384 78224 82424
rect 78224 82384 78266 82424
rect 78266 82384 78306 82424
rect 78306 82384 78346 82424
rect 78390 82384 78430 82424
rect 78430 82384 78470 82424
rect 78470 82384 78512 82424
rect 78512 82384 78514 82424
rect 78222 82342 78346 82384
rect 78390 82342 78514 82384
rect 93342 82424 93466 82466
rect 93510 82424 93634 82466
rect 93342 82384 93344 82424
rect 93344 82384 93386 82424
rect 93386 82384 93426 82424
rect 93426 82384 93466 82424
rect 93510 82384 93550 82424
rect 93550 82384 93590 82424
rect 93590 82384 93632 82424
rect 93632 82384 93634 82424
rect 93342 82342 93466 82384
rect 93510 82342 93634 82384
rect 108462 82424 108586 82466
rect 108630 82424 108754 82466
rect 108462 82384 108464 82424
rect 108464 82384 108506 82424
rect 108506 82384 108546 82424
rect 108546 82384 108586 82424
rect 108630 82384 108670 82424
rect 108670 82384 108710 82424
rect 108710 82384 108752 82424
rect 108752 82384 108754 82424
rect 108462 82342 108586 82384
rect 108630 82342 108754 82384
rect 123582 82424 123706 82466
rect 123750 82424 123874 82466
rect 123582 82384 123584 82424
rect 123584 82384 123626 82424
rect 123626 82384 123666 82424
rect 123666 82384 123706 82424
rect 123750 82384 123790 82424
rect 123790 82384 123830 82424
rect 123830 82384 123872 82424
rect 123872 82384 123874 82424
rect 123582 82342 123706 82384
rect 123750 82342 123874 82384
rect 138702 82424 138826 82466
rect 138870 82424 138994 82466
rect 138702 82384 138704 82424
rect 138704 82384 138746 82424
rect 138746 82384 138786 82424
rect 138786 82384 138826 82424
rect 138870 82384 138910 82424
rect 138910 82384 138950 82424
rect 138950 82384 138992 82424
rect 138992 82384 138994 82424
rect 138702 82342 138826 82384
rect 138870 82342 138994 82384
rect 79462 81668 79586 81710
rect 79630 81668 79754 81710
rect 79462 81628 79464 81668
rect 79464 81628 79506 81668
rect 79506 81628 79546 81668
rect 79546 81628 79586 81668
rect 79630 81628 79670 81668
rect 79670 81628 79710 81668
rect 79710 81628 79752 81668
rect 79752 81628 79754 81668
rect 79462 81586 79586 81628
rect 79630 81586 79754 81628
rect 94582 81668 94706 81710
rect 94750 81668 94874 81710
rect 94582 81628 94584 81668
rect 94584 81628 94626 81668
rect 94626 81628 94666 81668
rect 94666 81628 94706 81668
rect 94750 81628 94790 81668
rect 94790 81628 94830 81668
rect 94830 81628 94872 81668
rect 94872 81628 94874 81668
rect 94582 81586 94706 81628
rect 94750 81586 94874 81628
rect 109702 81668 109826 81710
rect 109870 81668 109994 81710
rect 109702 81628 109704 81668
rect 109704 81628 109746 81668
rect 109746 81628 109786 81668
rect 109786 81628 109826 81668
rect 109870 81628 109910 81668
rect 109910 81628 109950 81668
rect 109950 81628 109992 81668
rect 109992 81628 109994 81668
rect 109702 81586 109826 81628
rect 109870 81586 109994 81628
rect 124822 81668 124946 81710
rect 124990 81668 125114 81710
rect 124822 81628 124824 81668
rect 124824 81628 124866 81668
rect 124866 81628 124906 81668
rect 124906 81628 124946 81668
rect 124990 81628 125030 81668
rect 125030 81628 125070 81668
rect 125070 81628 125112 81668
rect 125112 81628 125114 81668
rect 124822 81586 124946 81628
rect 124990 81586 125114 81628
rect 139942 81668 140066 81710
rect 140110 81668 140234 81710
rect 139942 81628 139944 81668
rect 139944 81628 139986 81668
rect 139986 81628 140026 81668
rect 140026 81628 140066 81668
rect 140110 81628 140150 81668
rect 140150 81628 140190 81668
rect 140190 81628 140232 81668
rect 140232 81628 140234 81668
rect 139942 81586 140066 81628
rect 140110 81586 140234 81628
rect 78222 80912 78346 80954
rect 78390 80912 78514 80954
rect 78222 80872 78224 80912
rect 78224 80872 78266 80912
rect 78266 80872 78306 80912
rect 78306 80872 78346 80912
rect 78390 80872 78430 80912
rect 78430 80872 78470 80912
rect 78470 80872 78512 80912
rect 78512 80872 78514 80912
rect 78222 80830 78346 80872
rect 78390 80830 78514 80872
rect 93342 80912 93466 80954
rect 93510 80912 93634 80954
rect 93342 80872 93344 80912
rect 93344 80872 93386 80912
rect 93386 80872 93426 80912
rect 93426 80872 93466 80912
rect 93510 80872 93550 80912
rect 93550 80872 93590 80912
rect 93590 80872 93632 80912
rect 93632 80872 93634 80912
rect 93342 80830 93466 80872
rect 93510 80830 93634 80872
rect 108462 80912 108586 80954
rect 108630 80912 108754 80954
rect 108462 80872 108464 80912
rect 108464 80872 108506 80912
rect 108506 80872 108546 80912
rect 108546 80872 108586 80912
rect 108630 80872 108670 80912
rect 108670 80872 108710 80912
rect 108710 80872 108752 80912
rect 108752 80872 108754 80912
rect 108462 80830 108586 80872
rect 108630 80830 108754 80872
rect 123582 80912 123706 80954
rect 123750 80912 123874 80954
rect 123582 80872 123584 80912
rect 123584 80872 123626 80912
rect 123626 80872 123666 80912
rect 123666 80872 123706 80912
rect 123750 80872 123790 80912
rect 123790 80872 123830 80912
rect 123830 80872 123872 80912
rect 123872 80872 123874 80912
rect 123582 80830 123706 80872
rect 123750 80830 123874 80872
rect 138702 80912 138826 80954
rect 138870 80912 138994 80954
rect 138702 80872 138704 80912
rect 138704 80872 138746 80912
rect 138746 80872 138786 80912
rect 138786 80872 138826 80912
rect 138870 80872 138910 80912
rect 138910 80872 138950 80912
rect 138950 80872 138992 80912
rect 138992 80872 138994 80912
rect 138702 80830 138826 80872
rect 138870 80830 138994 80872
rect 79462 80156 79586 80198
rect 79630 80156 79754 80198
rect 79462 80116 79464 80156
rect 79464 80116 79506 80156
rect 79506 80116 79546 80156
rect 79546 80116 79586 80156
rect 79630 80116 79670 80156
rect 79670 80116 79710 80156
rect 79710 80116 79752 80156
rect 79752 80116 79754 80156
rect 79462 80074 79586 80116
rect 79630 80074 79754 80116
rect 94582 80156 94706 80198
rect 94750 80156 94874 80198
rect 94582 80116 94584 80156
rect 94584 80116 94626 80156
rect 94626 80116 94666 80156
rect 94666 80116 94706 80156
rect 94750 80116 94790 80156
rect 94790 80116 94830 80156
rect 94830 80116 94872 80156
rect 94872 80116 94874 80156
rect 94582 80074 94706 80116
rect 94750 80074 94874 80116
rect 109702 80156 109826 80198
rect 109870 80156 109994 80198
rect 109702 80116 109704 80156
rect 109704 80116 109746 80156
rect 109746 80116 109786 80156
rect 109786 80116 109826 80156
rect 109870 80116 109910 80156
rect 109910 80116 109950 80156
rect 109950 80116 109992 80156
rect 109992 80116 109994 80156
rect 109702 80074 109826 80116
rect 109870 80074 109994 80116
rect 124822 80156 124946 80198
rect 124990 80156 125114 80198
rect 124822 80116 124824 80156
rect 124824 80116 124866 80156
rect 124866 80116 124906 80156
rect 124906 80116 124946 80156
rect 124990 80116 125030 80156
rect 125030 80116 125070 80156
rect 125070 80116 125112 80156
rect 125112 80116 125114 80156
rect 124822 80074 124946 80116
rect 124990 80074 125114 80116
rect 139942 80156 140066 80198
rect 140110 80156 140234 80198
rect 139942 80116 139944 80156
rect 139944 80116 139986 80156
rect 139986 80116 140026 80156
rect 140026 80116 140066 80156
rect 140110 80116 140150 80156
rect 140150 80116 140190 80156
rect 140190 80116 140232 80156
rect 140232 80116 140234 80156
rect 139942 80074 140066 80116
rect 140110 80074 140234 80116
rect 78222 79400 78346 79442
rect 78390 79400 78514 79442
rect 78222 79360 78224 79400
rect 78224 79360 78266 79400
rect 78266 79360 78306 79400
rect 78306 79360 78346 79400
rect 78390 79360 78430 79400
rect 78430 79360 78470 79400
rect 78470 79360 78512 79400
rect 78512 79360 78514 79400
rect 78222 79318 78346 79360
rect 78390 79318 78514 79360
rect 93342 79400 93466 79442
rect 93510 79400 93634 79442
rect 93342 79360 93344 79400
rect 93344 79360 93386 79400
rect 93386 79360 93426 79400
rect 93426 79360 93466 79400
rect 93510 79360 93550 79400
rect 93550 79360 93590 79400
rect 93590 79360 93632 79400
rect 93632 79360 93634 79400
rect 93342 79318 93466 79360
rect 93510 79318 93634 79360
rect 108462 79400 108586 79442
rect 108630 79400 108754 79442
rect 108462 79360 108464 79400
rect 108464 79360 108506 79400
rect 108506 79360 108546 79400
rect 108546 79360 108586 79400
rect 108630 79360 108670 79400
rect 108670 79360 108710 79400
rect 108710 79360 108752 79400
rect 108752 79360 108754 79400
rect 108462 79318 108586 79360
rect 108630 79318 108754 79360
rect 123582 79400 123706 79442
rect 123750 79400 123874 79442
rect 123582 79360 123584 79400
rect 123584 79360 123626 79400
rect 123626 79360 123666 79400
rect 123666 79360 123706 79400
rect 123750 79360 123790 79400
rect 123790 79360 123830 79400
rect 123830 79360 123872 79400
rect 123872 79360 123874 79400
rect 123582 79318 123706 79360
rect 123750 79318 123874 79360
rect 138702 79400 138826 79442
rect 138870 79400 138994 79442
rect 138702 79360 138704 79400
rect 138704 79360 138746 79400
rect 138746 79360 138786 79400
rect 138786 79360 138826 79400
rect 138870 79360 138910 79400
rect 138910 79360 138950 79400
rect 138950 79360 138992 79400
rect 138992 79360 138994 79400
rect 138702 79318 138826 79360
rect 138870 79318 138994 79360
rect 79462 78644 79586 78686
rect 79630 78644 79754 78686
rect 79462 78604 79464 78644
rect 79464 78604 79506 78644
rect 79506 78604 79546 78644
rect 79546 78604 79586 78644
rect 79630 78604 79670 78644
rect 79670 78604 79710 78644
rect 79710 78604 79752 78644
rect 79752 78604 79754 78644
rect 79462 78562 79586 78604
rect 79630 78562 79754 78604
rect 94582 78644 94706 78686
rect 94750 78644 94874 78686
rect 94582 78604 94584 78644
rect 94584 78604 94626 78644
rect 94626 78604 94666 78644
rect 94666 78604 94706 78644
rect 94750 78604 94790 78644
rect 94790 78604 94830 78644
rect 94830 78604 94872 78644
rect 94872 78604 94874 78644
rect 94582 78562 94706 78604
rect 94750 78562 94874 78604
rect 109702 78644 109826 78686
rect 109870 78644 109994 78686
rect 109702 78604 109704 78644
rect 109704 78604 109746 78644
rect 109746 78604 109786 78644
rect 109786 78604 109826 78644
rect 109870 78604 109910 78644
rect 109910 78604 109950 78644
rect 109950 78604 109992 78644
rect 109992 78604 109994 78644
rect 109702 78562 109826 78604
rect 109870 78562 109994 78604
rect 124822 78644 124946 78686
rect 124990 78644 125114 78686
rect 124822 78604 124824 78644
rect 124824 78604 124866 78644
rect 124866 78604 124906 78644
rect 124906 78604 124946 78644
rect 124990 78604 125030 78644
rect 125030 78604 125070 78644
rect 125070 78604 125112 78644
rect 125112 78604 125114 78644
rect 124822 78562 124946 78604
rect 124990 78562 125114 78604
rect 139942 78644 140066 78686
rect 140110 78644 140234 78686
rect 139942 78604 139944 78644
rect 139944 78604 139986 78644
rect 139986 78604 140026 78644
rect 140026 78604 140066 78644
rect 140110 78604 140150 78644
rect 140150 78604 140190 78644
rect 140190 78604 140232 78644
rect 140232 78604 140234 78644
rect 139942 78562 140066 78604
rect 140110 78562 140234 78604
rect 78222 77888 78346 77930
rect 78390 77888 78514 77930
rect 78222 77848 78224 77888
rect 78224 77848 78266 77888
rect 78266 77848 78306 77888
rect 78306 77848 78346 77888
rect 78390 77848 78430 77888
rect 78430 77848 78470 77888
rect 78470 77848 78512 77888
rect 78512 77848 78514 77888
rect 78222 77806 78346 77848
rect 78390 77806 78514 77848
rect 93342 77888 93466 77930
rect 93510 77888 93634 77930
rect 93342 77848 93344 77888
rect 93344 77848 93386 77888
rect 93386 77848 93426 77888
rect 93426 77848 93466 77888
rect 93510 77848 93550 77888
rect 93550 77848 93590 77888
rect 93590 77848 93632 77888
rect 93632 77848 93634 77888
rect 93342 77806 93466 77848
rect 93510 77806 93634 77848
rect 108462 77888 108586 77930
rect 108630 77888 108754 77930
rect 108462 77848 108464 77888
rect 108464 77848 108506 77888
rect 108506 77848 108546 77888
rect 108546 77848 108586 77888
rect 108630 77848 108670 77888
rect 108670 77848 108710 77888
rect 108710 77848 108752 77888
rect 108752 77848 108754 77888
rect 108462 77806 108586 77848
rect 108630 77806 108754 77848
rect 123582 77888 123706 77930
rect 123750 77888 123874 77930
rect 123582 77848 123584 77888
rect 123584 77848 123626 77888
rect 123626 77848 123666 77888
rect 123666 77848 123706 77888
rect 123750 77848 123790 77888
rect 123790 77848 123830 77888
rect 123830 77848 123872 77888
rect 123872 77848 123874 77888
rect 123582 77806 123706 77848
rect 123750 77806 123874 77848
rect 138702 77888 138826 77930
rect 138870 77888 138994 77930
rect 138702 77848 138704 77888
rect 138704 77848 138746 77888
rect 138746 77848 138786 77888
rect 138786 77848 138826 77888
rect 138870 77848 138910 77888
rect 138910 77848 138950 77888
rect 138950 77848 138992 77888
rect 138992 77848 138994 77888
rect 138702 77806 138826 77848
rect 138870 77806 138994 77848
rect 79462 77132 79586 77174
rect 79630 77132 79754 77174
rect 79462 77092 79464 77132
rect 79464 77092 79506 77132
rect 79506 77092 79546 77132
rect 79546 77092 79586 77132
rect 79630 77092 79670 77132
rect 79670 77092 79710 77132
rect 79710 77092 79752 77132
rect 79752 77092 79754 77132
rect 79462 77050 79586 77092
rect 79630 77050 79754 77092
rect 94582 77132 94706 77174
rect 94750 77132 94874 77174
rect 94582 77092 94584 77132
rect 94584 77092 94626 77132
rect 94626 77092 94666 77132
rect 94666 77092 94706 77132
rect 94750 77092 94790 77132
rect 94790 77092 94830 77132
rect 94830 77092 94872 77132
rect 94872 77092 94874 77132
rect 94582 77050 94706 77092
rect 94750 77050 94874 77092
rect 109702 77132 109826 77174
rect 109870 77132 109994 77174
rect 109702 77092 109704 77132
rect 109704 77092 109746 77132
rect 109746 77092 109786 77132
rect 109786 77092 109826 77132
rect 109870 77092 109910 77132
rect 109910 77092 109950 77132
rect 109950 77092 109992 77132
rect 109992 77092 109994 77132
rect 109702 77050 109826 77092
rect 109870 77050 109994 77092
rect 124822 77132 124946 77174
rect 124990 77132 125114 77174
rect 124822 77092 124824 77132
rect 124824 77092 124866 77132
rect 124866 77092 124906 77132
rect 124906 77092 124946 77132
rect 124990 77092 125030 77132
rect 125030 77092 125070 77132
rect 125070 77092 125112 77132
rect 125112 77092 125114 77132
rect 124822 77050 124946 77092
rect 124990 77050 125114 77092
rect 139942 77132 140066 77174
rect 140110 77132 140234 77174
rect 139942 77092 139944 77132
rect 139944 77092 139986 77132
rect 139986 77092 140026 77132
rect 140026 77092 140066 77132
rect 140110 77092 140150 77132
rect 140150 77092 140190 77132
rect 140190 77092 140232 77132
rect 140232 77092 140234 77132
rect 139942 77050 140066 77092
rect 140110 77050 140234 77092
rect 78222 76376 78346 76418
rect 78390 76376 78514 76418
rect 78222 76336 78224 76376
rect 78224 76336 78266 76376
rect 78266 76336 78306 76376
rect 78306 76336 78346 76376
rect 78390 76336 78430 76376
rect 78430 76336 78470 76376
rect 78470 76336 78512 76376
rect 78512 76336 78514 76376
rect 78222 76294 78346 76336
rect 78390 76294 78514 76336
rect 93342 76376 93466 76418
rect 93510 76376 93634 76418
rect 93342 76336 93344 76376
rect 93344 76336 93386 76376
rect 93386 76336 93426 76376
rect 93426 76336 93466 76376
rect 93510 76336 93550 76376
rect 93550 76336 93590 76376
rect 93590 76336 93632 76376
rect 93632 76336 93634 76376
rect 93342 76294 93466 76336
rect 93510 76294 93634 76336
rect 108462 76376 108586 76418
rect 108630 76376 108754 76418
rect 108462 76336 108464 76376
rect 108464 76336 108506 76376
rect 108506 76336 108546 76376
rect 108546 76336 108586 76376
rect 108630 76336 108670 76376
rect 108670 76336 108710 76376
rect 108710 76336 108752 76376
rect 108752 76336 108754 76376
rect 108462 76294 108586 76336
rect 108630 76294 108754 76336
rect 123582 76376 123706 76418
rect 123750 76376 123874 76418
rect 123582 76336 123584 76376
rect 123584 76336 123626 76376
rect 123626 76336 123666 76376
rect 123666 76336 123706 76376
rect 123750 76336 123790 76376
rect 123790 76336 123830 76376
rect 123830 76336 123872 76376
rect 123872 76336 123874 76376
rect 123582 76294 123706 76336
rect 123750 76294 123874 76336
rect 138702 76376 138826 76418
rect 138870 76376 138994 76418
rect 138702 76336 138704 76376
rect 138704 76336 138746 76376
rect 138746 76336 138786 76376
rect 138786 76336 138826 76376
rect 138870 76336 138910 76376
rect 138910 76336 138950 76376
rect 138950 76336 138992 76376
rect 138992 76336 138994 76376
rect 138702 76294 138826 76336
rect 138870 76294 138994 76336
rect 79462 75620 79586 75662
rect 79630 75620 79754 75662
rect 79462 75580 79464 75620
rect 79464 75580 79506 75620
rect 79506 75580 79546 75620
rect 79546 75580 79586 75620
rect 79630 75580 79670 75620
rect 79670 75580 79710 75620
rect 79710 75580 79752 75620
rect 79752 75580 79754 75620
rect 79462 75538 79586 75580
rect 79630 75538 79754 75580
rect 94582 75620 94706 75662
rect 94750 75620 94874 75662
rect 94582 75580 94584 75620
rect 94584 75580 94626 75620
rect 94626 75580 94666 75620
rect 94666 75580 94706 75620
rect 94750 75580 94790 75620
rect 94790 75580 94830 75620
rect 94830 75580 94872 75620
rect 94872 75580 94874 75620
rect 94582 75538 94706 75580
rect 94750 75538 94874 75580
rect 109702 75620 109826 75662
rect 109870 75620 109994 75662
rect 109702 75580 109704 75620
rect 109704 75580 109746 75620
rect 109746 75580 109786 75620
rect 109786 75580 109826 75620
rect 109870 75580 109910 75620
rect 109910 75580 109950 75620
rect 109950 75580 109992 75620
rect 109992 75580 109994 75620
rect 109702 75538 109826 75580
rect 109870 75538 109994 75580
rect 124822 75620 124946 75662
rect 124990 75620 125114 75662
rect 124822 75580 124824 75620
rect 124824 75580 124866 75620
rect 124866 75580 124906 75620
rect 124906 75580 124946 75620
rect 124990 75580 125030 75620
rect 125030 75580 125070 75620
rect 125070 75580 125112 75620
rect 125112 75580 125114 75620
rect 124822 75538 124946 75580
rect 124990 75538 125114 75580
rect 139942 75620 140066 75662
rect 140110 75620 140234 75662
rect 139942 75580 139944 75620
rect 139944 75580 139986 75620
rect 139986 75580 140026 75620
rect 140026 75580 140066 75620
rect 140110 75580 140150 75620
rect 140150 75580 140190 75620
rect 140190 75580 140232 75620
rect 140232 75580 140234 75620
rect 139942 75538 140066 75580
rect 140110 75538 140234 75580
<< metal6 >>
rect 67748 155942 70748 156076
rect 67748 155562 67882 155942
rect 68262 155562 68274 155942
rect 68654 155562 68666 155942
rect 69046 155562 69058 155942
rect 69438 155562 69450 155942
rect 69830 155562 69842 155942
rect 70222 155562 70234 155942
rect 70614 155562 70748 155942
rect 67748 155550 70748 155562
rect 67748 155170 67882 155550
rect 68262 155170 68274 155550
rect 68654 155170 68666 155550
rect 69046 155170 69058 155550
rect 69438 155170 69450 155550
rect 69830 155170 69842 155550
rect 70222 155170 70234 155550
rect 70614 155170 70748 155550
rect 67748 155158 70748 155170
rect 67748 154778 67882 155158
rect 68262 154778 68274 155158
rect 68654 154778 68666 155158
rect 69046 154778 69058 155158
rect 69438 154778 69450 155158
rect 69830 154778 69842 155158
rect 70222 154778 70234 155158
rect 70614 154778 70748 155158
rect 67748 154766 70748 154778
rect 67748 154386 67882 154766
rect 68262 154386 68274 154766
rect 68654 154386 68666 154766
rect 69046 154386 69058 154766
rect 69438 154386 69450 154766
rect 69830 154386 69842 154766
rect 70222 154386 70234 154766
rect 70614 154386 70748 154766
rect 67748 154374 70748 154386
rect 67748 153994 67882 154374
rect 68262 153994 68274 154374
rect 68654 153994 68666 154374
rect 69046 153994 69058 154374
rect 69438 153994 69450 154374
rect 69830 153994 69842 154374
rect 70222 153994 70234 154374
rect 70614 153994 70748 154374
rect 67748 153982 70748 153994
rect 67748 153602 67882 153982
rect 68262 153602 68274 153982
rect 68654 153602 68666 153982
rect 69046 153602 69058 153982
rect 69438 153602 69450 153982
rect 69830 153602 69842 153982
rect 70222 153602 70234 153982
rect 70614 153602 70748 153982
rect 67748 153590 70748 153602
rect 67748 153210 67882 153590
rect 68262 153210 68274 153590
rect 68654 153210 68666 153590
rect 69046 153210 69058 153590
rect 69438 153210 69450 153590
rect 69830 153210 69842 153590
rect 70222 153210 70234 153590
rect 70614 153210 70748 153590
rect 67748 140230 70748 153210
rect 79388 155942 79828 156076
rect 79388 155562 79418 155942
rect 79798 155562 79828 155942
rect 79388 155550 79828 155562
rect 79388 155170 79418 155550
rect 79798 155170 79828 155550
rect 79388 155158 79828 155170
rect 79388 154778 79418 155158
rect 79798 154778 79828 155158
rect 79388 154766 79828 154778
rect 79388 154386 79418 154766
rect 79798 154386 79828 154766
rect 79388 154374 79828 154386
rect 79388 153994 79418 154374
rect 79798 153994 79828 154374
rect 79388 153982 79828 153994
rect 79388 153602 79418 153982
rect 79798 153602 79828 153982
rect 79388 153590 79828 153602
rect 79388 153210 79418 153590
rect 79798 153210 79828 153590
rect 67748 139850 67882 140230
rect 68262 139850 68274 140230
rect 68654 139850 68666 140230
rect 69046 139850 69058 140230
rect 69438 139850 69450 140230
rect 69830 139850 69842 140230
rect 70222 139850 70234 140230
rect 70614 139850 70748 140230
rect 56000 133169 59600 133332
rect 56000 132789 56042 133169
rect 56422 132789 56434 133169
rect 56814 132789 56826 133169
rect 57206 132789 57218 133169
rect 57598 132789 57610 133169
rect 57990 132789 58002 133169
rect 58382 132789 58394 133169
rect 58774 132789 58786 133169
rect 59166 132789 59178 133169
rect 59558 132789 59600 133169
rect 56000 132777 59600 132789
rect 56000 132397 56042 132777
rect 56422 132397 56434 132777
rect 56814 132397 56826 132777
rect 57206 132397 57218 132777
rect 57598 132397 57610 132777
rect 57990 132397 58002 132777
rect 58382 132397 58394 132777
rect 58774 132397 58786 132777
rect 59166 132397 59178 132777
rect 59558 132397 59600 132777
rect 56000 132385 59600 132397
rect 56000 132005 56042 132385
rect 56422 132005 56434 132385
rect 56814 132005 56826 132385
rect 57206 132005 57218 132385
rect 57598 132005 57610 132385
rect 57990 132005 58002 132385
rect 58382 132005 58394 132385
rect 58774 132005 58786 132385
rect 59166 132005 59178 132385
rect 59558 132005 59600 132385
rect 56000 131993 59600 132005
rect 56000 131613 56042 131993
rect 56422 131613 56434 131993
rect 56814 131613 56826 131993
rect 57206 131613 57218 131993
rect 57598 131613 57610 131993
rect 57990 131613 58002 131993
rect 58382 131613 58394 131993
rect 58774 131613 58786 131993
rect 59166 131613 59178 131993
rect 59558 131613 59600 131993
rect 56000 131601 59600 131613
rect 56000 131221 56042 131601
rect 56422 131221 56434 131601
rect 56814 131221 56826 131601
rect 57206 131221 57218 131601
rect 57598 131221 57610 131601
rect 57990 131221 58002 131601
rect 58382 131221 58394 131601
rect 58774 131221 58786 131601
rect 59166 131221 59178 131601
rect 59558 131221 59600 131601
rect 56000 131209 59600 131221
rect 56000 130829 56042 131209
rect 56422 130829 56434 131209
rect 56814 130829 56826 131209
rect 57206 130829 57218 131209
rect 57598 130829 57610 131209
rect 57990 130829 58002 131209
rect 58382 130829 58394 131209
rect 58774 130829 58786 131209
rect 59166 130829 59178 131209
rect 59558 130829 59600 131209
rect 56000 130666 59600 130829
rect 67748 125110 70748 139850
rect 67748 124730 67882 125110
rect 68262 124730 68274 125110
rect 68654 124730 68666 125110
rect 69046 124730 69058 125110
rect 69438 124730 69450 125110
rect 69830 124730 69842 125110
rect 70222 124730 70234 125110
rect 70614 124730 70748 125110
rect 56000 117169 59600 117332
rect 56000 116789 56042 117169
rect 56422 116789 56434 117169
rect 56814 116789 56826 117169
rect 57206 116789 57218 117169
rect 57598 116789 57610 117169
rect 57990 116789 58002 117169
rect 58382 116789 58394 117169
rect 58774 116789 58786 117169
rect 59166 116789 59178 117169
rect 59558 116789 59600 117169
rect 56000 116777 59600 116789
rect 56000 116397 56042 116777
rect 56422 116397 56434 116777
rect 56814 116397 56826 116777
rect 57206 116397 57218 116777
rect 57598 116397 57610 116777
rect 57990 116397 58002 116777
rect 58382 116397 58394 116777
rect 58774 116397 58786 116777
rect 59166 116397 59178 116777
rect 59558 116397 59600 116777
rect 56000 116385 59600 116397
rect 56000 116005 56042 116385
rect 56422 116005 56434 116385
rect 56814 116005 56826 116385
rect 57206 116005 57218 116385
rect 57598 116005 57610 116385
rect 57990 116005 58002 116385
rect 58382 116005 58394 116385
rect 58774 116005 58786 116385
rect 59166 116005 59178 116385
rect 59558 116005 59600 116385
rect 56000 115993 59600 116005
rect 56000 115613 56042 115993
rect 56422 115613 56434 115993
rect 56814 115613 56826 115993
rect 57206 115613 57218 115993
rect 57598 115613 57610 115993
rect 57990 115613 58002 115993
rect 58382 115613 58394 115993
rect 58774 115613 58786 115993
rect 59166 115613 59178 115993
rect 59558 115613 59600 115993
rect 56000 115601 59600 115613
rect 56000 115221 56042 115601
rect 56422 115221 56434 115601
rect 56814 115221 56826 115601
rect 57206 115221 57218 115601
rect 57598 115221 57610 115601
rect 57990 115221 58002 115601
rect 58382 115221 58394 115601
rect 58774 115221 58786 115601
rect 59166 115221 59178 115601
rect 59558 115221 59600 115601
rect 56000 115209 59600 115221
rect 56000 114829 56042 115209
rect 56422 114829 56434 115209
rect 56814 114829 56826 115209
rect 57206 114829 57218 115209
rect 57598 114829 57610 115209
rect 57990 114829 58002 115209
rect 58382 114829 58394 115209
rect 58774 114829 58786 115209
rect 59166 114829 59178 115209
rect 59558 114829 59600 115209
rect 56000 114666 59600 114829
rect 67748 109990 70748 124730
rect 67748 109610 67882 109990
rect 68262 109610 68274 109990
rect 68654 109610 68666 109990
rect 69046 109610 69058 109990
rect 69438 109610 69450 109990
rect 69830 109610 69842 109990
rect 70222 109610 70234 109990
rect 70614 109610 70748 109990
rect 60000 106501 63600 106664
rect 60000 106121 60042 106501
rect 60422 106121 60434 106501
rect 60814 106121 60826 106501
rect 61206 106121 61218 106501
rect 61598 106121 61610 106501
rect 61990 106121 62002 106501
rect 62382 106121 62394 106501
rect 62774 106121 62786 106501
rect 63166 106121 63178 106501
rect 63558 106121 63600 106501
rect 60000 106109 63600 106121
rect 60000 105729 60042 106109
rect 60422 105729 60434 106109
rect 60814 105729 60826 106109
rect 61206 105729 61218 106109
rect 61598 105729 61610 106109
rect 61990 105729 62002 106109
rect 62382 105729 62394 106109
rect 62774 105729 62786 106109
rect 63166 105729 63178 106109
rect 63558 105729 63600 106109
rect 60000 105717 63600 105729
rect 60000 105337 60042 105717
rect 60422 105337 60434 105717
rect 60814 105337 60826 105717
rect 61206 105337 61218 105717
rect 61598 105337 61610 105717
rect 61990 105337 62002 105717
rect 62382 105337 62394 105717
rect 62774 105337 62786 105717
rect 63166 105337 63178 105717
rect 63558 105337 63600 105717
rect 60000 105325 63600 105337
rect 60000 104945 60042 105325
rect 60422 104945 60434 105325
rect 60814 104945 60826 105325
rect 61206 104945 61218 105325
rect 61598 104945 61610 105325
rect 61990 104945 62002 105325
rect 62382 104945 62394 105325
rect 62774 104945 62786 105325
rect 63166 104945 63178 105325
rect 63558 104945 63600 105325
rect 60000 104933 63600 104945
rect 60000 104553 60042 104933
rect 60422 104553 60434 104933
rect 60814 104553 60826 104933
rect 61206 104553 61218 104933
rect 61598 104553 61610 104933
rect 61990 104553 62002 104933
rect 62382 104553 62394 104933
rect 62774 104553 62786 104933
rect 63166 104553 63178 104933
rect 63558 104553 63600 104933
rect 60000 104541 63600 104553
rect 60000 104161 60042 104541
rect 60422 104161 60434 104541
rect 60814 104161 60826 104541
rect 61206 104161 61218 104541
rect 61598 104161 61610 104541
rect 61990 104161 62002 104541
rect 62382 104161 62394 104541
rect 62774 104161 62786 104541
rect 63166 104161 63178 104541
rect 63558 104161 63600 104541
rect 60000 103998 63600 104161
rect 67748 106501 70748 109610
rect 67748 106121 67882 106501
rect 68262 106121 68274 106501
rect 68654 106121 68666 106501
rect 69046 106121 69058 106501
rect 69438 106121 69450 106501
rect 69830 106121 69842 106501
rect 70222 106121 70234 106501
rect 70614 106121 70748 106501
rect 67748 106109 70748 106121
rect 67748 105729 67882 106109
rect 68262 105729 68274 106109
rect 68654 105729 68666 106109
rect 69046 105729 69058 106109
rect 69438 105729 69450 106109
rect 69830 105729 69842 106109
rect 70222 105729 70234 106109
rect 70614 105729 70748 106109
rect 67748 105717 70748 105729
rect 67748 105337 67882 105717
rect 68262 105337 68274 105717
rect 68654 105337 68666 105717
rect 69046 105337 69058 105717
rect 69438 105337 69450 105717
rect 69830 105337 69842 105717
rect 70222 105337 70234 105717
rect 70614 105337 70748 105717
rect 67748 105325 70748 105337
rect 67748 104945 67882 105325
rect 68262 104945 68274 105325
rect 68654 104945 68666 105325
rect 69046 104945 69058 105325
rect 69438 104945 69450 105325
rect 69830 104945 69842 105325
rect 70222 104945 70234 105325
rect 70614 104945 70748 105325
rect 67748 104933 70748 104945
rect 67748 104553 67882 104933
rect 68262 104553 68274 104933
rect 68654 104553 68666 104933
rect 69046 104553 69058 104933
rect 69438 104553 69450 104933
rect 69830 104553 69842 104933
rect 70222 104553 70234 104933
rect 70614 104553 70748 104933
rect 67748 104541 70748 104553
rect 67748 104161 67882 104541
rect 68262 104161 68274 104541
rect 68654 104161 68666 104541
rect 69046 104161 69058 104541
rect 69438 104161 69450 104541
rect 69830 104161 69842 104541
rect 70222 104161 70234 104541
rect 70614 104161 70748 104541
rect 56000 101169 59600 101332
rect 56000 100789 56042 101169
rect 56422 100789 56434 101169
rect 56814 100789 56826 101169
rect 57206 100789 57218 101169
rect 57598 100789 57610 101169
rect 57990 100789 58002 101169
rect 58382 100789 58394 101169
rect 58774 100789 58786 101169
rect 59166 100789 59178 101169
rect 59558 100789 59600 101169
rect 56000 100777 59600 100789
rect 56000 100397 56042 100777
rect 56422 100397 56434 100777
rect 56814 100397 56826 100777
rect 57206 100397 57218 100777
rect 57598 100397 57610 100777
rect 57990 100397 58002 100777
rect 58382 100397 58394 100777
rect 58774 100397 58786 100777
rect 59166 100397 59178 100777
rect 59558 100397 59600 100777
rect 56000 100385 59600 100397
rect 56000 100005 56042 100385
rect 56422 100005 56434 100385
rect 56814 100005 56826 100385
rect 57206 100005 57218 100385
rect 57598 100005 57610 100385
rect 57990 100005 58002 100385
rect 58382 100005 58394 100385
rect 58774 100005 58786 100385
rect 59166 100005 59178 100385
rect 59558 100005 59600 100385
rect 56000 99993 59600 100005
rect 56000 99613 56042 99993
rect 56422 99613 56434 99993
rect 56814 99613 56826 99993
rect 57206 99613 57218 99993
rect 57598 99613 57610 99993
rect 57990 99613 58002 99993
rect 58382 99613 58394 99993
rect 58774 99613 58786 99993
rect 59166 99613 59178 99993
rect 59558 99613 59600 99993
rect 56000 99601 59600 99613
rect 56000 99221 56042 99601
rect 56422 99221 56434 99601
rect 56814 99221 56826 99601
rect 57206 99221 57218 99601
rect 57598 99221 57610 99601
rect 57990 99221 58002 99601
rect 58382 99221 58394 99601
rect 58774 99221 58786 99601
rect 59166 99221 59178 99601
rect 59558 99221 59600 99601
rect 56000 99209 59600 99221
rect 56000 98829 56042 99209
rect 56422 98829 56434 99209
rect 56814 98829 56826 99209
rect 57206 98829 57218 99209
rect 57598 98829 57610 99209
rect 57990 98829 58002 99209
rect 58382 98829 58394 99209
rect 58774 98829 58786 99209
rect 59166 98829 59178 99209
rect 59558 98829 59600 99209
rect 56000 98666 59600 98829
rect 67748 94870 70748 104161
rect 67748 94490 67882 94870
rect 68262 94490 68274 94870
rect 68654 94490 68666 94870
rect 69046 94490 69058 94870
rect 69438 94490 69450 94870
rect 69830 94490 69842 94870
rect 70222 94490 70234 94870
rect 70614 94490 70748 94870
rect 60000 90501 63600 90664
rect 60000 90121 60042 90501
rect 60422 90121 60434 90501
rect 60814 90121 60826 90501
rect 61206 90121 61218 90501
rect 61598 90121 61610 90501
rect 61990 90121 62002 90501
rect 62382 90121 62394 90501
rect 62774 90121 62786 90501
rect 63166 90121 63178 90501
rect 63558 90121 63600 90501
rect 60000 90109 63600 90121
rect 60000 89729 60042 90109
rect 60422 89729 60434 90109
rect 60814 89729 60826 90109
rect 61206 89729 61218 90109
rect 61598 89729 61610 90109
rect 61990 89729 62002 90109
rect 62382 89729 62394 90109
rect 62774 89729 62786 90109
rect 63166 89729 63178 90109
rect 63558 89729 63600 90109
rect 60000 89717 63600 89729
rect 60000 89337 60042 89717
rect 60422 89337 60434 89717
rect 60814 89337 60826 89717
rect 61206 89337 61218 89717
rect 61598 89337 61610 89717
rect 61990 89337 62002 89717
rect 62382 89337 62394 89717
rect 62774 89337 62786 89717
rect 63166 89337 63178 89717
rect 63558 89337 63600 89717
rect 60000 89325 63600 89337
rect 60000 88945 60042 89325
rect 60422 88945 60434 89325
rect 60814 88945 60826 89325
rect 61206 88945 61218 89325
rect 61598 88945 61610 89325
rect 61990 88945 62002 89325
rect 62382 88945 62394 89325
rect 62774 88945 62786 89325
rect 63166 88945 63178 89325
rect 63558 88945 63600 89325
rect 60000 88933 63600 88945
rect 60000 88553 60042 88933
rect 60422 88553 60434 88933
rect 60814 88553 60826 88933
rect 61206 88553 61218 88933
rect 61598 88553 61610 88933
rect 61990 88553 62002 88933
rect 62382 88553 62394 88933
rect 62774 88553 62786 88933
rect 63166 88553 63178 88933
rect 63558 88553 63600 88933
rect 60000 88541 63600 88553
rect 60000 88161 60042 88541
rect 60422 88161 60434 88541
rect 60814 88161 60826 88541
rect 61206 88161 61218 88541
rect 61598 88161 61610 88541
rect 61990 88161 62002 88541
rect 62382 88161 62394 88541
rect 62774 88161 62786 88541
rect 63166 88161 63178 88541
rect 63558 88161 63600 88541
rect 60000 87998 63600 88161
rect 67748 90501 70748 94490
rect 67748 90121 67882 90501
rect 68262 90121 68274 90501
rect 68654 90121 68666 90501
rect 69046 90121 69058 90501
rect 69438 90121 69450 90501
rect 69830 90121 69842 90501
rect 70222 90121 70234 90501
rect 70614 90121 70748 90501
rect 67748 90109 70748 90121
rect 67748 89729 67882 90109
rect 68262 89729 68274 90109
rect 68654 89729 68666 90109
rect 69046 89729 69058 90109
rect 69438 89729 69450 90109
rect 69830 89729 69842 90109
rect 70222 89729 70234 90109
rect 70614 89729 70748 90109
rect 67748 89717 70748 89729
rect 67748 89337 67882 89717
rect 68262 89337 68274 89717
rect 68654 89337 68666 89717
rect 69046 89337 69058 89717
rect 69438 89337 69450 89717
rect 69830 89337 69842 89717
rect 70222 89337 70234 89717
rect 70614 89337 70748 89717
rect 67748 89325 70748 89337
rect 67748 88945 67882 89325
rect 68262 88945 68274 89325
rect 68654 88945 68666 89325
rect 69046 88945 69058 89325
rect 69438 88945 69450 89325
rect 69830 88945 69842 89325
rect 70222 88945 70234 89325
rect 70614 88945 70748 89325
rect 67748 88933 70748 88945
rect 67748 88553 67882 88933
rect 68262 88553 68274 88933
rect 68654 88553 68666 88933
rect 69046 88553 69058 88933
rect 69438 88553 69450 88933
rect 69830 88553 69842 88933
rect 70222 88553 70234 88933
rect 70614 88553 70748 88933
rect 67748 88541 70748 88553
rect 67748 88161 67882 88541
rect 68262 88161 68274 88541
rect 68654 88161 68666 88541
rect 69046 88161 69058 88541
rect 69438 88161 69450 88541
rect 69830 88161 69842 88541
rect 70222 88161 70234 88541
rect 70614 88161 70748 88541
rect 56000 85169 59600 85332
rect 56000 84789 56042 85169
rect 56422 84789 56434 85169
rect 56814 84789 56826 85169
rect 57206 84789 57218 85169
rect 57598 84789 57610 85169
rect 57990 84789 58002 85169
rect 58382 84789 58394 85169
rect 58774 84789 58786 85169
rect 59166 84789 59178 85169
rect 59558 84789 59600 85169
rect 56000 84777 59600 84789
rect 56000 84397 56042 84777
rect 56422 84397 56434 84777
rect 56814 84397 56826 84777
rect 57206 84397 57218 84777
rect 57598 84397 57610 84777
rect 57990 84397 58002 84777
rect 58382 84397 58394 84777
rect 58774 84397 58786 84777
rect 59166 84397 59178 84777
rect 59558 84397 59600 84777
rect 56000 84385 59600 84397
rect 56000 84005 56042 84385
rect 56422 84005 56434 84385
rect 56814 84005 56826 84385
rect 57206 84005 57218 84385
rect 57598 84005 57610 84385
rect 57990 84005 58002 84385
rect 58382 84005 58394 84385
rect 58774 84005 58786 84385
rect 59166 84005 59178 84385
rect 59558 84005 59600 84385
rect 56000 83993 59600 84005
rect 56000 83613 56042 83993
rect 56422 83613 56434 83993
rect 56814 83613 56826 83993
rect 57206 83613 57218 83993
rect 57598 83613 57610 83993
rect 57990 83613 58002 83993
rect 58382 83613 58394 83993
rect 58774 83613 58786 83993
rect 59166 83613 59178 83993
rect 59558 83613 59600 83993
rect 56000 83601 59600 83613
rect 56000 83221 56042 83601
rect 56422 83221 56434 83601
rect 56814 83221 56826 83601
rect 57206 83221 57218 83601
rect 57598 83221 57610 83601
rect 57990 83221 58002 83601
rect 58382 83221 58394 83601
rect 58774 83221 58786 83601
rect 59166 83221 59178 83601
rect 59558 83221 59600 83601
rect 56000 83209 59600 83221
rect 56000 82829 56042 83209
rect 56422 82829 56434 83209
rect 56814 82829 56826 83209
rect 57206 82829 57218 83209
rect 57598 82829 57610 83209
rect 57990 82829 58002 83209
rect 58382 82829 58394 83209
rect 58774 82829 58786 83209
rect 59166 82829 59178 83209
rect 59558 82829 59600 83209
rect 56000 82666 59600 82829
rect 67748 79750 70748 88161
rect 67748 79370 67882 79750
rect 68262 79370 68274 79750
rect 68654 79370 68666 79750
rect 69046 79370 69058 79750
rect 69438 79370 69450 79750
rect 69830 79370 69842 79750
rect 70222 79370 70234 79750
rect 70614 79370 70748 79750
rect 60000 74501 63600 74664
rect 60000 74121 60042 74501
rect 60422 74121 60434 74501
rect 60814 74121 60826 74501
rect 61206 74121 61218 74501
rect 61598 74121 61610 74501
rect 61990 74121 62002 74501
rect 62382 74121 62394 74501
rect 62774 74121 62786 74501
rect 63166 74121 63178 74501
rect 63558 74121 63600 74501
rect 60000 74109 63600 74121
rect 60000 73729 60042 74109
rect 60422 73729 60434 74109
rect 60814 73729 60826 74109
rect 61206 73729 61218 74109
rect 61598 73729 61610 74109
rect 61990 73729 62002 74109
rect 62382 73729 62394 74109
rect 62774 73729 62786 74109
rect 63166 73729 63178 74109
rect 63558 73729 63600 74109
rect 60000 73717 63600 73729
rect 60000 73337 60042 73717
rect 60422 73337 60434 73717
rect 60814 73337 60826 73717
rect 61206 73337 61218 73717
rect 61598 73337 61610 73717
rect 61990 73337 62002 73717
rect 62382 73337 62394 73717
rect 62774 73337 62786 73717
rect 63166 73337 63178 73717
rect 63558 73337 63600 73717
rect 60000 73325 63600 73337
rect 60000 72945 60042 73325
rect 60422 72945 60434 73325
rect 60814 72945 60826 73325
rect 61206 72945 61218 73325
rect 61598 72945 61610 73325
rect 61990 72945 62002 73325
rect 62382 72945 62394 73325
rect 62774 72945 62786 73325
rect 63166 72945 63178 73325
rect 63558 72945 63600 73325
rect 60000 72933 63600 72945
rect 60000 72553 60042 72933
rect 60422 72553 60434 72933
rect 60814 72553 60826 72933
rect 61206 72553 61218 72933
rect 61598 72553 61610 72933
rect 61990 72553 62002 72933
rect 62382 72553 62394 72933
rect 62774 72553 62786 72933
rect 63166 72553 63178 72933
rect 63558 72553 63600 72933
rect 60000 72541 63600 72553
rect 60000 72161 60042 72541
rect 60422 72161 60434 72541
rect 60814 72161 60826 72541
rect 61206 72161 61218 72541
rect 61598 72161 61610 72541
rect 61990 72161 62002 72541
rect 62382 72161 62394 72541
rect 62774 72161 62786 72541
rect 63166 72161 63178 72541
rect 63558 72161 63600 72541
rect 60000 71998 63600 72161
rect 67748 74501 70748 79370
rect 67748 74121 67882 74501
rect 68262 74121 68274 74501
rect 68654 74121 68666 74501
rect 69046 74121 69058 74501
rect 69438 74121 69450 74501
rect 69830 74121 69842 74501
rect 70222 74121 70234 74501
rect 70614 74121 70748 74501
rect 67748 74109 70748 74121
rect 67748 73729 67882 74109
rect 68262 73729 68274 74109
rect 68654 73729 68666 74109
rect 69046 73729 69058 74109
rect 69438 73729 69450 74109
rect 69830 73729 69842 74109
rect 70222 73729 70234 74109
rect 70614 73729 70748 74109
rect 67748 73717 70748 73729
rect 67748 73337 67882 73717
rect 68262 73337 68274 73717
rect 68654 73337 68666 73717
rect 69046 73337 69058 73717
rect 69438 73337 69450 73717
rect 69830 73337 69842 73717
rect 70222 73337 70234 73717
rect 70614 73337 70748 73717
rect 67748 73325 70748 73337
rect 67748 72945 67882 73325
rect 68262 72945 68274 73325
rect 68654 72945 68666 73325
rect 69046 72945 69058 73325
rect 69438 72945 69450 73325
rect 69830 72945 69842 73325
rect 70222 72945 70234 73325
rect 70614 72945 70748 73325
rect 67748 72933 70748 72945
rect 67748 72553 67882 72933
rect 68262 72553 68274 72933
rect 68654 72553 68666 72933
rect 69046 72553 69058 72933
rect 69438 72553 69450 72933
rect 69830 72553 69842 72933
rect 70222 72553 70234 72933
rect 70614 72553 70748 72933
rect 67748 72541 70748 72553
rect 67748 72161 67882 72541
rect 68262 72161 68274 72541
rect 68654 72161 68666 72541
rect 69046 72161 69058 72541
rect 69438 72161 69450 72541
rect 69830 72161 69842 72541
rect 70222 72161 70234 72541
rect 70614 72161 70748 72541
rect 67748 70566 70748 72161
rect 71748 151942 74748 152076
rect 71748 151562 71882 151942
rect 72262 151562 72274 151942
rect 72654 151562 72666 151942
rect 73046 151562 73058 151942
rect 73438 151562 73450 151942
rect 73830 151562 73842 151942
rect 74222 151562 74234 151942
rect 74614 151562 74748 151942
rect 71748 151550 74748 151562
rect 71748 151170 71882 151550
rect 72262 151170 72274 151550
rect 72654 151170 72666 151550
rect 73046 151170 73058 151550
rect 73438 151170 73450 151550
rect 73830 151170 73842 151550
rect 74222 151170 74234 151550
rect 74614 151170 74748 151550
rect 71748 151158 74748 151170
rect 71748 150778 71882 151158
rect 72262 150778 72274 151158
rect 72654 150778 72666 151158
rect 73046 150778 73058 151158
rect 73438 150778 73450 151158
rect 73830 150778 73842 151158
rect 74222 150778 74234 151158
rect 74614 150778 74748 151158
rect 71748 150766 74748 150778
rect 71748 150386 71882 150766
rect 72262 150386 72274 150766
rect 72654 150386 72666 150766
rect 73046 150386 73058 150766
rect 73438 150386 73450 150766
rect 73830 150386 73842 150766
rect 74222 150386 74234 150766
rect 74614 150386 74748 150766
rect 71748 150374 74748 150386
rect 71748 149994 71882 150374
rect 72262 149994 72274 150374
rect 72654 149994 72666 150374
rect 73046 149994 73058 150374
rect 73438 149994 73450 150374
rect 73830 149994 73842 150374
rect 74222 149994 74234 150374
rect 74614 149994 74748 150374
rect 71748 149982 74748 149994
rect 71748 149602 71882 149982
rect 72262 149602 72274 149982
rect 72654 149602 72666 149982
rect 73046 149602 73058 149982
rect 73438 149602 73450 149982
rect 73830 149602 73842 149982
rect 74222 149602 74234 149982
rect 74614 149602 74748 149982
rect 71748 149590 74748 149602
rect 71748 149210 71882 149590
rect 72262 149210 72274 149590
rect 72654 149210 72666 149590
rect 73046 149210 73058 149590
rect 73438 149210 73450 149590
rect 73830 149210 73842 149590
rect 74222 149210 74234 149590
rect 74614 149210 74748 149590
rect 71748 138990 74748 149210
rect 71748 138610 71882 138990
rect 72262 138610 72274 138990
rect 72654 138610 72666 138990
rect 73046 138610 73058 138990
rect 73438 138610 73450 138990
rect 73830 138610 73842 138990
rect 74222 138610 74234 138990
rect 74614 138610 74748 138990
rect 71748 133169 74748 138610
rect 71748 132789 71882 133169
rect 72262 132789 72274 133169
rect 72654 132789 72666 133169
rect 73046 132789 73058 133169
rect 73438 132789 73450 133169
rect 73830 132789 73842 133169
rect 74222 132789 74234 133169
rect 74614 132789 74748 133169
rect 71748 132777 74748 132789
rect 71748 132397 71882 132777
rect 72262 132397 72274 132777
rect 72654 132397 72666 132777
rect 73046 132397 73058 132777
rect 73438 132397 73450 132777
rect 73830 132397 73842 132777
rect 74222 132397 74234 132777
rect 74614 132397 74748 132777
rect 71748 132385 74748 132397
rect 71748 132005 71882 132385
rect 72262 132005 72274 132385
rect 72654 132005 72666 132385
rect 73046 132005 73058 132385
rect 73438 132005 73450 132385
rect 73830 132005 73842 132385
rect 74222 132005 74234 132385
rect 74614 132005 74748 132385
rect 71748 131993 74748 132005
rect 71748 131613 71882 131993
rect 72262 131613 72274 131993
rect 72654 131613 72666 131993
rect 73046 131613 73058 131993
rect 73438 131613 73450 131993
rect 73830 131613 73842 131993
rect 74222 131613 74234 131993
rect 74614 131613 74748 131993
rect 71748 131601 74748 131613
rect 71748 131221 71882 131601
rect 72262 131221 72274 131601
rect 72654 131221 72666 131601
rect 73046 131221 73058 131601
rect 73438 131221 73450 131601
rect 73830 131221 73842 131601
rect 74222 131221 74234 131601
rect 74614 131221 74748 131601
rect 71748 131209 74748 131221
rect 71748 130829 71882 131209
rect 72262 130829 72274 131209
rect 72654 130829 72666 131209
rect 73046 130829 73058 131209
rect 73438 130829 73450 131209
rect 73830 130829 73842 131209
rect 74222 130829 74234 131209
rect 74614 130829 74748 131209
rect 71748 123870 74748 130829
rect 71748 123490 71882 123870
rect 72262 123490 72274 123870
rect 72654 123490 72666 123870
rect 73046 123490 73058 123870
rect 73438 123490 73450 123870
rect 73830 123490 73842 123870
rect 74222 123490 74234 123870
rect 74614 123490 74748 123870
rect 71748 117169 74748 123490
rect 71748 116789 71882 117169
rect 72262 116789 72274 117169
rect 72654 116789 72666 117169
rect 73046 116789 73058 117169
rect 73438 116789 73450 117169
rect 73830 116789 73842 117169
rect 74222 116789 74234 117169
rect 74614 116789 74748 117169
rect 71748 116777 74748 116789
rect 71748 116397 71882 116777
rect 72262 116397 72274 116777
rect 72654 116397 72666 116777
rect 73046 116397 73058 116777
rect 73438 116397 73450 116777
rect 73830 116397 73842 116777
rect 74222 116397 74234 116777
rect 74614 116397 74748 116777
rect 71748 116385 74748 116397
rect 71748 116005 71882 116385
rect 72262 116005 72274 116385
rect 72654 116005 72666 116385
rect 73046 116005 73058 116385
rect 73438 116005 73450 116385
rect 73830 116005 73842 116385
rect 74222 116005 74234 116385
rect 74614 116005 74748 116385
rect 71748 115993 74748 116005
rect 71748 115613 71882 115993
rect 72262 115613 72274 115993
rect 72654 115613 72666 115993
rect 73046 115613 73058 115993
rect 73438 115613 73450 115993
rect 73830 115613 73842 115993
rect 74222 115613 74234 115993
rect 74614 115613 74748 115993
rect 71748 115601 74748 115613
rect 71748 115221 71882 115601
rect 72262 115221 72274 115601
rect 72654 115221 72666 115601
rect 73046 115221 73058 115601
rect 73438 115221 73450 115601
rect 73830 115221 73842 115601
rect 74222 115221 74234 115601
rect 74614 115221 74748 115601
rect 71748 115209 74748 115221
rect 71748 114829 71882 115209
rect 72262 114829 72274 115209
rect 72654 114829 72666 115209
rect 73046 114829 73058 115209
rect 73438 114829 73450 115209
rect 73830 114829 73842 115209
rect 74222 114829 74234 115209
rect 74614 114829 74748 115209
rect 71748 108750 74748 114829
rect 71748 108370 71882 108750
rect 72262 108370 72274 108750
rect 72654 108370 72666 108750
rect 73046 108370 73058 108750
rect 73438 108370 73450 108750
rect 73830 108370 73842 108750
rect 74222 108370 74234 108750
rect 74614 108370 74748 108750
rect 71748 101169 74748 108370
rect 71748 100789 71882 101169
rect 72262 100789 72274 101169
rect 72654 100789 72666 101169
rect 73046 100789 73058 101169
rect 73438 100789 73450 101169
rect 73830 100789 73842 101169
rect 74222 100789 74234 101169
rect 74614 100789 74748 101169
rect 71748 100777 74748 100789
rect 71748 100397 71882 100777
rect 72262 100397 72274 100777
rect 72654 100397 72666 100777
rect 73046 100397 73058 100777
rect 73438 100397 73450 100777
rect 73830 100397 73842 100777
rect 74222 100397 74234 100777
rect 74614 100397 74748 100777
rect 71748 100385 74748 100397
rect 71748 100005 71882 100385
rect 72262 100005 72274 100385
rect 72654 100005 72666 100385
rect 73046 100005 73058 100385
rect 73438 100005 73450 100385
rect 73830 100005 73842 100385
rect 74222 100005 74234 100385
rect 74614 100005 74748 100385
rect 71748 99993 74748 100005
rect 71748 99613 71882 99993
rect 72262 99613 72274 99993
rect 72654 99613 72666 99993
rect 73046 99613 73058 99993
rect 73438 99613 73450 99993
rect 73830 99613 73842 99993
rect 74222 99613 74234 99993
rect 74614 99613 74748 99993
rect 71748 99601 74748 99613
rect 71748 99221 71882 99601
rect 72262 99221 72274 99601
rect 72654 99221 72666 99601
rect 73046 99221 73058 99601
rect 73438 99221 73450 99601
rect 73830 99221 73842 99601
rect 74222 99221 74234 99601
rect 74614 99221 74748 99601
rect 71748 99209 74748 99221
rect 71748 98829 71882 99209
rect 72262 98829 72274 99209
rect 72654 98829 72666 99209
rect 73046 98829 73058 99209
rect 73438 98829 73450 99209
rect 73830 98829 73842 99209
rect 74222 98829 74234 99209
rect 74614 98829 74748 99209
rect 71748 93630 74748 98829
rect 71748 93250 71882 93630
rect 72262 93250 72274 93630
rect 72654 93250 72666 93630
rect 73046 93250 73058 93630
rect 73438 93250 73450 93630
rect 73830 93250 73842 93630
rect 74222 93250 74234 93630
rect 74614 93250 74748 93630
rect 71748 85169 74748 93250
rect 71748 84789 71882 85169
rect 72262 84789 72274 85169
rect 72654 84789 72666 85169
rect 73046 84789 73058 85169
rect 73438 84789 73450 85169
rect 73830 84789 73842 85169
rect 74222 84789 74234 85169
rect 74614 84789 74748 85169
rect 71748 84777 74748 84789
rect 71748 84397 71882 84777
rect 72262 84397 72274 84777
rect 72654 84397 72666 84777
rect 73046 84397 73058 84777
rect 73438 84397 73450 84777
rect 73830 84397 73842 84777
rect 74222 84397 74234 84777
rect 74614 84397 74748 84777
rect 71748 84385 74748 84397
rect 71748 84005 71882 84385
rect 72262 84005 72274 84385
rect 72654 84005 72666 84385
rect 73046 84005 73058 84385
rect 73438 84005 73450 84385
rect 73830 84005 73842 84385
rect 74222 84005 74234 84385
rect 74614 84005 74748 84385
rect 71748 83993 74748 84005
rect 71748 83613 71882 83993
rect 72262 83613 72274 83993
rect 72654 83613 72666 83993
rect 73046 83613 73058 83993
rect 73438 83613 73450 83993
rect 73830 83613 73842 83993
rect 74222 83613 74234 83993
rect 74614 83613 74748 83993
rect 71748 83601 74748 83613
rect 71748 83221 71882 83601
rect 72262 83221 72274 83601
rect 72654 83221 72666 83601
rect 73046 83221 73058 83601
rect 73438 83221 73450 83601
rect 73830 83221 73842 83601
rect 74222 83221 74234 83601
rect 74614 83221 74748 83601
rect 71748 83209 74748 83221
rect 71748 82829 71882 83209
rect 72262 82829 72274 83209
rect 72654 82829 72666 83209
rect 73046 82829 73058 83209
rect 73438 82829 73450 83209
rect 73830 82829 73842 83209
rect 74222 82829 74234 83209
rect 74614 82829 74748 83209
rect 71748 78510 74748 82829
rect 71748 78130 71882 78510
rect 72262 78130 72274 78510
rect 72654 78130 72666 78510
rect 73046 78130 73058 78510
rect 73438 78130 73450 78510
rect 73830 78130 73842 78510
rect 74222 78130 74234 78510
rect 74614 78130 74748 78510
rect 71748 74566 74748 78130
rect 71748 74186 71882 74566
rect 72262 74186 72274 74566
rect 72654 74186 72666 74566
rect 73046 74186 73058 74566
rect 73438 74186 73450 74566
rect 73830 74186 73842 74566
rect 74222 74186 74234 74566
rect 74614 74186 74748 74566
rect 71748 74174 74748 74186
rect 71748 73794 71882 74174
rect 72262 73794 72274 74174
rect 72654 73794 72666 74174
rect 73046 73794 73058 74174
rect 73438 73794 73450 74174
rect 73830 73794 73842 74174
rect 74222 73794 74234 74174
rect 74614 73794 74748 74174
rect 71748 73782 74748 73794
rect 71748 73402 71882 73782
rect 72262 73402 72274 73782
rect 72654 73402 72666 73782
rect 73046 73402 73058 73782
rect 73438 73402 73450 73782
rect 73830 73402 73842 73782
rect 74222 73402 74234 73782
rect 74614 73402 74748 73782
rect 71748 73390 74748 73402
rect 71748 73010 71882 73390
rect 72262 73010 72274 73390
rect 72654 73010 72666 73390
rect 73046 73010 73058 73390
rect 73438 73010 73450 73390
rect 73830 73010 73842 73390
rect 74222 73010 74234 73390
rect 74614 73010 74748 73390
rect 71748 72998 74748 73010
rect 71748 72618 71882 72998
rect 72262 72618 72274 72998
rect 72654 72618 72666 72998
rect 73046 72618 73058 72998
rect 73438 72618 73450 72998
rect 73830 72618 73842 72998
rect 74222 72618 74234 72998
rect 74614 72618 74748 72998
rect 71748 72606 74748 72618
rect 71748 72226 71882 72606
rect 72262 72226 72274 72606
rect 72654 72226 72666 72606
rect 73046 72226 73058 72606
rect 73438 72226 73450 72606
rect 73830 72226 73842 72606
rect 74222 72226 74234 72606
rect 74614 72226 74748 72606
rect 71748 72214 74748 72226
rect 71748 71834 71882 72214
rect 72262 71834 72274 72214
rect 72654 71834 72666 72214
rect 73046 71834 73058 72214
rect 73438 71834 73450 72214
rect 73830 71834 73842 72214
rect 74222 71834 74234 72214
rect 74614 71834 74748 72214
rect 71748 71700 74748 71834
rect 78148 151942 78588 152076
rect 78148 151562 78178 151942
rect 78558 151562 78588 151942
rect 78148 151550 78588 151562
rect 78148 151170 78178 151550
rect 78558 151170 78588 151550
rect 78148 151158 78588 151170
rect 78148 150778 78178 151158
rect 78558 150778 78588 151158
rect 78148 150766 78588 150778
rect 78148 150386 78178 150766
rect 78558 150386 78588 150766
rect 78148 150374 78588 150386
rect 78148 149994 78178 150374
rect 78558 149994 78588 150374
rect 78148 149982 78588 149994
rect 78148 149602 78178 149982
rect 78558 149602 78588 149982
rect 78148 149590 78588 149602
rect 78148 149210 78178 149590
rect 78558 149210 78588 149590
rect 78148 147482 78588 149210
rect 78148 147358 78222 147482
rect 78346 147358 78390 147482
rect 78514 147358 78588 147482
rect 78148 145970 78588 147358
rect 78148 145846 78222 145970
rect 78346 145846 78390 145970
rect 78514 145846 78588 145970
rect 78148 144458 78588 145846
rect 78148 144334 78222 144458
rect 78346 144334 78390 144458
rect 78514 144334 78588 144458
rect 78148 142946 78588 144334
rect 78148 142822 78222 142946
rect 78346 142822 78390 142946
rect 78514 142822 78588 142946
rect 78148 141434 78588 142822
rect 78148 141310 78222 141434
rect 78346 141310 78390 141434
rect 78514 141310 78588 141434
rect 78148 139922 78588 141310
rect 78148 139798 78222 139922
rect 78346 139798 78390 139922
rect 78514 139798 78588 139922
rect 78148 138990 78588 139798
rect 78148 138610 78178 138990
rect 78558 138610 78588 138990
rect 78148 138410 78588 138610
rect 78148 138286 78222 138410
rect 78346 138286 78390 138410
rect 78514 138286 78588 138410
rect 78148 136898 78588 138286
rect 78148 136774 78222 136898
rect 78346 136774 78390 136898
rect 78514 136774 78588 136898
rect 78148 135386 78588 136774
rect 78148 135262 78222 135386
rect 78346 135262 78390 135386
rect 78514 135262 78588 135386
rect 78148 133874 78588 135262
rect 78148 133750 78222 133874
rect 78346 133750 78390 133874
rect 78514 133750 78588 133874
rect 78148 132362 78588 133750
rect 78148 132238 78222 132362
rect 78346 132238 78390 132362
rect 78514 132238 78588 132362
rect 78148 130850 78588 132238
rect 78148 130726 78222 130850
rect 78346 130726 78390 130850
rect 78514 130726 78588 130850
rect 78148 129338 78588 130726
rect 78148 129214 78222 129338
rect 78346 129214 78390 129338
rect 78514 129214 78588 129338
rect 78148 127826 78588 129214
rect 78148 127702 78222 127826
rect 78346 127702 78390 127826
rect 78514 127702 78588 127826
rect 78148 126314 78588 127702
rect 78148 126190 78222 126314
rect 78346 126190 78390 126314
rect 78514 126190 78588 126314
rect 78148 124802 78588 126190
rect 78148 124678 78222 124802
rect 78346 124678 78390 124802
rect 78514 124678 78588 124802
rect 78148 123870 78588 124678
rect 78148 123490 78178 123870
rect 78558 123490 78588 123870
rect 78148 123290 78588 123490
rect 78148 123166 78222 123290
rect 78346 123166 78390 123290
rect 78514 123166 78588 123290
rect 78148 121778 78588 123166
rect 78148 121654 78222 121778
rect 78346 121654 78390 121778
rect 78514 121654 78588 121778
rect 78148 120266 78588 121654
rect 78148 120142 78222 120266
rect 78346 120142 78390 120266
rect 78514 120142 78588 120266
rect 78148 118754 78588 120142
rect 78148 118630 78222 118754
rect 78346 118630 78390 118754
rect 78514 118630 78588 118754
rect 78148 117242 78588 118630
rect 78148 117118 78222 117242
rect 78346 117118 78390 117242
rect 78514 117118 78588 117242
rect 78148 115730 78588 117118
rect 78148 115606 78222 115730
rect 78346 115606 78390 115730
rect 78514 115606 78588 115730
rect 78148 114218 78588 115606
rect 78148 114094 78222 114218
rect 78346 114094 78390 114218
rect 78514 114094 78588 114218
rect 78148 112706 78588 114094
rect 78148 112582 78222 112706
rect 78346 112582 78390 112706
rect 78514 112582 78588 112706
rect 78148 111194 78588 112582
rect 78148 111070 78222 111194
rect 78346 111070 78390 111194
rect 78514 111070 78588 111194
rect 78148 109682 78588 111070
rect 78148 109558 78222 109682
rect 78346 109558 78390 109682
rect 78514 109558 78588 109682
rect 78148 108750 78588 109558
rect 78148 108370 78178 108750
rect 78558 108370 78588 108750
rect 78148 108170 78588 108370
rect 78148 108046 78222 108170
rect 78346 108046 78390 108170
rect 78514 108046 78588 108170
rect 78148 106658 78588 108046
rect 78148 106534 78222 106658
rect 78346 106534 78390 106658
rect 78514 106534 78588 106658
rect 78148 105146 78588 106534
rect 78148 105022 78222 105146
rect 78346 105022 78390 105146
rect 78514 105022 78588 105146
rect 78148 103634 78588 105022
rect 78148 103510 78222 103634
rect 78346 103510 78390 103634
rect 78514 103510 78588 103634
rect 78148 102122 78588 103510
rect 78148 101998 78222 102122
rect 78346 101998 78390 102122
rect 78514 101998 78588 102122
rect 78148 100610 78588 101998
rect 78148 100486 78222 100610
rect 78346 100486 78390 100610
rect 78514 100486 78588 100610
rect 78148 99098 78588 100486
rect 78148 98974 78222 99098
rect 78346 98974 78390 99098
rect 78514 98974 78588 99098
rect 78148 97586 78588 98974
rect 78148 97462 78222 97586
rect 78346 97462 78390 97586
rect 78514 97462 78588 97586
rect 78148 96074 78588 97462
rect 78148 95950 78222 96074
rect 78346 95950 78390 96074
rect 78514 95950 78588 96074
rect 78148 94562 78588 95950
rect 78148 94438 78222 94562
rect 78346 94438 78390 94562
rect 78514 94438 78588 94562
rect 78148 93630 78588 94438
rect 78148 93250 78178 93630
rect 78558 93250 78588 93630
rect 78148 93050 78588 93250
rect 78148 92926 78222 93050
rect 78346 92926 78390 93050
rect 78514 92926 78588 93050
rect 78148 91538 78588 92926
rect 78148 91414 78222 91538
rect 78346 91414 78390 91538
rect 78514 91414 78588 91538
rect 78148 90026 78588 91414
rect 78148 89902 78222 90026
rect 78346 89902 78390 90026
rect 78514 89902 78588 90026
rect 78148 88514 78588 89902
rect 78148 88390 78222 88514
rect 78346 88390 78390 88514
rect 78514 88390 78588 88514
rect 78148 87002 78588 88390
rect 78148 86878 78222 87002
rect 78346 86878 78390 87002
rect 78514 86878 78588 87002
rect 78148 85490 78588 86878
rect 78148 85366 78222 85490
rect 78346 85366 78390 85490
rect 78514 85366 78588 85490
rect 78148 83978 78588 85366
rect 78148 83854 78222 83978
rect 78346 83854 78390 83978
rect 78514 83854 78588 83978
rect 78148 82466 78588 83854
rect 78148 82342 78222 82466
rect 78346 82342 78390 82466
rect 78514 82342 78588 82466
rect 78148 80954 78588 82342
rect 78148 80830 78222 80954
rect 78346 80830 78390 80954
rect 78514 80830 78588 80954
rect 78148 79442 78588 80830
rect 78148 79318 78222 79442
rect 78346 79318 78390 79442
rect 78514 79318 78588 79442
rect 78148 78510 78588 79318
rect 78148 78130 78178 78510
rect 78558 78130 78588 78510
rect 78148 77930 78588 78130
rect 78148 77806 78222 77930
rect 78346 77806 78390 77930
rect 78514 77806 78588 77930
rect 78148 76418 78588 77806
rect 78148 76294 78222 76418
rect 78346 76294 78390 76418
rect 78514 76294 78588 76418
rect 78148 74566 78588 76294
rect 78148 74186 78178 74566
rect 78558 74186 78588 74566
rect 78148 74174 78588 74186
rect 78148 73794 78178 74174
rect 78558 73794 78588 74174
rect 78148 73782 78588 73794
rect 78148 73402 78178 73782
rect 78558 73402 78588 73782
rect 78148 73390 78588 73402
rect 78148 73010 78178 73390
rect 78558 73010 78588 73390
rect 78148 72998 78588 73010
rect 78148 72618 78178 72998
rect 78558 72618 78588 72998
rect 78148 72606 78588 72618
rect 78148 72226 78178 72606
rect 78558 72226 78588 72606
rect 78148 72214 78588 72226
rect 78148 71834 78178 72214
rect 78558 71834 78588 72214
rect 78148 71700 78588 71834
rect 79388 148238 79828 153210
rect 94508 155942 94948 156076
rect 94508 155562 94538 155942
rect 94918 155562 94948 155942
rect 94508 155550 94948 155562
rect 94508 155170 94538 155550
rect 94918 155170 94948 155550
rect 94508 155158 94948 155170
rect 94508 154778 94538 155158
rect 94918 154778 94948 155158
rect 94508 154766 94948 154778
rect 94508 154386 94538 154766
rect 94918 154386 94948 154766
rect 94508 154374 94948 154386
rect 94508 153994 94538 154374
rect 94918 153994 94948 154374
rect 94508 153982 94948 153994
rect 94508 153602 94538 153982
rect 94918 153602 94948 153982
rect 94508 153590 94948 153602
rect 94508 153210 94538 153590
rect 94918 153210 94948 153590
rect 79388 148114 79462 148238
rect 79586 148114 79630 148238
rect 79754 148114 79828 148238
rect 79388 146726 79828 148114
rect 79388 146602 79462 146726
rect 79586 146602 79630 146726
rect 79754 146602 79828 146726
rect 79388 145214 79828 146602
rect 79388 145090 79462 145214
rect 79586 145090 79630 145214
rect 79754 145090 79828 145214
rect 79388 143702 79828 145090
rect 79388 143578 79462 143702
rect 79586 143578 79630 143702
rect 79754 143578 79828 143702
rect 79388 142190 79828 143578
rect 79388 142066 79462 142190
rect 79586 142066 79630 142190
rect 79754 142066 79828 142190
rect 79388 140678 79828 142066
rect 79388 140554 79462 140678
rect 79586 140554 79630 140678
rect 79754 140554 79828 140678
rect 79388 140230 79828 140554
rect 79388 139850 79418 140230
rect 79798 139850 79828 140230
rect 79388 139166 79828 139850
rect 79388 139042 79462 139166
rect 79586 139042 79630 139166
rect 79754 139042 79828 139166
rect 79388 137654 79828 139042
rect 79388 137530 79462 137654
rect 79586 137530 79630 137654
rect 79754 137530 79828 137654
rect 79388 136142 79828 137530
rect 79388 136018 79462 136142
rect 79586 136018 79630 136142
rect 79754 136018 79828 136142
rect 79388 134630 79828 136018
rect 79388 134506 79462 134630
rect 79586 134506 79630 134630
rect 79754 134506 79828 134630
rect 79388 133118 79828 134506
rect 79388 132994 79462 133118
rect 79586 132994 79630 133118
rect 79754 132994 79828 133118
rect 79388 131606 79828 132994
rect 79388 131482 79462 131606
rect 79586 131482 79630 131606
rect 79754 131482 79828 131606
rect 79388 130094 79828 131482
rect 79388 129970 79462 130094
rect 79586 129970 79630 130094
rect 79754 129970 79828 130094
rect 79388 128582 79828 129970
rect 79388 128458 79462 128582
rect 79586 128458 79630 128582
rect 79754 128458 79828 128582
rect 79388 127070 79828 128458
rect 79388 126946 79462 127070
rect 79586 126946 79630 127070
rect 79754 126946 79828 127070
rect 79388 125558 79828 126946
rect 79388 125434 79462 125558
rect 79586 125434 79630 125558
rect 79754 125434 79828 125558
rect 79388 125110 79828 125434
rect 79388 124730 79418 125110
rect 79798 124730 79828 125110
rect 79388 124046 79828 124730
rect 79388 123922 79462 124046
rect 79586 123922 79630 124046
rect 79754 123922 79828 124046
rect 79388 122534 79828 123922
rect 79388 122410 79462 122534
rect 79586 122410 79630 122534
rect 79754 122410 79828 122534
rect 79388 121022 79828 122410
rect 79388 120898 79462 121022
rect 79586 120898 79630 121022
rect 79754 120898 79828 121022
rect 79388 119510 79828 120898
rect 79388 119386 79462 119510
rect 79586 119386 79630 119510
rect 79754 119386 79828 119510
rect 79388 117998 79828 119386
rect 79388 117874 79462 117998
rect 79586 117874 79630 117998
rect 79754 117874 79828 117998
rect 79388 116486 79828 117874
rect 79388 116362 79462 116486
rect 79586 116362 79630 116486
rect 79754 116362 79828 116486
rect 79388 114974 79828 116362
rect 79388 114850 79462 114974
rect 79586 114850 79630 114974
rect 79754 114850 79828 114974
rect 79388 113462 79828 114850
rect 79388 113338 79462 113462
rect 79586 113338 79630 113462
rect 79754 113338 79828 113462
rect 79388 111950 79828 113338
rect 79388 111826 79462 111950
rect 79586 111826 79630 111950
rect 79754 111826 79828 111950
rect 79388 110438 79828 111826
rect 79388 110314 79462 110438
rect 79586 110314 79630 110438
rect 79754 110314 79828 110438
rect 79388 109990 79828 110314
rect 79388 109610 79418 109990
rect 79798 109610 79828 109990
rect 79388 108926 79828 109610
rect 79388 108802 79462 108926
rect 79586 108802 79630 108926
rect 79754 108802 79828 108926
rect 79388 107414 79828 108802
rect 79388 107290 79462 107414
rect 79586 107290 79630 107414
rect 79754 107290 79828 107414
rect 79388 105902 79828 107290
rect 79388 105778 79462 105902
rect 79586 105778 79630 105902
rect 79754 105778 79828 105902
rect 79388 104390 79828 105778
rect 79388 104266 79462 104390
rect 79586 104266 79630 104390
rect 79754 104266 79828 104390
rect 79388 102878 79828 104266
rect 79388 102754 79462 102878
rect 79586 102754 79630 102878
rect 79754 102754 79828 102878
rect 79388 101366 79828 102754
rect 79388 101242 79462 101366
rect 79586 101242 79630 101366
rect 79754 101242 79828 101366
rect 79388 99854 79828 101242
rect 79388 99730 79462 99854
rect 79586 99730 79630 99854
rect 79754 99730 79828 99854
rect 79388 98342 79828 99730
rect 79388 98218 79462 98342
rect 79586 98218 79630 98342
rect 79754 98218 79828 98342
rect 79388 96830 79828 98218
rect 79388 96706 79462 96830
rect 79586 96706 79630 96830
rect 79754 96706 79828 96830
rect 79388 95318 79828 96706
rect 79388 95194 79462 95318
rect 79586 95194 79630 95318
rect 79754 95194 79828 95318
rect 79388 94870 79828 95194
rect 79388 94490 79418 94870
rect 79798 94490 79828 94870
rect 79388 93806 79828 94490
rect 79388 93682 79462 93806
rect 79586 93682 79630 93806
rect 79754 93682 79828 93806
rect 79388 92294 79828 93682
rect 79388 92170 79462 92294
rect 79586 92170 79630 92294
rect 79754 92170 79828 92294
rect 79388 90782 79828 92170
rect 79388 90658 79462 90782
rect 79586 90658 79630 90782
rect 79754 90658 79828 90782
rect 79388 89270 79828 90658
rect 79388 89146 79462 89270
rect 79586 89146 79630 89270
rect 79754 89146 79828 89270
rect 79388 87758 79828 89146
rect 79388 87634 79462 87758
rect 79586 87634 79630 87758
rect 79754 87634 79828 87758
rect 79388 86246 79828 87634
rect 79388 86122 79462 86246
rect 79586 86122 79630 86246
rect 79754 86122 79828 86246
rect 79388 84734 79828 86122
rect 79388 84610 79462 84734
rect 79586 84610 79630 84734
rect 79754 84610 79828 84734
rect 79388 83222 79828 84610
rect 79388 83098 79462 83222
rect 79586 83098 79630 83222
rect 79754 83098 79828 83222
rect 79388 81710 79828 83098
rect 79388 81586 79462 81710
rect 79586 81586 79630 81710
rect 79754 81586 79828 81710
rect 79388 80198 79828 81586
rect 79388 80074 79462 80198
rect 79586 80074 79630 80198
rect 79754 80074 79828 80198
rect 79388 79750 79828 80074
rect 79388 79370 79418 79750
rect 79798 79370 79828 79750
rect 79388 78686 79828 79370
rect 79388 78562 79462 78686
rect 79586 78562 79630 78686
rect 79754 78562 79828 78686
rect 79388 77174 79828 78562
rect 79388 77050 79462 77174
rect 79586 77050 79630 77174
rect 79754 77050 79828 77174
rect 79388 75662 79828 77050
rect 79388 75538 79462 75662
rect 79586 75538 79630 75662
rect 79754 75538 79828 75662
rect 67748 70186 67882 70566
rect 68262 70186 68274 70566
rect 68654 70186 68666 70566
rect 69046 70186 69058 70566
rect 69438 70186 69450 70566
rect 69830 70186 69842 70566
rect 70222 70186 70234 70566
rect 70614 70186 70748 70566
rect 67748 70174 70748 70186
rect 67748 69794 67882 70174
rect 68262 69794 68274 70174
rect 68654 69794 68666 70174
rect 69046 69794 69058 70174
rect 69438 69794 69450 70174
rect 69830 69794 69842 70174
rect 70222 69794 70234 70174
rect 70614 69794 70748 70174
rect 67748 69782 70748 69794
rect 67748 69402 67882 69782
rect 68262 69402 68274 69782
rect 68654 69402 68666 69782
rect 69046 69402 69058 69782
rect 69438 69402 69450 69782
rect 69830 69402 69842 69782
rect 70222 69402 70234 69782
rect 70614 69402 70748 69782
rect 67748 69390 70748 69402
rect 67748 69010 67882 69390
rect 68262 69010 68274 69390
rect 68654 69010 68666 69390
rect 69046 69010 69058 69390
rect 69438 69010 69450 69390
rect 69830 69010 69842 69390
rect 70222 69010 70234 69390
rect 70614 69010 70748 69390
rect 67748 68998 70748 69010
rect 67748 68618 67882 68998
rect 68262 68618 68274 68998
rect 68654 68618 68666 68998
rect 69046 68618 69058 68998
rect 69438 68618 69450 68998
rect 69830 68618 69842 68998
rect 70222 68618 70234 68998
rect 70614 68618 70748 68998
rect 67748 68606 70748 68618
rect 67748 68226 67882 68606
rect 68262 68226 68274 68606
rect 68654 68226 68666 68606
rect 69046 68226 69058 68606
rect 69438 68226 69450 68606
rect 69830 68226 69842 68606
rect 70222 68226 70234 68606
rect 70614 68226 70748 68606
rect 67748 68214 70748 68226
rect 67748 67834 67882 68214
rect 68262 67834 68274 68214
rect 68654 67834 68666 68214
rect 69046 67834 69058 68214
rect 69438 67834 69450 68214
rect 69830 67834 69842 68214
rect 70222 67834 70234 68214
rect 70614 67834 70748 68214
rect 67748 67700 70748 67834
rect 79388 70566 79828 75538
rect 93268 151942 93708 152076
rect 93268 151562 93298 151942
rect 93678 151562 93708 151942
rect 93268 151550 93708 151562
rect 93268 151170 93298 151550
rect 93678 151170 93708 151550
rect 93268 151158 93708 151170
rect 93268 150778 93298 151158
rect 93678 150778 93708 151158
rect 93268 150766 93708 150778
rect 93268 150386 93298 150766
rect 93678 150386 93708 150766
rect 93268 150374 93708 150386
rect 93268 149994 93298 150374
rect 93678 149994 93708 150374
rect 93268 149982 93708 149994
rect 93268 149602 93298 149982
rect 93678 149602 93708 149982
rect 93268 149590 93708 149602
rect 93268 149210 93298 149590
rect 93678 149210 93708 149590
rect 93268 147482 93708 149210
rect 93268 147358 93342 147482
rect 93466 147358 93510 147482
rect 93634 147358 93708 147482
rect 93268 145970 93708 147358
rect 93268 145846 93342 145970
rect 93466 145846 93510 145970
rect 93634 145846 93708 145970
rect 93268 144458 93708 145846
rect 93268 144334 93342 144458
rect 93466 144334 93510 144458
rect 93634 144334 93708 144458
rect 93268 142946 93708 144334
rect 93268 142822 93342 142946
rect 93466 142822 93510 142946
rect 93634 142822 93708 142946
rect 93268 141434 93708 142822
rect 93268 141310 93342 141434
rect 93466 141310 93510 141434
rect 93634 141310 93708 141434
rect 93268 139922 93708 141310
rect 93268 139798 93342 139922
rect 93466 139798 93510 139922
rect 93634 139798 93708 139922
rect 93268 138990 93708 139798
rect 93268 138610 93298 138990
rect 93678 138610 93708 138990
rect 93268 138410 93708 138610
rect 93268 138286 93342 138410
rect 93466 138286 93510 138410
rect 93634 138286 93708 138410
rect 93268 136898 93708 138286
rect 93268 136774 93342 136898
rect 93466 136774 93510 136898
rect 93634 136774 93708 136898
rect 93268 135386 93708 136774
rect 93268 135262 93342 135386
rect 93466 135262 93510 135386
rect 93634 135262 93708 135386
rect 93268 133874 93708 135262
rect 93268 133750 93342 133874
rect 93466 133750 93510 133874
rect 93634 133750 93708 133874
rect 93268 132362 93708 133750
rect 93268 132238 93342 132362
rect 93466 132238 93510 132362
rect 93634 132238 93708 132362
rect 93268 130850 93708 132238
rect 93268 130726 93342 130850
rect 93466 130726 93510 130850
rect 93634 130726 93708 130850
rect 93268 129338 93708 130726
rect 93268 129214 93342 129338
rect 93466 129214 93510 129338
rect 93634 129214 93708 129338
rect 93268 127826 93708 129214
rect 93268 127702 93342 127826
rect 93466 127702 93510 127826
rect 93634 127702 93708 127826
rect 93268 126314 93708 127702
rect 93268 126190 93342 126314
rect 93466 126190 93510 126314
rect 93634 126190 93708 126314
rect 93268 124802 93708 126190
rect 93268 124678 93342 124802
rect 93466 124678 93510 124802
rect 93634 124678 93708 124802
rect 93268 123870 93708 124678
rect 93268 123490 93298 123870
rect 93678 123490 93708 123870
rect 93268 123290 93708 123490
rect 93268 123166 93342 123290
rect 93466 123166 93510 123290
rect 93634 123166 93708 123290
rect 93268 121778 93708 123166
rect 93268 121654 93342 121778
rect 93466 121654 93510 121778
rect 93634 121654 93708 121778
rect 93268 120266 93708 121654
rect 93268 120142 93342 120266
rect 93466 120142 93510 120266
rect 93634 120142 93708 120266
rect 93268 118754 93708 120142
rect 93268 118630 93342 118754
rect 93466 118630 93510 118754
rect 93634 118630 93708 118754
rect 93268 117242 93708 118630
rect 93268 117118 93342 117242
rect 93466 117118 93510 117242
rect 93634 117118 93708 117242
rect 93268 115730 93708 117118
rect 93268 115606 93342 115730
rect 93466 115606 93510 115730
rect 93634 115606 93708 115730
rect 93268 114218 93708 115606
rect 93268 114094 93342 114218
rect 93466 114094 93510 114218
rect 93634 114094 93708 114218
rect 93268 112706 93708 114094
rect 93268 112582 93342 112706
rect 93466 112582 93510 112706
rect 93634 112582 93708 112706
rect 93268 111194 93708 112582
rect 93268 111070 93342 111194
rect 93466 111070 93510 111194
rect 93634 111070 93708 111194
rect 93268 109682 93708 111070
rect 93268 109558 93342 109682
rect 93466 109558 93510 109682
rect 93634 109558 93708 109682
rect 93268 108750 93708 109558
rect 93268 108370 93298 108750
rect 93678 108370 93708 108750
rect 93268 108170 93708 108370
rect 93268 108046 93342 108170
rect 93466 108046 93510 108170
rect 93634 108046 93708 108170
rect 93268 106658 93708 108046
rect 93268 106534 93342 106658
rect 93466 106534 93510 106658
rect 93634 106534 93708 106658
rect 93268 105146 93708 106534
rect 93268 105022 93342 105146
rect 93466 105022 93510 105146
rect 93634 105022 93708 105146
rect 93268 103634 93708 105022
rect 93268 103510 93342 103634
rect 93466 103510 93510 103634
rect 93634 103510 93708 103634
rect 93268 102122 93708 103510
rect 93268 101998 93342 102122
rect 93466 101998 93510 102122
rect 93634 101998 93708 102122
rect 93268 100610 93708 101998
rect 93268 100486 93342 100610
rect 93466 100486 93510 100610
rect 93634 100486 93708 100610
rect 93268 99098 93708 100486
rect 93268 98974 93342 99098
rect 93466 98974 93510 99098
rect 93634 98974 93708 99098
rect 93268 97586 93708 98974
rect 93268 97462 93342 97586
rect 93466 97462 93510 97586
rect 93634 97462 93708 97586
rect 93268 96074 93708 97462
rect 93268 95950 93342 96074
rect 93466 95950 93510 96074
rect 93634 95950 93708 96074
rect 93268 94562 93708 95950
rect 93268 94438 93342 94562
rect 93466 94438 93510 94562
rect 93634 94438 93708 94562
rect 93268 93630 93708 94438
rect 93268 93250 93298 93630
rect 93678 93250 93708 93630
rect 93268 93050 93708 93250
rect 93268 92926 93342 93050
rect 93466 92926 93510 93050
rect 93634 92926 93708 93050
rect 93268 91538 93708 92926
rect 93268 91414 93342 91538
rect 93466 91414 93510 91538
rect 93634 91414 93708 91538
rect 93268 90026 93708 91414
rect 93268 89902 93342 90026
rect 93466 89902 93510 90026
rect 93634 89902 93708 90026
rect 93268 88514 93708 89902
rect 93268 88390 93342 88514
rect 93466 88390 93510 88514
rect 93634 88390 93708 88514
rect 93268 87002 93708 88390
rect 93268 86878 93342 87002
rect 93466 86878 93510 87002
rect 93634 86878 93708 87002
rect 93268 85490 93708 86878
rect 93268 85366 93342 85490
rect 93466 85366 93510 85490
rect 93634 85366 93708 85490
rect 93268 83978 93708 85366
rect 93268 83854 93342 83978
rect 93466 83854 93510 83978
rect 93634 83854 93708 83978
rect 93268 82466 93708 83854
rect 93268 82342 93342 82466
rect 93466 82342 93510 82466
rect 93634 82342 93708 82466
rect 93268 80954 93708 82342
rect 93268 80830 93342 80954
rect 93466 80830 93510 80954
rect 93634 80830 93708 80954
rect 93268 79442 93708 80830
rect 93268 79318 93342 79442
rect 93466 79318 93510 79442
rect 93634 79318 93708 79442
rect 93268 78510 93708 79318
rect 93268 78130 93298 78510
rect 93678 78130 93708 78510
rect 93268 77930 93708 78130
rect 93268 77806 93342 77930
rect 93466 77806 93510 77930
rect 93634 77806 93708 77930
rect 93268 76418 93708 77806
rect 93268 76294 93342 76418
rect 93466 76294 93510 76418
rect 93634 76294 93708 76418
rect 93268 74566 93708 76294
rect 93268 74186 93298 74566
rect 93678 74186 93708 74566
rect 93268 74174 93708 74186
rect 93268 73794 93298 74174
rect 93678 73794 93708 74174
rect 93268 73782 93708 73794
rect 93268 73402 93298 73782
rect 93678 73402 93708 73782
rect 93268 73390 93708 73402
rect 93268 73010 93298 73390
rect 93678 73010 93708 73390
rect 93268 72998 93708 73010
rect 93268 72618 93298 72998
rect 93678 72618 93708 72998
rect 93268 72606 93708 72618
rect 93268 72226 93298 72606
rect 93678 72226 93708 72606
rect 93268 72214 93708 72226
rect 93268 71834 93298 72214
rect 93678 71834 93708 72214
rect 93268 71700 93708 71834
rect 94508 148238 94948 153210
rect 109628 155942 110068 156076
rect 109628 155562 109658 155942
rect 110038 155562 110068 155942
rect 109628 155550 110068 155562
rect 109628 155170 109658 155550
rect 110038 155170 110068 155550
rect 109628 155158 110068 155170
rect 109628 154778 109658 155158
rect 110038 154778 110068 155158
rect 109628 154766 110068 154778
rect 109628 154386 109658 154766
rect 110038 154386 110068 154766
rect 109628 154374 110068 154386
rect 109628 153994 109658 154374
rect 110038 153994 110068 154374
rect 109628 153982 110068 153994
rect 109628 153602 109658 153982
rect 110038 153602 110068 153982
rect 109628 153590 110068 153602
rect 109628 153210 109658 153590
rect 110038 153210 110068 153590
rect 94508 148114 94582 148238
rect 94706 148114 94750 148238
rect 94874 148114 94948 148238
rect 94508 146726 94948 148114
rect 94508 146602 94582 146726
rect 94706 146602 94750 146726
rect 94874 146602 94948 146726
rect 94508 145214 94948 146602
rect 94508 145090 94582 145214
rect 94706 145090 94750 145214
rect 94874 145090 94948 145214
rect 94508 143702 94948 145090
rect 94508 143578 94582 143702
rect 94706 143578 94750 143702
rect 94874 143578 94948 143702
rect 94508 142190 94948 143578
rect 94508 142066 94582 142190
rect 94706 142066 94750 142190
rect 94874 142066 94948 142190
rect 94508 140678 94948 142066
rect 94508 140554 94582 140678
rect 94706 140554 94750 140678
rect 94874 140554 94948 140678
rect 94508 140230 94948 140554
rect 94508 139850 94538 140230
rect 94918 139850 94948 140230
rect 94508 139166 94948 139850
rect 94508 139042 94582 139166
rect 94706 139042 94750 139166
rect 94874 139042 94948 139166
rect 94508 137654 94948 139042
rect 94508 137530 94582 137654
rect 94706 137530 94750 137654
rect 94874 137530 94948 137654
rect 94508 136142 94948 137530
rect 94508 136018 94582 136142
rect 94706 136018 94750 136142
rect 94874 136018 94948 136142
rect 94508 134630 94948 136018
rect 94508 134506 94582 134630
rect 94706 134506 94750 134630
rect 94874 134506 94948 134630
rect 94508 133118 94948 134506
rect 94508 132994 94582 133118
rect 94706 132994 94750 133118
rect 94874 132994 94948 133118
rect 94508 131606 94948 132994
rect 94508 131482 94582 131606
rect 94706 131482 94750 131606
rect 94874 131482 94948 131606
rect 94508 130094 94948 131482
rect 94508 129970 94582 130094
rect 94706 129970 94750 130094
rect 94874 129970 94948 130094
rect 94508 128582 94948 129970
rect 94508 128458 94582 128582
rect 94706 128458 94750 128582
rect 94874 128458 94948 128582
rect 94508 127070 94948 128458
rect 94508 126946 94582 127070
rect 94706 126946 94750 127070
rect 94874 126946 94948 127070
rect 94508 125558 94948 126946
rect 94508 125434 94582 125558
rect 94706 125434 94750 125558
rect 94874 125434 94948 125558
rect 94508 125110 94948 125434
rect 94508 124730 94538 125110
rect 94918 124730 94948 125110
rect 94508 124046 94948 124730
rect 94508 123922 94582 124046
rect 94706 123922 94750 124046
rect 94874 123922 94948 124046
rect 94508 122534 94948 123922
rect 94508 122410 94582 122534
rect 94706 122410 94750 122534
rect 94874 122410 94948 122534
rect 94508 121022 94948 122410
rect 94508 120898 94582 121022
rect 94706 120898 94750 121022
rect 94874 120898 94948 121022
rect 94508 119510 94948 120898
rect 94508 119386 94582 119510
rect 94706 119386 94750 119510
rect 94874 119386 94948 119510
rect 94508 117998 94948 119386
rect 94508 117874 94582 117998
rect 94706 117874 94750 117998
rect 94874 117874 94948 117998
rect 94508 116486 94948 117874
rect 94508 116362 94582 116486
rect 94706 116362 94750 116486
rect 94874 116362 94948 116486
rect 94508 114974 94948 116362
rect 94508 114850 94582 114974
rect 94706 114850 94750 114974
rect 94874 114850 94948 114974
rect 94508 113462 94948 114850
rect 94508 113338 94582 113462
rect 94706 113338 94750 113462
rect 94874 113338 94948 113462
rect 94508 111950 94948 113338
rect 94508 111826 94582 111950
rect 94706 111826 94750 111950
rect 94874 111826 94948 111950
rect 94508 110438 94948 111826
rect 94508 110314 94582 110438
rect 94706 110314 94750 110438
rect 94874 110314 94948 110438
rect 94508 109990 94948 110314
rect 94508 109610 94538 109990
rect 94918 109610 94948 109990
rect 94508 108926 94948 109610
rect 94508 108802 94582 108926
rect 94706 108802 94750 108926
rect 94874 108802 94948 108926
rect 94508 107414 94948 108802
rect 94508 107290 94582 107414
rect 94706 107290 94750 107414
rect 94874 107290 94948 107414
rect 94508 105902 94948 107290
rect 94508 105778 94582 105902
rect 94706 105778 94750 105902
rect 94874 105778 94948 105902
rect 94508 104390 94948 105778
rect 94508 104266 94582 104390
rect 94706 104266 94750 104390
rect 94874 104266 94948 104390
rect 94508 102878 94948 104266
rect 94508 102754 94582 102878
rect 94706 102754 94750 102878
rect 94874 102754 94948 102878
rect 94508 101366 94948 102754
rect 94508 101242 94582 101366
rect 94706 101242 94750 101366
rect 94874 101242 94948 101366
rect 94508 99854 94948 101242
rect 94508 99730 94582 99854
rect 94706 99730 94750 99854
rect 94874 99730 94948 99854
rect 94508 98342 94948 99730
rect 94508 98218 94582 98342
rect 94706 98218 94750 98342
rect 94874 98218 94948 98342
rect 94508 96830 94948 98218
rect 94508 96706 94582 96830
rect 94706 96706 94750 96830
rect 94874 96706 94948 96830
rect 94508 95318 94948 96706
rect 94508 95194 94582 95318
rect 94706 95194 94750 95318
rect 94874 95194 94948 95318
rect 94508 94870 94948 95194
rect 94508 94490 94538 94870
rect 94918 94490 94948 94870
rect 94508 93806 94948 94490
rect 94508 93682 94582 93806
rect 94706 93682 94750 93806
rect 94874 93682 94948 93806
rect 94508 92294 94948 93682
rect 94508 92170 94582 92294
rect 94706 92170 94750 92294
rect 94874 92170 94948 92294
rect 94508 90782 94948 92170
rect 94508 90658 94582 90782
rect 94706 90658 94750 90782
rect 94874 90658 94948 90782
rect 94508 89270 94948 90658
rect 94508 89146 94582 89270
rect 94706 89146 94750 89270
rect 94874 89146 94948 89270
rect 94508 87758 94948 89146
rect 94508 87634 94582 87758
rect 94706 87634 94750 87758
rect 94874 87634 94948 87758
rect 94508 86246 94948 87634
rect 94508 86122 94582 86246
rect 94706 86122 94750 86246
rect 94874 86122 94948 86246
rect 94508 84734 94948 86122
rect 94508 84610 94582 84734
rect 94706 84610 94750 84734
rect 94874 84610 94948 84734
rect 94508 83222 94948 84610
rect 94508 83098 94582 83222
rect 94706 83098 94750 83222
rect 94874 83098 94948 83222
rect 94508 81710 94948 83098
rect 94508 81586 94582 81710
rect 94706 81586 94750 81710
rect 94874 81586 94948 81710
rect 94508 80198 94948 81586
rect 94508 80074 94582 80198
rect 94706 80074 94750 80198
rect 94874 80074 94948 80198
rect 94508 79750 94948 80074
rect 94508 79370 94538 79750
rect 94918 79370 94948 79750
rect 94508 78686 94948 79370
rect 94508 78562 94582 78686
rect 94706 78562 94750 78686
rect 94874 78562 94948 78686
rect 94508 77174 94948 78562
rect 94508 77050 94582 77174
rect 94706 77050 94750 77174
rect 94874 77050 94948 77174
rect 94508 75662 94948 77050
rect 94508 75538 94582 75662
rect 94706 75538 94750 75662
rect 94874 75538 94948 75662
rect 79388 70186 79418 70566
rect 79798 70186 79828 70566
rect 79388 70174 79828 70186
rect 79388 69794 79418 70174
rect 79798 69794 79828 70174
rect 79388 69782 79828 69794
rect 79388 69402 79418 69782
rect 79798 69402 79828 69782
rect 79388 69390 79828 69402
rect 79388 69010 79418 69390
rect 79798 69010 79828 69390
rect 79388 68998 79828 69010
rect 79388 68618 79418 68998
rect 79798 68618 79828 68998
rect 79388 68606 79828 68618
rect 79388 68226 79418 68606
rect 79798 68226 79828 68606
rect 79388 68214 79828 68226
rect 79388 67834 79418 68214
rect 79798 67834 79828 68214
rect 79388 67700 79828 67834
rect 94508 70566 94948 75538
rect 108388 151942 108828 152076
rect 108388 151562 108418 151942
rect 108798 151562 108828 151942
rect 108388 151550 108828 151562
rect 108388 151170 108418 151550
rect 108798 151170 108828 151550
rect 108388 151158 108828 151170
rect 108388 150778 108418 151158
rect 108798 150778 108828 151158
rect 108388 150766 108828 150778
rect 108388 150386 108418 150766
rect 108798 150386 108828 150766
rect 108388 150374 108828 150386
rect 108388 149994 108418 150374
rect 108798 149994 108828 150374
rect 108388 149982 108828 149994
rect 108388 149602 108418 149982
rect 108798 149602 108828 149982
rect 108388 149590 108828 149602
rect 108388 149210 108418 149590
rect 108798 149210 108828 149590
rect 108388 147482 108828 149210
rect 108388 147358 108462 147482
rect 108586 147358 108630 147482
rect 108754 147358 108828 147482
rect 108388 145970 108828 147358
rect 108388 145846 108462 145970
rect 108586 145846 108630 145970
rect 108754 145846 108828 145970
rect 108388 144458 108828 145846
rect 108388 144334 108462 144458
rect 108586 144334 108630 144458
rect 108754 144334 108828 144458
rect 108388 142946 108828 144334
rect 108388 142822 108462 142946
rect 108586 142822 108630 142946
rect 108754 142822 108828 142946
rect 108388 141434 108828 142822
rect 108388 141310 108462 141434
rect 108586 141310 108630 141434
rect 108754 141310 108828 141434
rect 108388 139922 108828 141310
rect 108388 139798 108462 139922
rect 108586 139798 108630 139922
rect 108754 139798 108828 139922
rect 108388 138990 108828 139798
rect 108388 138610 108418 138990
rect 108798 138610 108828 138990
rect 108388 138410 108828 138610
rect 108388 138286 108462 138410
rect 108586 138286 108630 138410
rect 108754 138286 108828 138410
rect 108388 136898 108828 138286
rect 108388 136774 108462 136898
rect 108586 136774 108630 136898
rect 108754 136774 108828 136898
rect 108388 135386 108828 136774
rect 108388 135262 108462 135386
rect 108586 135262 108630 135386
rect 108754 135262 108828 135386
rect 108388 133874 108828 135262
rect 108388 133750 108462 133874
rect 108586 133750 108630 133874
rect 108754 133750 108828 133874
rect 108388 132362 108828 133750
rect 108388 132238 108462 132362
rect 108586 132238 108630 132362
rect 108754 132238 108828 132362
rect 108388 130850 108828 132238
rect 108388 130726 108462 130850
rect 108586 130726 108630 130850
rect 108754 130726 108828 130850
rect 108388 129338 108828 130726
rect 108388 129214 108462 129338
rect 108586 129214 108630 129338
rect 108754 129214 108828 129338
rect 108388 127826 108828 129214
rect 108388 127702 108462 127826
rect 108586 127702 108630 127826
rect 108754 127702 108828 127826
rect 108388 126314 108828 127702
rect 108388 126190 108462 126314
rect 108586 126190 108630 126314
rect 108754 126190 108828 126314
rect 108388 124802 108828 126190
rect 108388 124678 108462 124802
rect 108586 124678 108630 124802
rect 108754 124678 108828 124802
rect 108388 123870 108828 124678
rect 108388 123490 108418 123870
rect 108798 123490 108828 123870
rect 108388 123290 108828 123490
rect 108388 123166 108462 123290
rect 108586 123166 108630 123290
rect 108754 123166 108828 123290
rect 108388 121778 108828 123166
rect 108388 121654 108462 121778
rect 108586 121654 108630 121778
rect 108754 121654 108828 121778
rect 108388 120266 108828 121654
rect 108388 120142 108462 120266
rect 108586 120142 108630 120266
rect 108754 120142 108828 120266
rect 108388 118754 108828 120142
rect 108388 118630 108462 118754
rect 108586 118630 108630 118754
rect 108754 118630 108828 118754
rect 108388 117242 108828 118630
rect 108388 117118 108462 117242
rect 108586 117118 108630 117242
rect 108754 117118 108828 117242
rect 108388 115730 108828 117118
rect 108388 115606 108462 115730
rect 108586 115606 108630 115730
rect 108754 115606 108828 115730
rect 108388 114218 108828 115606
rect 108388 114094 108462 114218
rect 108586 114094 108630 114218
rect 108754 114094 108828 114218
rect 108388 112706 108828 114094
rect 108388 112582 108462 112706
rect 108586 112582 108630 112706
rect 108754 112582 108828 112706
rect 108388 111194 108828 112582
rect 108388 111070 108462 111194
rect 108586 111070 108630 111194
rect 108754 111070 108828 111194
rect 108388 109682 108828 111070
rect 108388 109558 108462 109682
rect 108586 109558 108630 109682
rect 108754 109558 108828 109682
rect 108388 108750 108828 109558
rect 108388 108370 108418 108750
rect 108798 108370 108828 108750
rect 108388 108170 108828 108370
rect 108388 108046 108462 108170
rect 108586 108046 108630 108170
rect 108754 108046 108828 108170
rect 108388 106658 108828 108046
rect 108388 106534 108462 106658
rect 108586 106534 108630 106658
rect 108754 106534 108828 106658
rect 108388 105146 108828 106534
rect 108388 105022 108462 105146
rect 108586 105022 108630 105146
rect 108754 105022 108828 105146
rect 108388 103634 108828 105022
rect 108388 103510 108462 103634
rect 108586 103510 108630 103634
rect 108754 103510 108828 103634
rect 108388 102122 108828 103510
rect 108388 101998 108462 102122
rect 108586 101998 108630 102122
rect 108754 101998 108828 102122
rect 108388 100610 108828 101998
rect 108388 100486 108462 100610
rect 108586 100486 108630 100610
rect 108754 100486 108828 100610
rect 108388 99098 108828 100486
rect 108388 98974 108462 99098
rect 108586 98974 108630 99098
rect 108754 98974 108828 99098
rect 108388 97586 108828 98974
rect 108388 97462 108462 97586
rect 108586 97462 108630 97586
rect 108754 97462 108828 97586
rect 108388 96074 108828 97462
rect 108388 95950 108462 96074
rect 108586 95950 108630 96074
rect 108754 95950 108828 96074
rect 108388 94562 108828 95950
rect 108388 94438 108462 94562
rect 108586 94438 108630 94562
rect 108754 94438 108828 94562
rect 108388 93630 108828 94438
rect 108388 93250 108418 93630
rect 108798 93250 108828 93630
rect 108388 93050 108828 93250
rect 108388 92926 108462 93050
rect 108586 92926 108630 93050
rect 108754 92926 108828 93050
rect 108388 91538 108828 92926
rect 108388 91414 108462 91538
rect 108586 91414 108630 91538
rect 108754 91414 108828 91538
rect 108388 90026 108828 91414
rect 108388 89902 108462 90026
rect 108586 89902 108630 90026
rect 108754 89902 108828 90026
rect 108388 88514 108828 89902
rect 108388 88390 108462 88514
rect 108586 88390 108630 88514
rect 108754 88390 108828 88514
rect 108388 87002 108828 88390
rect 108388 86878 108462 87002
rect 108586 86878 108630 87002
rect 108754 86878 108828 87002
rect 108388 85490 108828 86878
rect 108388 85366 108462 85490
rect 108586 85366 108630 85490
rect 108754 85366 108828 85490
rect 108388 83978 108828 85366
rect 108388 83854 108462 83978
rect 108586 83854 108630 83978
rect 108754 83854 108828 83978
rect 108388 82466 108828 83854
rect 108388 82342 108462 82466
rect 108586 82342 108630 82466
rect 108754 82342 108828 82466
rect 108388 80954 108828 82342
rect 108388 80830 108462 80954
rect 108586 80830 108630 80954
rect 108754 80830 108828 80954
rect 108388 79442 108828 80830
rect 108388 79318 108462 79442
rect 108586 79318 108630 79442
rect 108754 79318 108828 79442
rect 108388 78510 108828 79318
rect 108388 78130 108418 78510
rect 108798 78130 108828 78510
rect 108388 77930 108828 78130
rect 108388 77806 108462 77930
rect 108586 77806 108630 77930
rect 108754 77806 108828 77930
rect 108388 76418 108828 77806
rect 108388 76294 108462 76418
rect 108586 76294 108630 76418
rect 108754 76294 108828 76418
rect 108388 74566 108828 76294
rect 108388 74186 108418 74566
rect 108798 74186 108828 74566
rect 108388 74174 108828 74186
rect 108388 73794 108418 74174
rect 108798 73794 108828 74174
rect 108388 73782 108828 73794
rect 108388 73402 108418 73782
rect 108798 73402 108828 73782
rect 108388 73390 108828 73402
rect 108388 73010 108418 73390
rect 108798 73010 108828 73390
rect 108388 72998 108828 73010
rect 108388 72618 108418 72998
rect 108798 72618 108828 72998
rect 108388 72606 108828 72618
rect 108388 72226 108418 72606
rect 108798 72226 108828 72606
rect 108388 72214 108828 72226
rect 108388 71834 108418 72214
rect 108798 71834 108828 72214
rect 108388 71700 108828 71834
rect 109628 148238 110068 153210
rect 124748 155942 125188 156076
rect 124748 155562 124778 155942
rect 125158 155562 125188 155942
rect 124748 155550 125188 155562
rect 124748 155170 124778 155550
rect 125158 155170 125188 155550
rect 124748 155158 125188 155170
rect 124748 154778 124778 155158
rect 125158 154778 125188 155158
rect 124748 154766 125188 154778
rect 124748 154386 124778 154766
rect 125158 154386 125188 154766
rect 124748 154374 125188 154386
rect 124748 153994 124778 154374
rect 125158 153994 125188 154374
rect 124748 153982 125188 153994
rect 124748 153602 124778 153982
rect 125158 153602 125188 153982
rect 124748 153590 125188 153602
rect 124748 153210 124778 153590
rect 125158 153210 125188 153590
rect 109628 148114 109702 148238
rect 109826 148114 109870 148238
rect 109994 148114 110068 148238
rect 109628 146726 110068 148114
rect 109628 146602 109702 146726
rect 109826 146602 109870 146726
rect 109994 146602 110068 146726
rect 109628 145214 110068 146602
rect 109628 145090 109702 145214
rect 109826 145090 109870 145214
rect 109994 145090 110068 145214
rect 109628 143702 110068 145090
rect 109628 143578 109702 143702
rect 109826 143578 109870 143702
rect 109994 143578 110068 143702
rect 109628 142190 110068 143578
rect 109628 142066 109702 142190
rect 109826 142066 109870 142190
rect 109994 142066 110068 142190
rect 109628 140678 110068 142066
rect 109628 140554 109702 140678
rect 109826 140554 109870 140678
rect 109994 140554 110068 140678
rect 109628 140230 110068 140554
rect 109628 139850 109658 140230
rect 110038 139850 110068 140230
rect 109628 139166 110068 139850
rect 109628 139042 109702 139166
rect 109826 139042 109870 139166
rect 109994 139042 110068 139166
rect 109628 137654 110068 139042
rect 109628 137530 109702 137654
rect 109826 137530 109870 137654
rect 109994 137530 110068 137654
rect 109628 136142 110068 137530
rect 109628 136018 109702 136142
rect 109826 136018 109870 136142
rect 109994 136018 110068 136142
rect 109628 134630 110068 136018
rect 109628 134506 109702 134630
rect 109826 134506 109870 134630
rect 109994 134506 110068 134630
rect 109628 133118 110068 134506
rect 109628 132994 109702 133118
rect 109826 132994 109870 133118
rect 109994 132994 110068 133118
rect 109628 131606 110068 132994
rect 109628 131482 109702 131606
rect 109826 131482 109870 131606
rect 109994 131482 110068 131606
rect 109628 130094 110068 131482
rect 109628 129970 109702 130094
rect 109826 129970 109870 130094
rect 109994 129970 110068 130094
rect 109628 128582 110068 129970
rect 109628 128458 109702 128582
rect 109826 128458 109870 128582
rect 109994 128458 110068 128582
rect 109628 127070 110068 128458
rect 109628 126946 109702 127070
rect 109826 126946 109870 127070
rect 109994 126946 110068 127070
rect 109628 125558 110068 126946
rect 109628 125434 109702 125558
rect 109826 125434 109870 125558
rect 109994 125434 110068 125558
rect 109628 125110 110068 125434
rect 109628 124730 109658 125110
rect 110038 124730 110068 125110
rect 109628 124046 110068 124730
rect 109628 123922 109702 124046
rect 109826 123922 109870 124046
rect 109994 123922 110068 124046
rect 109628 122534 110068 123922
rect 109628 122410 109702 122534
rect 109826 122410 109870 122534
rect 109994 122410 110068 122534
rect 109628 121022 110068 122410
rect 109628 120898 109702 121022
rect 109826 120898 109870 121022
rect 109994 120898 110068 121022
rect 109628 119510 110068 120898
rect 109628 119386 109702 119510
rect 109826 119386 109870 119510
rect 109994 119386 110068 119510
rect 109628 117998 110068 119386
rect 109628 117874 109702 117998
rect 109826 117874 109870 117998
rect 109994 117874 110068 117998
rect 109628 116486 110068 117874
rect 109628 116362 109702 116486
rect 109826 116362 109870 116486
rect 109994 116362 110068 116486
rect 109628 114974 110068 116362
rect 109628 114850 109702 114974
rect 109826 114850 109870 114974
rect 109994 114850 110068 114974
rect 109628 113462 110068 114850
rect 109628 113338 109702 113462
rect 109826 113338 109870 113462
rect 109994 113338 110068 113462
rect 109628 111950 110068 113338
rect 109628 111826 109702 111950
rect 109826 111826 109870 111950
rect 109994 111826 110068 111950
rect 109628 110438 110068 111826
rect 109628 110314 109702 110438
rect 109826 110314 109870 110438
rect 109994 110314 110068 110438
rect 109628 109990 110068 110314
rect 109628 109610 109658 109990
rect 110038 109610 110068 109990
rect 109628 108926 110068 109610
rect 109628 108802 109702 108926
rect 109826 108802 109870 108926
rect 109994 108802 110068 108926
rect 109628 107414 110068 108802
rect 109628 107290 109702 107414
rect 109826 107290 109870 107414
rect 109994 107290 110068 107414
rect 109628 105902 110068 107290
rect 109628 105778 109702 105902
rect 109826 105778 109870 105902
rect 109994 105778 110068 105902
rect 109628 104390 110068 105778
rect 109628 104266 109702 104390
rect 109826 104266 109870 104390
rect 109994 104266 110068 104390
rect 109628 102878 110068 104266
rect 109628 102754 109702 102878
rect 109826 102754 109870 102878
rect 109994 102754 110068 102878
rect 109628 101366 110068 102754
rect 109628 101242 109702 101366
rect 109826 101242 109870 101366
rect 109994 101242 110068 101366
rect 109628 99854 110068 101242
rect 109628 99730 109702 99854
rect 109826 99730 109870 99854
rect 109994 99730 110068 99854
rect 109628 98342 110068 99730
rect 109628 98218 109702 98342
rect 109826 98218 109870 98342
rect 109994 98218 110068 98342
rect 109628 96830 110068 98218
rect 109628 96706 109702 96830
rect 109826 96706 109870 96830
rect 109994 96706 110068 96830
rect 109628 95318 110068 96706
rect 109628 95194 109702 95318
rect 109826 95194 109870 95318
rect 109994 95194 110068 95318
rect 109628 94870 110068 95194
rect 109628 94490 109658 94870
rect 110038 94490 110068 94870
rect 109628 93806 110068 94490
rect 109628 93682 109702 93806
rect 109826 93682 109870 93806
rect 109994 93682 110068 93806
rect 109628 92294 110068 93682
rect 109628 92170 109702 92294
rect 109826 92170 109870 92294
rect 109994 92170 110068 92294
rect 109628 90782 110068 92170
rect 109628 90658 109702 90782
rect 109826 90658 109870 90782
rect 109994 90658 110068 90782
rect 109628 89270 110068 90658
rect 109628 89146 109702 89270
rect 109826 89146 109870 89270
rect 109994 89146 110068 89270
rect 109628 87758 110068 89146
rect 109628 87634 109702 87758
rect 109826 87634 109870 87758
rect 109994 87634 110068 87758
rect 109628 86246 110068 87634
rect 109628 86122 109702 86246
rect 109826 86122 109870 86246
rect 109994 86122 110068 86246
rect 109628 84734 110068 86122
rect 109628 84610 109702 84734
rect 109826 84610 109870 84734
rect 109994 84610 110068 84734
rect 109628 83222 110068 84610
rect 109628 83098 109702 83222
rect 109826 83098 109870 83222
rect 109994 83098 110068 83222
rect 109628 81710 110068 83098
rect 109628 81586 109702 81710
rect 109826 81586 109870 81710
rect 109994 81586 110068 81710
rect 109628 80198 110068 81586
rect 109628 80074 109702 80198
rect 109826 80074 109870 80198
rect 109994 80074 110068 80198
rect 109628 79750 110068 80074
rect 109628 79370 109658 79750
rect 110038 79370 110068 79750
rect 109628 78686 110068 79370
rect 109628 78562 109702 78686
rect 109826 78562 109870 78686
rect 109994 78562 110068 78686
rect 109628 77174 110068 78562
rect 109628 77050 109702 77174
rect 109826 77050 109870 77174
rect 109994 77050 110068 77174
rect 109628 75662 110068 77050
rect 109628 75538 109702 75662
rect 109826 75538 109870 75662
rect 109994 75538 110068 75662
rect 94508 70186 94538 70566
rect 94918 70186 94948 70566
rect 94508 70174 94948 70186
rect 94508 69794 94538 70174
rect 94918 69794 94948 70174
rect 94508 69782 94948 69794
rect 94508 69402 94538 69782
rect 94918 69402 94948 69782
rect 94508 69390 94948 69402
rect 94508 69010 94538 69390
rect 94918 69010 94948 69390
rect 94508 68998 94948 69010
rect 94508 68618 94538 68998
rect 94918 68618 94948 68998
rect 94508 68606 94948 68618
rect 94508 68226 94538 68606
rect 94918 68226 94948 68606
rect 94508 68214 94948 68226
rect 94508 67834 94538 68214
rect 94918 67834 94948 68214
rect 94508 67700 94948 67834
rect 109628 70566 110068 75538
rect 123508 151942 123948 152076
rect 123508 151562 123538 151942
rect 123918 151562 123948 151942
rect 123508 151550 123948 151562
rect 123508 151170 123538 151550
rect 123918 151170 123948 151550
rect 123508 151158 123948 151170
rect 123508 150778 123538 151158
rect 123918 150778 123948 151158
rect 123508 150766 123948 150778
rect 123508 150386 123538 150766
rect 123918 150386 123948 150766
rect 123508 150374 123948 150386
rect 123508 149994 123538 150374
rect 123918 149994 123948 150374
rect 123508 149982 123948 149994
rect 123508 149602 123538 149982
rect 123918 149602 123948 149982
rect 123508 149590 123948 149602
rect 123508 149210 123538 149590
rect 123918 149210 123948 149590
rect 123508 147482 123948 149210
rect 123508 147358 123582 147482
rect 123706 147358 123750 147482
rect 123874 147358 123948 147482
rect 123508 145970 123948 147358
rect 123508 145846 123582 145970
rect 123706 145846 123750 145970
rect 123874 145846 123948 145970
rect 123508 144458 123948 145846
rect 123508 144334 123582 144458
rect 123706 144334 123750 144458
rect 123874 144334 123948 144458
rect 123508 142946 123948 144334
rect 123508 142822 123582 142946
rect 123706 142822 123750 142946
rect 123874 142822 123948 142946
rect 123508 141434 123948 142822
rect 123508 141310 123582 141434
rect 123706 141310 123750 141434
rect 123874 141310 123948 141434
rect 123508 139922 123948 141310
rect 123508 139798 123582 139922
rect 123706 139798 123750 139922
rect 123874 139798 123948 139922
rect 123508 138990 123948 139798
rect 123508 138610 123538 138990
rect 123918 138610 123948 138990
rect 123508 138410 123948 138610
rect 123508 138286 123582 138410
rect 123706 138286 123750 138410
rect 123874 138286 123948 138410
rect 123508 136898 123948 138286
rect 123508 136774 123582 136898
rect 123706 136774 123750 136898
rect 123874 136774 123948 136898
rect 123508 135386 123948 136774
rect 123508 135262 123582 135386
rect 123706 135262 123750 135386
rect 123874 135262 123948 135386
rect 123508 133874 123948 135262
rect 123508 133750 123582 133874
rect 123706 133750 123750 133874
rect 123874 133750 123948 133874
rect 123508 132362 123948 133750
rect 123508 132238 123582 132362
rect 123706 132238 123750 132362
rect 123874 132238 123948 132362
rect 123508 130850 123948 132238
rect 123508 130726 123582 130850
rect 123706 130726 123750 130850
rect 123874 130726 123948 130850
rect 123508 129338 123948 130726
rect 123508 129214 123582 129338
rect 123706 129214 123750 129338
rect 123874 129214 123948 129338
rect 123508 127826 123948 129214
rect 123508 127702 123582 127826
rect 123706 127702 123750 127826
rect 123874 127702 123948 127826
rect 123508 126314 123948 127702
rect 123508 126190 123582 126314
rect 123706 126190 123750 126314
rect 123874 126190 123948 126314
rect 123508 124802 123948 126190
rect 123508 124678 123582 124802
rect 123706 124678 123750 124802
rect 123874 124678 123948 124802
rect 123508 123870 123948 124678
rect 123508 123490 123538 123870
rect 123918 123490 123948 123870
rect 123508 123290 123948 123490
rect 123508 123166 123582 123290
rect 123706 123166 123750 123290
rect 123874 123166 123948 123290
rect 123508 121778 123948 123166
rect 123508 121654 123582 121778
rect 123706 121654 123750 121778
rect 123874 121654 123948 121778
rect 123508 120266 123948 121654
rect 123508 120142 123582 120266
rect 123706 120142 123750 120266
rect 123874 120142 123948 120266
rect 123508 118754 123948 120142
rect 123508 118630 123582 118754
rect 123706 118630 123750 118754
rect 123874 118630 123948 118754
rect 123508 117242 123948 118630
rect 123508 117118 123582 117242
rect 123706 117118 123750 117242
rect 123874 117118 123948 117242
rect 123508 115730 123948 117118
rect 123508 115606 123582 115730
rect 123706 115606 123750 115730
rect 123874 115606 123948 115730
rect 123508 114218 123948 115606
rect 123508 114094 123582 114218
rect 123706 114094 123750 114218
rect 123874 114094 123948 114218
rect 123508 112706 123948 114094
rect 123508 112582 123582 112706
rect 123706 112582 123750 112706
rect 123874 112582 123948 112706
rect 123508 111194 123948 112582
rect 123508 111070 123582 111194
rect 123706 111070 123750 111194
rect 123874 111070 123948 111194
rect 123508 109682 123948 111070
rect 123508 109558 123582 109682
rect 123706 109558 123750 109682
rect 123874 109558 123948 109682
rect 123508 108750 123948 109558
rect 123508 108370 123538 108750
rect 123918 108370 123948 108750
rect 123508 108170 123948 108370
rect 123508 108046 123582 108170
rect 123706 108046 123750 108170
rect 123874 108046 123948 108170
rect 123508 106658 123948 108046
rect 123508 106534 123582 106658
rect 123706 106534 123750 106658
rect 123874 106534 123948 106658
rect 123508 105146 123948 106534
rect 123508 105022 123582 105146
rect 123706 105022 123750 105146
rect 123874 105022 123948 105146
rect 123508 103634 123948 105022
rect 123508 103510 123582 103634
rect 123706 103510 123750 103634
rect 123874 103510 123948 103634
rect 123508 102122 123948 103510
rect 123508 101998 123582 102122
rect 123706 101998 123750 102122
rect 123874 101998 123948 102122
rect 123508 100610 123948 101998
rect 123508 100486 123582 100610
rect 123706 100486 123750 100610
rect 123874 100486 123948 100610
rect 123508 99098 123948 100486
rect 123508 98974 123582 99098
rect 123706 98974 123750 99098
rect 123874 98974 123948 99098
rect 123508 97586 123948 98974
rect 123508 97462 123582 97586
rect 123706 97462 123750 97586
rect 123874 97462 123948 97586
rect 123508 96074 123948 97462
rect 123508 95950 123582 96074
rect 123706 95950 123750 96074
rect 123874 95950 123948 96074
rect 123508 94562 123948 95950
rect 123508 94438 123582 94562
rect 123706 94438 123750 94562
rect 123874 94438 123948 94562
rect 123508 93630 123948 94438
rect 123508 93250 123538 93630
rect 123918 93250 123948 93630
rect 123508 93050 123948 93250
rect 123508 92926 123582 93050
rect 123706 92926 123750 93050
rect 123874 92926 123948 93050
rect 123508 91538 123948 92926
rect 123508 91414 123582 91538
rect 123706 91414 123750 91538
rect 123874 91414 123948 91538
rect 123508 90026 123948 91414
rect 123508 89902 123582 90026
rect 123706 89902 123750 90026
rect 123874 89902 123948 90026
rect 123508 88514 123948 89902
rect 123508 88390 123582 88514
rect 123706 88390 123750 88514
rect 123874 88390 123948 88514
rect 123508 87002 123948 88390
rect 123508 86878 123582 87002
rect 123706 86878 123750 87002
rect 123874 86878 123948 87002
rect 123508 85490 123948 86878
rect 123508 85366 123582 85490
rect 123706 85366 123750 85490
rect 123874 85366 123948 85490
rect 123508 83978 123948 85366
rect 123508 83854 123582 83978
rect 123706 83854 123750 83978
rect 123874 83854 123948 83978
rect 123508 82466 123948 83854
rect 123508 82342 123582 82466
rect 123706 82342 123750 82466
rect 123874 82342 123948 82466
rect 123508 80954 123948 82342
rect 123508 80830 123582 80954
rect 123706 80830 123750 80954
rect 123874 80830 123948 80954
rect 123508 79442 123948 80830
rect 123508 79318 123582 79442
rect 123706 79318 123750 79442
rect 123874 79318 123948 79442
rect 123508 78510 123948 79318
rect 123508 78130 123538 78510
rect 123918 78130 123948 78510
rect 123508 77930 123948 78130
rect 123508 77806 123582 77930
rect 123706 77806 123750 77930
rect 123874 77806 123948 77930
rect 123508 76418 123948 77806
rect 123508 76294 123582 76418
rect 123706 76294 123750 76418
rect 123874 76294 123948 76418
rect 123508 74566 123948 76294
rect 123508 74186 123538 74566
rect 123918 74186 123948 74566
rect 123508 74174 123948 74186
rect 123508 73794 123538 74174
rect 123918 73794 123948 74174
rect 123508 73782 123948 73794
rect 123508 73402 123538 73782
rect 123918 73402 123948 73782
rect 123508 73390 123948 73402
rect 123508 73010 123538 73390
rect 123918 73010 123948 73390
rect 123508 72998 123948 73010
rect 123508 72618 123538 72998
rect 123918 72618 123948 72998
rect 123508 72606 123948 72618
rect 123508 72226 123538 72606
rect 123918 72226 123948 72606
rect 123508 72214 123948 72226
rect 123508 71834 123538 72214
rect 123918 71834 123948 72214
rect 123508 71700 123948 71834
rect 124748 148238 125188 153210
rect 139868 155942 140308 156076
rect 139868 155562 139898 155942
rect 140278 155562 140308 155942
rect 139868 155550 140308 155562
rect 139868 155170 139898 155550
rect 140278 155170 140308 155550
rect 139868 155158 140308 155170
rect 139868 154778 139898 155158
rect 140278 154778 140308 155158
rect 139868 154766 140308 154778
rect 139868 154386 139898 154766
rect 140278 154386 140308 154766
rect 139868 154374 140308 154386
rect 139868 153994 139898 154374
rect 140278 153994 140308 154374
rect 139868 153982 140308 153994
rect 139868 153602 139898 153982
rect 140278 153602 140308 153982
rect 139868 153590 140308 153602
rect 139868 153210 139898 153590
rect 140278 153210 140308 153590
rect 124748 148114 124822 148238
rect 124946 148114 124990 148238
rect 125114 148114 125188 148238
rect 124748 146726 125188 148114
rect 124748 146602 124822 146726
rect 124946 146602 124990 146726
rect 125114 146602 125188 146726
rect 124748 145214 125188 146602
rect 124748 145090 124822 145214
rect 124946 145090 124990 145214
rect 125114 145090 125188 145214
rect 124748 143702 125188 145090
rect 124748 143578 124822 143702
rect 124946 143578 124990 143702
rect 125114 143578 125188 143702
rect 124748 142190 125188 143578
rect 124748 142066 124822 142190
rect 124946 142066 124990 142190
rect 125114 142066 125188 142190
rect 124748 140678 125188 142066
rect 124748 140554 124822 140678
rect 124946 140554 124990 140678
rect 125114 140554 125188 140678
rect 124748 140230 125188 140554
rect 124748 139850 124778 140230
rect 125158 139850 125188 140230
rect 124748 139166 125188 139850
rect 124748 139042 124822 139166
rect 124946 139042 124990 139166
rect 125114 139042 125188 139166
rect 124748 137654 125188 139042
rect 124748 137530 124822 137654
rect 124946 137530 124990 137654
rect 125114 137530 125188 137654
rect 124748 136142 125188 137530
rect 124748 136018 124822 136142
rect 124946 136018 124990 136142
rect 125114 136018 125188 136142
rect 124748 134630 125188 136018
rect 124748 134506 124822 134630
rect 124946 134506 124990 134630
rect 125114 134506 125188 134630
rect 124748 133118 125188 134506
rect 124748 132994 124822 133118
rect 124946 132994 124990 133118
rect 125114 132994 125188 133118
rect 124748 131606 125188 132994
rect 124748 131482 124822 131606
rect 124946 131482 124990 131606
rect 125114 131482 125188 131606
rect 124748 130094 125188 131482
rect 124748 129970 124822 130094
rect 124946 129970 124990 130094
rect 125114 129970 125188 130094
rect 124748 128582 125188 129970
rect 124748 128458 124822 128582
rect 124946 128458 124990 128582
rect 125114 128458 125188 128582
rect 124748 127070 125188 128458
rect 124748 126946 124822 127070
rect 124946 126946 124990 127070
rect 125114 126946 125188 127070
rect 124748 125558 125188 126946
rect 124748 125434 124822 125558
rect 124946 125434 124990 125558
rect 125114 125434 125188 125558
rect 124748 125110 125188 125434
rect 124748 124730 124778 125110
rect 125158 124730 125188 125110
rect 124748 124046 125188 124730
rect 124748 123922 124822 124046
rect 124946 123922 124990 124046
rect 125114 123922 125188 124046
rect 124748 122534 125188 123922
rect 124748 122410 124822 122534
rect 124946 122410 124990 122534
rect 125114 122410 125188 122534
rect 124748 121022 125188 122410
rect 124748 120898 124822 121022
rect 124946 120898 124990 121022
rect 125114 120898 125188 121022
rect 124748 119510 125188 120898
rect 124748 119386 124822 119510
rect 124946 119386 124990 119510
rect 125114 119386 125188 119510
rect 124748 117998 125188 119386
rect 124748 117874 124822 117998
rect 124946 117874 124990 117998
rect 125114 117874 125188 117998
rect 124748 116486 125188 117874
rect 124748 116362 124822 116486
rect 124946 116362 124990 116486
rect 125114 116362 125188 116486
rect 124748 114974 125188 116362
rect 124748 114850 124822 114974
rect 124946 114850 124990 114974
rect 125114 114850 125188 114974
rect 124748 113462 125188 114850
rect 124748 113338 124822 113462
rect 124946 113338 124990 113462
rect 125114 113338 125188 113462
rect 124748 111950 125188 113338
rect 124748 111826 124822 111950
rect 124946 111826 124990 111950
rect 125114 111826 125188 111950
rect 124748 110438 125188 111826
rect 124748 110314 124822 110438
rect 124946 110314 124990 110438
rect 125114 110314 125188 110438
rect 124748 109990 125188 110314
rect 124748 109610 124778 109990
rect 125158 109610 125188 109990
rect 124748 108926 125188 109610
rect 124748 108802 124822 108926
rect 124946 108802 124990 108926
rect 125114 108802 125188 108926
rect 124748 107414 125188 108802
rect 124748 107290 124822 107414
rect 124946 107290 124990 107414
rect 125114 107290 125188 107414
rect 124748 105902 125188 107290
rect 124748 105778 124822 105902
rect 124946 105778 124990 105902
rect 125114 105778 125188 105902
rect 124748 104390 125188 105778
rect 124748 104266 124822 104390
rect 124946 104266 124990 104390
rect 125114 104266 125188 104390
rect 124748 102878 125188 104266
rect 124748 102754 124822 102878
rect 124946 102754 124990 102878
rect 125114 102754 125188 102878
rect 124748 101366 125188 102754
rect 124748 101242 124822 101366
rect 124946 101242 124990 101366
rect 125114 101242 125188 101366
rect 124748 99854 125188 101242
rect 124748 99730 124822 99854
rect 124946 99730 124990 99854
rect 125114 99730 125188 99854
rect 124748 98342 125188 99730
rect 124748 98218 124822 98342
rect 124946 98218 124990 98342
rect 125114 98218 125188 98342
rect 124748 96830 125188 98218
rect 124748 96706 124822 96830
rect 124946 96706 124990 96830
rect 125114 96706 125188 96830
rect 124748 95318 125188 96706
rect 124748 95194 124822 95318
rect 124946 95194 124990 95318
rect 125114 95194 125188 95318
rect 124748 94870 125188 95194
rect 124748 94490 124778 94870
rect 125158 94490 125188 94870
rect 124748 93806 125188 94490
rect 124748 93682 124822 93806
rect 124946 93682 124990 93806
rect 125114 93682 125188 93806
rect 124748 92294 125188 93682
rect 124748 92170 124822 92294
rect 124946 92170 124990 92294
rect 125114 92170 125188 92294
rect 124748 90782 125188 92170
rect 124748 90658 124822 90782
rect 124946 90658 124990 90782
rect 125114 90658 125188 90782
rect 124748 89270 125188 90658
rect 124748 89146 124822 89270
rect 124946 89146 124990 89270
rect 125114 89146 125188 89270
rect 124748 87758 125188 89146
rect 124748 87634 124822 87758
rect 124946 87634 124990 87758
rect 125114 87634 125188 87758
rect 124748 86246 125188 87634
rect 124748 86122 124822 86246
rect 124946 86122 124990 86246
rect 125114 86122 125188 86246
rect 124748 84734 125188 86122
rect 124748 84610 124822 84734
rect 124946 84610 124990 84734
rect 125114 84610 125188 84734
rect 124748 83222 125188 84610
rect 124748 83098 124822 83222
rect 124946 83098 124990 83222
rect 125114 83098 125188 83222
rect 124748 81710 125188 83098
rect 124748 81586 124822 81710
rect 124946 81586 124990 81710
rect 125114 81586 125188 81710
rect 124748 80198 125188 81586
rect 124748 80074 124822 80198
rect 124946 80074 124990 80198
rect 125114 80074 125188 80198
rect 124748 79750 125188 80074
rect 124748 79370 124778 79750
rect 125158 79370 125188 79750
rect 124748 78686 125188 79370
rect 124748 78562 124822 78686
rect 124946 78562 124990 78686
rect 125114 78562 125188 78686
rect 124748 77174 125188 78562
rect 124748 77050 124822 77174
rect 124946 77050 124990 77174
rect 125114 77050 125188 77174
rect 124748 75662 125188 77050
rect 124748 75538 124822 75662
rect 124946 75538 124990 75662
rect 125114 75538 125188 75662
rect 109628 70186 109658 70566
rect 110038 70186 110068 70566
rect 109628 70174 110068 70186
rect 109628 69794 109658 70174
rect 110038 69794 110068 70174
rect 109628 69782 110068 69794
rect 109628 69402 109658 69782
rect 110038 69402 110068 69782
rect 109628 69390 110068 69402
rect 109628 69010 109658 69390
rect 110038 69010 110068 69390
rect 109628 68998 110068 69010
rect 109628 68618 109658 68998
rect 110038 68618 110068 68998
rect 109628 68606 110068 68618
rect 109628 68226 109658 68606
rect 110038 68226 110068 68606
rect 109628 68214 110068 68226
rect 109628 67834 109658 68214
rect 110038 67834 110068 68214
rect 109628 67700 110068 67834
rect 124748 70566 125188 75538
rect 138628 151942 139068 152076
rect 138628 151562 138658 151942
rect 139038 151562 139068 151942
rect 138628 151550 139068 151562
rect 138628 151170 138658 151550
rect 139038 151170 139068 151550
rect 138628 151158 139068 151170
rect 138628 150778 138658 151158
rect 139038 150778 139068 151158
rect 138628 150766 139068 150778
rect 138628 150386 138658 150766
rect 139038 150386 139068 150766
rect 138628 150374 139068 150386
rect 138628 149994 138658 150374
rect 139038 149994 139068 150374
rect 138628 149982 139068 149994
rect 138628 149602 138658 149982
rect 139038 149602 139068 149982
rect 138628 149590 139068 149602
rect 138628 149210 138658 149590
rect 139038 149210 139068 149590
rect 138628 147482 139068 149210
rect 138628 147358 138702 147482
rect 138826 147358 138870 147482
rect 138994 147358 139068 147482
rect 138628 145970 139068 147358
rect 138628 145846 138702 145970
rect 138826 145846 138870 145970
rect 138994 145846 139068 145970
rect 138628 144458 139068 145846
rect 138628 144334 138702 144458
rect 138826 144334 138870 144458
rect 138994 144334 139068 144458
rect 138628 142946 139068 144334
rect 138628 142822 138702 142946
rect 138826 142822 138870 142946
rect 138994 142822 139068 142946
rect 138628 141434 139068 142822
rect 138628 141310 138702 141434
rect 138826 141310 138870 141434
rect 138994 141310 139068 141434
rect 138628 139922 139068 141310
rect 138628 139798 138702 139922
rect 138826 139798 138870 139922
rect 138994 139798 139068 139922
rect 138628 138990 139068 139798
rect 138628 138610 138658 138990
rect 139038 138610 139068 138990
rect 138628 138410 139068 138610
rect 138628 138286 138702 138410
rect 138826 138286 138870 138410
rect 138994 138286 139068 138410
rect 138628 136898 139068 138286
rect 138628 136774 138702 136898
rect 138826 136774 138870 136898
rect 138994 136774 139068 136898
rect 138628 135386 139068 136774
rect 138628 135262 138702 135386
rect 138826 135262 138870 135386
rect 138994 135262 139068 135386
rect 138628 133874 139068 135262
rect 138628 133750 138702 133874
rect 138826 133750 138870 133874
rect 138994 133750 139068 133874
rect 138628 132362 139068 133750
rect 138628 132238 138702 132362
rect 138826 132238 138870 132362
rect 138994 132238 139068 132362
rect 138628 130850 139068 132238
rect 138628 130726 138702 130850
rect 138826 130726 138870 130850
rect 138994 130726 139068 130850
rect 138628 129338 139068 130726
rect 138628 129214 138702 129338
rect 138826 129214 138870 129338
rect 138994 129214 139068 129338
rect 138628 127826 139068 129214
rect 138628 127702 138702 127826
rect 138826 127702 138870 127826
rect 138994 127702 139068 127826
rect 138628 126314 139068 127702
rect 138628 126190 138702 126314
rect 138826 126190 138870 126314
rect 138994 126190 139068 126314
rect 138628 124802 139068 126190
rect 138628 124678 138702 124802
rect 138826 124678 138870 124802
rect 138994 124678 139068 124802
rect 138628 123870 139068 124678
rect 138628 123490 138658 123870
rect 139038 123490 139068 123870
rect 138628 123290 139068 123490
rect 138628 123166 138702 123290
rect 138826 123166 138870 123290
rect 138994 123166 139068 123290
rect 138628 121778 139068 123166
rect 138628 121654 138702 121778
rect 138826 121654 138870 121778
rect 138994 121654 139068 121778
rect 138628 120266 139068 121654
rect 138628 120142 138702 120266
rect 138826 120142 138870 120266
rect 138994 120142 139068 120266
rect 138628 118754 139068 120142
rect 138628 118630 138702 118754
rect 138826 118630 138870 118754
rect 138994 118630 139068 118754
rect 138628 117242 139068 118630
rect 138628 117118 138702 117242
rect 138826 117118 138870 117242
rect 138994 117118 139068 117242
rect 138628 115730 139068 117118
rect 138628 115606 138702 115730
rect 138826 115606 138870 115730
rect 138994 115606 139068 115730
rect 138628 114218 139068 115606
rect 138628 114094 138702 114218
rect 138826 114094 138870 114218
rect 138994 114094 139068 114218
rect 138628 112706 139068 114094
rect 138628 112582 138702 112706
rect 138826 112582 138870 112706
rect 138994 112582 139068 112706
rect 138628 111194 139068 112582
rect 138628 111070 138702 111194
rect 138826 111070 138870 111194
rect 138994 111070 139068 111194
rect 138628 109682 139068 111070
rect 138628 109558 138702 109682
rect 138826 109558 138870 109682
rect 138994 109558 139068 109682
rect 138628 108750 139068 109558
rect 138628 108370 138658 108750
rect 139038 108370 139068 108750
rect 138628 108170 139068 108370
rect 138628 108046 138702 108170
rect 138826 108046 138870 108170
rect 138994 108046 139068 108170
rect 138628 106658 139068 108046
rect 138628 106534 138702 106658
rect 138826 106534 138870 106658
rect 138994 106534 139068 106658
rect 138628 105146 139068 106534
rect 138628 105022 138702 105146
rect 138826 105022 138870 105146
rect 138994 105022 139068 105146
rect 138628 103634 139068 105022
rect 138628 103510 138702 103634
rect 138826 103510 138870 103634
rect 138994 103510 139068 103634
rect 138628 102122 139068 103510
rect 138628 101998 138702 102122
rect 138826 101998 138870 102122
rect 138994 101998 139068 102122
rect 138628 100610 139068 101998
rect 138628 100486 138702 100610
rect 138826 100486 138870 100610
rect 138994 100486 139068 100610
rect 138628 99098 139068 100486
rect 138628 98974 138702 99098
rect 138826 98974 138870 99098
rect 138994 98974 139068 99098
rect 138628 97586 139068 98974
rect 138628 97462 138702 97586
rect 138826 97462 138870 97586
rect 138994 97462 139068 97586
rect 138628 96074 139068 97462
rect 138628 95950 138702 96074
rect 138826 95950 138870 96074
rect 138994 95950 139068 96074
rect 138628 94562 139068 95950
rect 138628 94438 138702 94562
rect 138826 94438 138870 94562
rect 138994 94438 139068 94562
rect 138628 93630 139068 94438
rect 138628 93250 138658 93630
rect 139038 93250 139068 93630
rect 138628 93050 139068 93250
rect 138628 92926 138702 93050
rect 138826 92926 138870 93050
rect 138994 92926 139068 93050
rect 138628 91538 139068 92926
rect 138628 91414 138702 91538
rect 138826 91414 138870 91538
rect 138994 91414 139068 91538
rect 138628 90026 139068 91414
rect 138628 89902 138702 90026
rect 138826 89902 138870 90026
rect 138994 89902 139068 90026
rect 138628 88514 139068 89902
rect 138628 88390 138702 88514
rect 138826 88390 138870 88514
rect 138994 88390 139068 88514
rect 138628 87002 139068 88390
rect 138628 86878 138702 87002
rect 138826 86878 138870 87002
rect 138994 86878 139068 87002
rect 138628 85490 139068 86878
rect 138628 85366 138702 85490
rect 138826 85366 138870 85490
rect 138994 85366 139068 85490
rect 138628 83978 139068 85366
rect 138628 83854 138702 83978
rect 138826 83854 138870 83978
rect 138994 83854 139068 83978
rect 138628 82466 139068 83854
rect 138628 82342 138702 82466
rect 138826 82342 138870 82466
rect 138994 82342 139068 82466
rect 138628 80954 139068 82342
rect 138628 80830 138702 80954
rect 138826 80830 138870 80954
rect 138994 80830 139068 80954
rect 138628 79442 139068 80830
rect 138628 79318 138702 79442
rect 138826 79318 138870 79442
rect 138994 79318 139068 79442
rect 138628 78510 139068 79318
rect 138628 78130 138658 78510
rect 139038 78130 139068 78510
rect 138628 77930 139068 78130
rect 138628 77806 138702 77930
rect 138826 77806 138870 77930
rect 138994 77806 139068 77930
rect 138628 76418 139068 77806
rect 138628 76294 138702 76418
rect 138826 76294 138870 76418
rect 138994 76294 139068 76418
rect 138628 74566 139068 76294
rect 138628 74186 138658 74566
rect 139038 74186 139068 74566
rect 138628 74174 139068 74186
rect 138628 73794 138658 74174
rect 139038 73794 139068 74174
rect 138628 73782 139068 73794
rect 138628 73402 138658 73782
rect 139038 73402 139068 73782
rect 138628 73390 139068 73402
rect 138628 73010 138658 73390
rect 139038 73010 139068 73390
rect 138628 72998 139068 73010
rect 138628 72618 138658 72998
rect 139038 72618 139068 72998
rect 138628 72606 139068 72618
rect 138628 72226 138658 72606
rect 139038 72226 139068 72606
rect 138628 72214 139068 72226
rect 138628 71834 138658 72214
rect 139038 71834 139068 72214
rect 138628 71700 139068 71834
rect 139868 148238 140308 153210
rect 153220 155942 156220 156076
rect 153220 155562 153354 155942
rect 153734 155562 153746 155942
rect 154126 155562 154138 155942
rect 154518 155562 154530 155942
rect 154910 155562 154922 155942
rect 155302 155562 155314 155942
rect 155694 155562 155706 155942
rect 156086 155562 156220 155942
rect 153220 155550 156220 155562
rect 153220 155170 153354 155550
rect 153734 155170 153746 155550
rect 154126 155170 154138 155550
rect 154518 155170 154530 155550
rect 154910 155170 154922 155550
rect 155302 155170 155314 155550
rect 155694 155170 155706 155550
rect 156086 155170 156220 155550
rect 153220 155158 156220 155170
rect 153220 154778 153354 155158
rect 153734 154778 153746 155158
rect 154126 154778 154138 155158
rect 154518 154778 154530 155158
rect 154910 154778 154922 155158
rect 155302 154778 155314 155158
rect 155694 154778 155706 155158
rect 156086 154778 156220 155158
rect 153220 154766 156220 154778
rect 153220 154386 153354 154766
rect 153734 154386 153746 154766
rect 154126 154386 154138 154766
rect 154518 154386 154530 154766
rect 154910 154386 154922 154766
rect 155302 154386 155314 154766
rect 155694 154386 155706 154766
rect 156086 154386 156220 154766
rect 153220 154374 156220 154386
rect 153220 153994 153354 154374
rect 153734 153994 153746 154374
rect 154126 153994 154138 154374
rect 154518 153994 154530 154374
rect 154910 153994 154922 154374
rect 155302 153994 155314 154374
rect 155694 153994 155706 154374
rect 156086 153994 156220 154374
rect 153220 153982 156220 153994
rect 153220 153602 153354 153982
rect 153734 153602 153746 153982
rect 154126 153602 154138 153982
rect 154518 153602 154530 153982
rect 154910 153602 154922 153982
rect 155302 153602 155314 153982
rect 155694 153602 155706 153982
rect 156086 153602 156220 153982
rect 153220 153590 156220 153602
rect 153220 153210 153354 153590
rect 153734 153210 153746 153590
rect 154126 153210 154138 153590
rect 154518 153210 154530 153590
rect 154910 153210 154922 153590
rect 155302 153210 155314 153590
rect 155694 153210 155706 153590
rect 156086 153210 156220 153590
rect 139868 148114 139942 148238
rect 140066 148114 140110 148238
rect 140234 148114 140308 148238
rect 139868 146726 140308 148114
rect 139868 146602 139942 146726
rect 140066 146602 140110 146726
rect 140234 146602 140308 146726
rect 139868 145214 140308 146602
rect 139868 145090 139942 145214
rect 140066 145090 140110 145214
rect 140234 145090 140308 145214
rect 139868 143702 140308 145090
rect 139868 143578 139942 143702
rect 140066 143578 140110 143702
rect 140234 143578 140308 143702
rect 139868 142190 140308 143578
rect 139868 142066 139942 142190
rect 140066 142066 140110 142190
rect 140234 142066 140308 142190
rect 139868 140678 140308 142066
rect 139868 140554 139942 140678
rect 140066 140554 140110 140678
rect 140234 140554 140308 140678
rect 139868 140230 140308 140554
rect 139868 139850 139898 140230
rect 140278 139850 140308 140230
rect 139868 139166 140308 139850
rect 139868 139042 139942 139166
rect 140066 139042 140110 139166
rect 140234 139042 140308 139166
rect 139868 137654 140308 139042
rect 139868 137530 139942 137654
rect 140066 137530 140110 137654
rect 140234 137530 140308 137654
rect 139868 136142 140308 137530
rect 139868 136018 139942 136142
rect 140066 136018 140110 136142
rect 140234 136018 140308 136142
rect 139868 134630 140308 136018
rect 139868 134506 139942 134630
rect 140066 134506 140110 134630
rect 140234 134506 140308 134630
rect 139868 133118 140308 134506
rect 139868 132994 139942 133118
rect 140066 132994 140110 133118
rect 140234 132994 140308 133118
rect 139868 131606 140308 132994
rect 139868 131482 139942 131606
rect 140066 131482 140110 131606
rect 140234 131482 140308 131606
rect 139868 130094 140308 131482
rect 139868 129970 139942 130094
rect 140066 129970 140110 130094
rect 140234 129970 140308 130094
rect 139868 128582 140308 129970
rect 139868 128458 139942 128582
rect 140066 128458 140110 128582
rect 140234 128458 140308 128582
rect 139868 127070 140308 128458
rect 139868 126946 139942 127070
rect 140066 126946 140110 127070
rect 140234 126946 140308 127070
rect 139868 125558 140308 126946
rect 139868 125434 139942 125558
rect 140066 125434 140110 125558
rect 140234 125434 140308 125558
rect 139868 125110 140308 125434
rect 139868 124730 139898 125110
rect 140278 124730 140308 125110
rect 139868 124046 140308 124730
rect 139868 123922 139942 124046
rect 140066 123922 140110 124046
rect 140234 123922 140308 124046
rect 139868 122534 140308 123922
rect 139868 122410 139942 122534
rect 140066 122410 140110 122534
rect 140234 122410 140308 122534
rect 139868 121022 140308 122410
rect 139868 120898 139942 121022
rect 140066 120898 140110 121022
rect 140234 120898 140308 121022
rect 139868 119510 140308 120898
rect 139868 119386 139942 119510
rect 140066 119386 140110 119510
rect 140234 119386 140308 119510
rect 139868 117998 140308 119386
rect 139868 117874 139942 117998
rect 140066 117874 140110 117998
rect 140234 117874 140308 117998
rect 139868 116486 140308 117874
rect 139868 116362 139942 116486
rect 140066 116362 140110 116486
rect 140234 116362 140308 116486
rect 139868 114974 140308 116362
rect 139868 114850 139942 114974
rect 140066 114850 140110 114974
rect 140234 114850 140308 114974
rect 139868 113462 140308 114850
rect 139868 113338 139942 113462
rect 140066 113338 140110 113462
rect 140234 113338 140308 113462
rect 139868 111950 140308 113338
rect 139868 111826 139942 111950
rect 140066 111826 140110 111950
rect 140234 111826 140308 111950
rect 139868 110438 140308 111826
rect 139868 110314 139942 110438
rect 140066 110314 140110 110438
rect 140234 110314 140308 110438
rect 139868 109990 140308 110314
rect 139868 109610 139898 109990
rect 140278 109610 140308 109990
rect 139868 108926 140308 109610
rect 139868 108802 139942 108926
rect 140066 108802 140110 108926
rect 140234 108802 140308 108926
rect 139868 107414 140308 108802
rect 139868 107290 139942 107414
rect 140066 107290 140110 107414
rect 140234 107290 140308 107414
rect 139868 105902 140308 107290
rect 139868 105778 139942 105902
rect 140066 105778 140110 105902
rect 140234 105778 140308 105902
rect 139868 104390 140308 105778
rect 139868 104266 139942 104390
rect 140066 104266 140110 104390
rect 140234 104266 140308 104390
rect 139868 102878 140308 104266
rect 139868 102754 139942 102878
rect 140066 102754 140110 102878
rect 140234 102754 140308 102878
rect 139868 101366 140308 102754
rect 139868 101242 139942 101366
rect 140066 101242 140110 101366
rect 140234 101242 140308 101366
rect 139868 99854 140308 101242
rect 139868 99730 139942 99854
rect 140066 99730 140110 99854
rect 140234 99730 140308 99854
rect 139868 98342 140308 99730
rect 139868 98218 139942 98342
rect 140066 98218 140110 98342
rect 140234 98218 140308 98342
rect 139868 96830 140308 98218
rect 139868 96706 139942 96830
rect 140066 96706 140110 96830
rect 140234 96706 140308 96830
rect 139868 95318 140308 96706
rect 139868 95194 139942 95318
rect 140066 95194 140110 95318
rect 140234 95194 140308 95318
rect 139868 94870 140308 95194
rect 139868 94490 139898 94870
rect 140278 94490 140308 94870
rect 139868 93806 140308 94490
rect 139868 93682 139942 93806
rect 140066 93682 140110 93806
rect 140234 93682 140308 93806
rect 139868 92294 140308 93682
rect 139868 92170 139942 92294
rect 140066 92170 140110 92294
rect 140234 92170 140308 92294
rect 139868 90782 140308 92170
rect 139868 90658 139942 90782
rect 140066 90658 140110 90782
rect 140234 90658 140308 90782
rect 139868 89270 140308 90658
rect 139868 89146 139942 89270
rect 140066 89146 140110 89270
rect 140234 89146 140308 89270
rect 139868 87758 140308 89146
rect 139868 87634 139942 87758
rect 140066 87634 140110 87758
rect 140234 87634 140308 87758
rect 139868 86246 140308 87634
rect 139868 86122 139942 86246
rect 140066 86122 140110 86246
rect 140234 86122 140308 86246
rect 139868 84734 140308 86122
rect 139868 84610 139942 84734
rect 140066 84610 140110 84734
rect 140234 84610 140308 84734
rect 139868 83222 140308 84610
rect 139868 83098 139942 83222
rect 140066 83098 140110 83222
rect 140234 83098 140308 83222
rect 139868 81710 140308 83098
rect 139868 81586 139942 81710
rect 140066 81586 140110 81710
rect 140234 81586 140308 81710
rect 139868 80198 140308 81586
rect 139868 80074 139942 80198
rect 140066 80074 140110 80198
rect 140234 80074 140308 80198
rect 139868 79750 140308 80074
rect 139868 79370 139898 79750
rect 140278 79370 140308 79750
rect 139868 78686 140308 79370
rect 139868 78562 139942 78686
rect 140066 78562 140110 78686
rect 140234 78562 140308 78686
rect 139868 77174 140308 78562
rect 139868 77050 139942 77174
rect 140066 77050 140110 77174
rect 140234 77050 140308 77174
rect 139868 75662 140308 77050
rect 139868 75538 139942 75662
rect 140066 75538 140110 75662
rect 140234 75538 140308 75662
rect 124748 70186 124778 70566
rect 125158 70186 125188 70566
rect 124748 70174 125188 70186
rect 124748 69794 124778 70174
rect 125158 69794 125188 70174
rect 124748 69782 125188 69794
rect 124748 69402 124778 69782
rect 125158 69402 125188 69782
rect 124748 69390 125188 69402
rect 124748 69010 124778 69390
rect 125158 69010 125188 69390
rect 124748 68998 125188 69010
rect 124748 68618 124778 68998
rect 125158 68618 125188 68998
rect 124748 68606 125188 68618
rect 124748 68226 124778 68606
rect 125158 68226 125188 68606
rect 124748 68214 125188 68226
rect 124748 67834 124778 68214
rect 125158 67834 125188 68214
rect 124748 67700 125188 67834
rect 139868 70566 140308 75538
rect 149220 151942 152220 152076
rect 149220 151562 149354 151942
rect 149734 151562 149746 151942
rect 150126 151562 150138 151942
rect 150518 151562 150530 151942
rect 150910 151562 150922 151942
rect 151302 151562 151314 151942
rect 151694 151562 151706 151942
rect 152086 151562 152220 151942
rect 149220 151550 152220 151562
rect 149220 151170 149354 151550
rect 149734 151170 149746 151550
rect 150126 151170 150138 151550
rect 150518 151170 150530 151550
rect 150910 151170 150922 151550
rect 151302 151170 151314 151550
rect 151694 151170 151706 151550
rect 152086 151170 152220 151550
rect 149220 151158 152220 151170
rect 149220 150778 149354 151158
rect 149734 150778 149746 151158
rect 150126 150778 150138 151158
rect 150518 150778 150530 151158
rect 150910 150778 150922 151158
rect 151302 150778 151314 151158
rect 151694 150778 151706 151158
rect 152086 150778 152220 151158
rect 149220 150766 152220 150778
rect 149220 150386 149354 150766
rect 149734 150386 149746 150766
rect 150126 150386 150138 150766
rect 150518 150386 150530 150766
rect 150910 150386 150922 150766
rect 151302 150386 151314 150766
rect 151694 150386 151706 150766
rect 152086 150386 152220 150766
rect 149220 150374 152220 150386
rect 149220 149994 149354 150374
rect 149734 149994 149746 150374
rect 150126 149994 150138 150374
rect 150518 149994 150530 150374
rect 150910 149994 150922 150374
rect 151302 149994 151314 150374
rect 151694 149994 151706 150374
rect 152086 149994 152220 150374
rect 149220 149982 152220 149994
rect 149220 149602 149354 149982
rect 149734 149602 149746 149982
rect 150126 149602 150138 149982
rect 150518 149602 150530 149982
rect 150910 149602 150922 149982
rect 151302 149602 151314 149982
rect 151694 149602 151706 149982
rect 152086 149602 152220 149982
rect 149220 149590 152220 149602
rect 149220 149210 149354 149590
rect 149734 149210 149746 149590
rect 150126 149210 150138 149590
rect 150518 149210 150530 149590
rect 150910 149210 150922 149590
rect 151302 149210 151314 149590
rect 151694 149210 151706 149590
rect 152086 149210 152220 149590
rect 149220 138990 152220 149210
rect 149220 138610 149354 138990
rect 149734 138610 149746 138990
rect 150126 138610 150138 138990
rect 150518 138610 150530 138990
rect 150910 138610 150922 138990
rect 151302 138610 151314 138990
rect 151694 138610 151706 138990
rect 152086 138610 152220 138990
rect 149220 133169 152220 138610
rect 149220 132789 149354 133169
rect 149734 132789 149746 133169
rect 150126 132789 150138 133169
rect 150518 132789 150530 133169
rect 150910 132789 150922 133169
rect 151302 132789 151314 133169
rect 151694 132789 151706 133169
rect 152086 132789 152220 133169
rect 149220 132777 152220 132789
rect 149220 132397 149354 132777
rect 149734 132397 149746 132777
rect 150126 132397 150138 132777
rect 150518 132397 150530 132777
rect 150910 132397 150922 132777
rect 151302 132397 151314 132777
rect 151694 132397 151706 132777
rect 152086 132397 152220 132777
rect 149220 132385 152220 132397
rect 149220 132005 149354 132385
rect 149734 132005 149746 132385
rect 150126 132005 150138 132385
rect 150518 132005 150530 132385
rect 150910 132005 150922 132385
rect 151302 132005 151314 132385
rect 151694 132005 151706 132385
rect 152086 132005 152220 132385
rect 149220 131993 152220 132005
rect 149220 131613 149354 131993
rect 149734 131613 149746 131993
rect 150126 131613 150138 131993
rect 150518 131613 150530 131993
rect 150910 131613 150922 131993
rect 151302 131613 151314 131993
rect 151694 131613 151706 131993
rect 152086 131613 152220 131993
rect 149220 131601 152220 131613
rect 149220 131221 149354 131601
rect 149734 131221 149746 131601
rect 150126 131221 150138 131601
rect 150518 131221 150530 131601
rect 150910 131221 150922 131601
rect 151302 131221 151314 131601
rect 151694 131221 151706 131601
rect 152086 131221 152220 131601
rect 149220 131209 152220 131221
rect 149220 130829 149354 131209
rect 149734 130829 149746 131209
rect 150126 130829 150138 131209
rect 150518 130829 150530 131209
rect 150910 130829 150922 131209
rect 151302 130829 151314 131209
rect 151694 130829 151706 131209
rect 152086 130829 152220 131209
rect 149220 123870 152220 130829
rect 149220 123490 149354 123870
rect 149734 123490 149746 123870
rect 150126 123490 150138 123870
rect 150518 123490 150530 123870
rect 150910 123490 150922 123870
rect 151302 123490 151314 123870
rect 151694 123490 151706 123870
rect 152086 123490 152220 123870
rect 149220 117169 152220 123490
rect 149220 116789 149354 117169
rect 149734 116789 149746 117169
rect 150126 116789 150138 117169
rect 150518 116789 150530 117169
rect 150910 116789 150922 117169
rect 151302 116789 151314 117169
rect 151694 116789 151706 117169
rect 152086 116789 152220 117169
rect 149220 116777 152220 116789
rect 149220 116397 149354 116777
rect 149734 116397 149746 116777
rect 150126 116397 150138 116777
rect 150518 116397 150530 116777
rect 150910 116397 150922 116777
rect 151302 116397 151314 116777
rect 151694 116397 151706 116777
rect 152086 116397 152220 116777
rect 149220 116385 152220 116397
rect 149220 116005 149354 116385
rect 149734 116005 149746 116385
rect 150126 116005 150138 116385
rect 150518 116005 150530 116385
rect 150910 116005 150922 116385
rect 151302 116005 151314 116385
rect 151694 116005 151706 116385
rect 152086 116005 152220 116385
rect 149220 115993 152220 116005
rect 149220 115613 149354 115993
rect 149734 115613 149746 115993
rect 150126 115613 150138 115993
rect 150518 115613 150530 115993
rect 150910 115613 150922 115993
rect 151302 115613 151314 115993
rect 151694 115613 151706 115993
rect 152086 115613 152220 115993
rect 149220 115601 152220 115613
rect 149220 115221 149354 115601
rect 149734 115221 149746 115601
rect 150126 115221 150138 115601
rect 150518 115221 150530 115601
rect 150910 115221 150922 115601
rect 151302 115221 151314 115601
rect 151694 115221 151706 115601
rect 152086 115221 152220 115601
rect 149220 115209 152220 115221
rect 149220 114829 149354 115209
rect 149734 114829 149746 115209
rect 150126 114829 150138 115209
rect 150518 114829 150530 115209
rect 150910 114829 150922 115209
rect 151302 114829 151314 115209
rect 151694 114829 151706 115209
rect 152086 114829 152220 115209
rect 149220 108750 152220 114829
rect 149220 108370 149354 108750
rect 149734 108370 149746 108750
rect 150126 108370 150138 108750
rect 150518 108370 150530 108750
rect 150910 108370 150922 108750
rect 151302 108370 151314 108750
rect 151694 108370 151706 108750
rect 152086 108370 152220 108750
rect 149220 101169 152220 108370
rect 149220 100789 149354 101169
rect 149734 100789 149746 101169
rect 150126 100789 150138 101169
rect 150518 100789 150530 101169
rect 150910 100789 150922 101169
rect 151302 100789 151314 101169
rect 151694 100789 151706 101169
rect 152086 100789 152220 101169
rect 149220 100777 152220 100789
rect 149220 100397 149354 100777
rect 149734 100397 149746 100777
rect 150126 100397 150138 100777
rect 150518 100397 150530 100777
rect 150910 100397 150922 100777
rect 151302 100397 151314 100777
rect 151694 100397 151706 100777
rect 152086 100397 152220 100777
rect 149220 100385 152220 100397
rect 149220 100005 149354 100385
rect 149734 100005 149746 100385
rect 150126 100005 150138 100385
rect 150518 100005 150530 100385
rect 150910 100005 150922 100385
rect 151302 100005 151314 100385
rect 151694 100005 151706 100385
rect 152086 100005 152220 100385
rect 149220 99993 152220 100005
rect 149220 99613 149354 99993
rect 149734 99613 149746 99993
rect 150126 99613 150138 99993
rect 150518 99613 150530 99993
rect 150910 99613 150922 99993
rect 151302 99613 151314 99993
rect 151694 99613 151706 99993
rect 152086 99613 152220 99993
rect 149220 99601 152220 99613
rect 149220 99221 149354 99601
rect 149734 99221 149746 99601
rect 150126 99221 150138 99601
rect 150518 99221 150530 99601
rect 150910 99221 150922 99601
rect 151302 99221 151314 99601
rect 151694 99221 151706 99601
rect 152086 99221 152220 99601
rect 149220 99209 152220 99221
rect 149220 98829 149354 99209
rect 149734 98829 149746 99209
rect 150126 98829 150138 99209
rect 150518 98829 150530 99209
rect 150910 98829 150922 99209
rect 151302 98829 151314 99209
rect 151694 98829 151706 99209
rect 152086 98829 152220 99209
rect 149220 93630 152220 98829
rect 149220 93250 149354 93630
rect 149734 93250 149746 93630
rect 150126 93250 150138 93630
rect 150518 93250 150530 93630
rect 150910 93250 150922 93630
rect 151302 93250 151314 93630
rect 151694 93250 151706 93630
rect 152086 93250 152220 93630
rect 149220 85169 152220 93250
rect 149220 84789 149354 85169
rect 149734 84789 149746 85169
rect 150126 84789 150138 85169
rect 150518 84789 150530 85169
rect 150910 84789 150922 85169
rect 151302 84789 151314 85169
rect 151694 84789 151706 85169
rect 152086 84789 152220 85169
rect 149220 84777 152220 84789
rect 149220 84397 149354 84777
rect 149734 84397 149746 84777
rect 150126 84397 150138 84777
rect 150518 84397 150530 84777
rect 150910 84397 150922 84777
rect 151302 84397 151314 84777
rect 151694 84397 151706 84777
rect 152086 84397 152220 84777
rect 149220 84385 152220 84397
rect 149220 84005 149354 84385
rect 149734 84005 149746 84385
rect 150126 84005 150138 84385
rect 150518 84005 150530 84385
rect 150910 84005 150922 84385
rect 151302 84005 151314 84385
rect 151694 84005 151706 84385
rect 152086 84005 152220 84385
rect 149220 83993 152220 84005
rect 149220 83613 149354 83993
rect 149734 83613 149746 83993
rect 150126 83613 150138 83993
rect 150518 83613 150530 83993
rect 150910 83613 150922 83993
rect 151302 83613 151314 83993
rect 151694 83613 151706 83993
rect 152086 83613 152220 83993
rect 149220 83601 152220 83613
rect 149220 83221 149354 83601
rect 149734 83221 149746 83601
rect 150126 83221 150138 83601
rect 150518 83221 150530 83601
rect 150910 83221 150922 83601
rect 151302 83221 151314 83601
rect 151694 83221 151706 83601
rect 152086 83221 152220 83601
rect 149220 83209 152220 83221
rect 149220 82829 149354 83209
rect 149734 82829 149746 83209
rect 150126 82829 150138 83209
rect 150518 82829 150530 83209
rect 150910 82829 150922 83209
rect 151302 82829 151314 83209
rect 151694 82829 151706 83209
rect 152086 82829 152220 83209
rect 149220 78510 152220 82829
rect 149220 78130 149354 78510
rect 149734 78130 149746 78510
rect 150126 78130 150138 78510
rect 150518 78130 150530 78510
rect 150910 78130 150922 78510
rect 151302 78130 151314 78510
rect 151694 78130 151706 78510
rect 152086 78130 152220 78510
rect 149220 74566 152220 78130
rect 149220 74186 149354 74566
rect 149734 74186 149746 74566
rect 150126 74186 150138 74566
rect 150518 74186 150530 74566
rect 150910 74186 150922 74566
rect 151302 74186 151314 74566
rect 151694 74186 151706 74566
rect 152086 74186 152220 74566
rect 149220 74174 152220 74186
rect 149220 73794 149354 74174
rect 149734 73794 149746 74174
rect 150126 73794 150138 74174
rect 150518 73794 150530 74174
rect 150910 73794 150922 74174
rect 151302 73794 151314 74174
rect 151694 73794 151706 74174
rect 152086 73794 152220 74174
rect 149220 73782 152220 73794
rect 149220 73402 149354 73782
rect 149734 73402 149746 73782
rect 150126 73402 150138 73782
rect 150518 73402 150530 73782
rect 150910 73402 150922 73782
rect 151302 73402 151314 73782
rect 151694 73402 151706 73782
rect 152086 73402 152220 73782
rect 149220 73390 152220 73402
rect 149220 73010 149354 73390
rect 149734 73010 149746 73390
rect 150126 73010 150138 73390
rect 150518 73010 150530 73390
rect 150910 73010 150922 73390
rect 151302 73010 151314 73390
rect 151694 73010 151706 73390
rect 152086 73010 152220 73390
rect 149220 72998 152220 73010
rect 149220 72618 149354 72998
rect 149734 72618 149746 72998
rect 150126 72618 150138 72998
rect 150518 72618 150530 72998
rect 150910 72618 150922 72998
rect 151302 72618 151314 72998
rect 151694 72618 151706 72998
rect 152086 72618 152220 72998
rect 149220 72606 152220 72618
rect 149220 72226 149354 72606
rect 149734 72226 149746 72606
rect 150126 72226 150138 72606
rect 150518 72226 150530 72606
rect 150910 72226 150922 72606
rect 151302 72226 151314 72606
rect 151694 72226 151706 72606
rect 152086 72226 152220 72606
rect 149220 72214 152220 72226
rect 149220 71834 149354 72214
rect 149734 71834 149746 72214
rect 150126 71834 150138 72214
rect 150518 71834 150530 72214
rect 150910 71834 150922 72214
rect 151302 71834 151314 72214
rect 151694 71834 151706 72214
rect 152086 71834 152220 72214
rect 149220 71700 152220 71834
rect 153220 140230 156220 153210
rect 153220 139850 153354 140230
rect 153734 139850 153746 140230
rect 154126 139850 154138 140230
rect 154518 139850 154530 140230
rect 154910 139850 154922 140230
rect 155302 139850 155314 140230
rect 155694 139850 155706 140230
rect 156086 139850 156220 140230
rect 153220 125110 156220 139850
rect 164400 133169 168000 133332
rect 164400 132789 164442 133169
rect 164822 132789 164834 133169
rect 165214 132789 165226 133169
rect 165606 132789 165618 133169
rect 165998 132789 166010 133169
rect 166390 132789 166402 133169
rect 166782 132789 166794 133169
rect 167174 132789 167186 133169
rect 167566 132789 167578 133169
rect 167958 132789 168000 133169
rect 164400 132777 168000 132789
rect 164400 132397 164442 132777
rect 164822 132397 164834 132777
rect 165214 132397 165226 132777
rect 165606 132397 165618 132777
rect 165998 132397 166010 132777
rect 166390 132397 166402 132777
rect 166782 132397 166794 132777
rect 167174 132397 167186 132777
rect 167566 132397 167578 132777
rect 167958 132397 168000 132777
rect 164400 132385 168000 132397
rect 164400 132005 164442 132385
rect 164822 132005 164834 132385
rect 165214 132005 165226 132385
rect 165606 132005 165618 132385
rect 165998 132005 166010 132385
rect 166390 132005 166402 132385
rect 166782 132005 166794 132385
rect 167174 132005 167186 132385
rect 167566 132005 167578 132385
rect 167958 132005 168000 132385
rect 164400 131993 168000 132005
rect 164400 131613 164442 131993
rect 164822 131613 164834 131993
rect 165214 131613 165226 131993
rect 165606 131613 165618 131993
rect 165998 131613 166010 131993
rect 166390 131613 166402 131993
rect 166782 131613 166794 131993
rect 167174 131613 167186 131993
rect 167566 131613 167578 131993
rect 167958 131613 168000 131993
rect 164400 131601 168000 131613
rect 164400 131221 164442 131601
rect 164822 131221 164834 131601
rect 165214 131221 165226 131601
rect 165606 131221 165618 131601
rect 165998 131221 166010 131601
rect 166390 131221 166402 131601
rect 166782 131221 166794 131601
rect 167174 131221 167186 131601
rect 167566 131221 167578 131601
rect 167958 131221 168000 131601
rect 164400 131209 168000 131221
rect 164400 130829 164442 131209
rect 164822 130829 164834 131209
rect 165214 130829 165226 131209
rect 165606 130829 165618 131209
rect 165998 130829 166010 131209
rect 166390 130829 166402 131209
rect 166782 130829 166794 131209
rect 167174 130829 167186 131209
rect 167566 130829 167578 131209
rect 167958 130829 168000 131209
rect 164400 130666 168000 130829
rect 153220 124730 153354 125110
rect 153734 124730 153746 125110
rect 154126 124730 154138 125110
rect 154518 124730 154530 125110
rect 154910 124730 154922 125110
rect 155302 124730 155314 125110
rect 155694 124730 155706 125110
rect 156086 124730 156220 125110
rect 153220 109990 156220 124730
rect 164400 117169 168000 117332
rect 164400 116789 164442 117169
rect 164822 116789 164834 117169
rect 165214 116789 165226 117169
rect 165606 116789 165618 117169
rect 165998 116789 166010 117169
rect 166390 116789 166402 117169
rect 166782 116789 166794 117169
rect 167174 116789 167186 117169
rect 167566 116789 167578 117169
rect 167958 116789 168000 117169
rect 164400 116777 168000 116789
rect 164400 116397 164442 116777
rect 164822 116397 164834 116777
rect 165214 116397 165226 116777
rect 165606 116397 165618 116777
rect 165998 116397 166010 116777
rect 166390 116397 166402 116777
rect 166782 116397 166794 116777
rect 167174 116397 167186 116777
rect 167566 116397 167578 116777
rect 167958 116397 168000 116777
rect 164400 116385 168000 116397
rect 164400 116005 164442 116385
rect 164822 116005 164834 116385
rect 165214 116005 165226 116385
rect 165606 116005 165618 116385
rect 165998 116005 166010 116385
rect 166390 116005 166402 116385
rect 166782 116005 166794 116385
rect 167174 116005 167186 116385
rect 167566 116005 167578 116385
rect 167958 116005 168000 116385
rect 164400 115993 168000 116005
rect 164400 115613 164442 115993
rect 164822 115613 164834 115993
rect 165214 115613 165226 115993
rect 165606 115613 165618 115993
rect 165998 115613 166010 115993
rect 166390 115613 166402 115993
rect 166782 115613 166794 115993
rect 167174 115613 167186 115993
rect 167566 115613 167578 115993
rect 167958 115613 168000 115993
rect 164400 115601 168000 115613
rect 164400 115221 164442 115601
rect 164822 115221 164834 115601
rect 165214 115221 165226 115601
rect 165606 115221 165618 115601
rect 165998 115221 166010 115601
rect 166390 115221 166402 115601
rect 166782 115221 166794 115601
rect 167174 115221 167186 115601
rect 167566 115221 167578 115601
rect 167958 115221 168000 115601
rect 164400 115209 168000 115221
rect 164400 114829 164442 115209
rect 164822 114829 164834 115209
rect 165214 114829 165226 115209
rect 165606 114829 165618 115209
rect 165998 114829 166010 115209
rect 166390 114829 166402 115209
rect 166782 114829 166794 115209
rect 167174 114829 167186 115209
rect 167566 114829 167578 115209
rect 167958 114829 168000 115209
rect 164400 114666 168000 114829
rect 153220 109610 153354 109990
rect 153734 109610 153746 109990
rect 154126 109610 154138 109990
rect 154518 109610 154530 109990
rect 154910 109610 154922 109990
rect 155302 109610 155314 109990
rect 155694 109610 155706 109990
rect 156086 109610 156220 109990
rect 153220 106501 156220 109610
rect 153220 106121 153354 106501
rect 153734 106121 153746 106501
rect 154126 106121 154138 106501
rect 154518 106121 154530 106501
rect 154910 106121 154922 106501
rect 155302 106121 155314 106501
rect 155694 106121 155706 106501
rect 156086 106121 156220 106501
rect 153220 106109 156220 106121
rect 153220 105729 153354 106109
rect 153734 105729 153746 106109
rect 154126 105729 154138 106109
rect 154518 105729 154530 106109
rect 154910 105729 154922 106109
rect 155302 105729 155314 106109
rect 155694 105729 155706 106109
rect 156086 105729 156220 106109
rect 153220 105717 156220 105729
rect 153220 105337 153354 105717
rect 153734 105337 153746 105717
rect 154126 105337 154138 105717
rect 154518 105337 154530 105717
rect 154910 105337 154922 105717
rect 155302 105337 155314 105717
rect 155694 105337 155706 105717
rect 156086 105337 156220 105717
rect 153220 105325 156220 105337
rect 153220 104945 153354 105325
rect 153734 104945 153746 105325
rect 154126 104945 154138 105325
rect 154518 104945 154530 105325
rect 154910 104945 154922 105325
rect 155302 104945 155314 105325
rect 155694 104945 155706 105325
rect 156086 104945 156220 105325
rect 153220 104933 156220 104945
rect 153220 104553 153354 104933
rect 153734 104553 153746 104933
rect 154126 104553 154138 104933
rect 154518 104553 154530 104933
rect 154910 104553 154922 104933
rect 155302 104553 155314 104933
rect 155694 104553 155706 104933
rect 156086 104553 156220 104933
rect 153220 104541 156220 104553
rect 153220 104161 153354 104541
rect 153734 104161 153746 104541
rect 154126 104161 154138 104541
rect 154518 104161 154530 104541
rect 154910 104161 154922 104541
rect 155302 104161 155314 104541
rect 155694 104161 155706 104541
rect 156086 104161 156220 104541
rect 153220 94870 156220 104161
rect 160400 106501 164000 106664
rect 160400 106121 160442 106501
rect 160822 106121 160834 106501
rect 161214 106121 161226 106501
rect 161606 106121 161618 106501
rect 161998 106121 162010 106501
rect 162390 106121 162402 106501
rect 162782 106121 162794 106501
rect 163174 106121 163186 106501
rect 163566 106121 163578 106501
rect 163958 106121 164000 106501
rect 160400 106109 164000 106121
rect 160400 105729 160442 106109
rect 160822 105729 160834 106109
rect 161214 105729 161226 106109
rect 161606 105729 161618 106109
rect 161998 105729 162010 106109
rect 162390 105729 162402 106109
rect 162782 105729 162794 106109
rect 163174 105729 163186 106109
rect 163566 105729 163578 106109
rect 163958 105729 164000 106109
rect 160400 105717 164000 105729
rect 160400 105337 160442 105717
rect 160822 105337 160834 105717
rect 161214 105337 161226 105717
rect 161606 105337 161618 105717
rect 161998 105337 162010 105717
rect 162390 105337 162402 105717
rect 162782 105337 162794 105717
rect 163174 105337 163186 105717
rect 163566 105337 163578 105717
rect 163958 105337 164000 105717
rect 160400 105325 164000 105337
rect 160400 104945 160442 105325
rect 160822 104945 160834 105325
rect 161214 104945 161226 105325
rect 161606 104945 161618 105325
rect 161998 104945 162010 105325
rect 162390 104945 162402 105325
rect 162782 104945 162794 105325
rect 163174 104945 163186 105325
rect 163566 104945 163578 105325
rect 163958 104945 164000 105325
rect 160400 104933 164000 104945
rect 160400 104553 160442 104933
rect 160822 104553 160834 104933
rect 161214 104553 161226 104933
rect 161606 104553 161618 104933
rect 161998 104553 162010 104933
rect 162390 104553 162402 104933
rect 162782 104553 162794 104933
rect 163174 104553 163186 104933
rect 163566 104553 163578 104933
rect 163958 104553 164000 104933
rect 160400 104541 164000 104553
rect 160400 104161 160442 104541
rect 160822 104161 160834 104541
rect 161214 104161 161226 104541
rect 161606 104161 161618 104541
rect 161998 104161 162010 104541
rect 162390 104161 162402 104541
rect 162782 104161 162794 104541
rect 163174 104161 163186 104541
rect 163566 104161 163578 104541
rect 163958 104161 164000 104541
rect 160400 103998 164000 104161
rect 164400 101169 168000 101332
rect 164400 100789 164442 101169
rect 164822 100789 164834 101169
rect 165214 100789 165226 101169
rect 165606 100789 165618 101169
rect 165998 100789 166010 101169
rect 166390 100789 166402 101169
rect 166782 100789 166794 101169
rect 167174 100789 167186 101169
rect 167566 100789 167578 101169
rect 167958 100789 168000 101169
rect 164400 100777 168000 100789
rect 164400 100397 164442 100777
rect 164822 100397 164834 100777
rect 165214 100397 165226 100777
rect 165606 100397 165618 100777
rect 165998 100397 166010 100777
rect 166390 100397 166402 100777
rect 166782 100397 166794 100777
rect 167174 100397 167186 100777
rect 167566 100397 167578 100777
rect 167958 100397 168000 100777
rect 164400 100385 168000 100397
rect 164400 100005 164442 100385
rect 164822 100005 164834 100385
rect 165214 100005 165226 100385
rect 165606 100005 165618 100385
rect 165998 100005 166010 100385
rect 166390 100005 166402 100385
rect 166782 100005 166794 100385
rect 167174 100005 167186 100385
rect 167566 100005 167578 100385
rect 167958 100005 168000 100385
rect 164400 99993 168000 100005
rect 164400 99613 164442 99993
rect 164822 99613 164834 99993
rect 165214 99613 165226 99993
rect 165606 99613 165618 99993
rect 165998 99613 166010 99993
rect 166390 99613 166402 99993
rect 166782 99613 166794 99993
rect 167174 99613 167186 99993
rect 167566 99613 167578 99993
rect 167958 99613 168000 99993
rect 164400 99601 168000 99613
rect 164400 99221 164442 99601
rect 164822 99221 164834 99601
rect 165214 99221 165226 99601
rect 165606 99221 165618 99601
rect 165998 99221 166010 99601
rect 166390 99221 166402 99601
rect 166782 99221 166794 99601
rect 167174 99221 167186 99601
rect 167566 99221 167578 99601
rect 167958 99221 168000 99601
rect 164400 99209 168000 99221
rect 164400 98829 164442 99209
rect 164822 98829 164834 99209
rect 165214 98829 165226 99209
rect 165606 98829 165618 99209
rect 165998 98829 166010 99209
rect 166390 98829 166402 99209
rect 166782 98829 166794 99209
rect 167174 98829 167186 99209
rect 167566 98829 167578 99209
rect 167958 98829 168000 99209
rect 164400 98666 168000 98829
rect 153220 94490 153354 94870
rect 153734 94490 153746 94870
rect 154126 94490 154138 94870
rect 154518 94490 154530 94870
rect 154910 94490 154922 94870
rect 155302 94490 155314 94870
rect 155694 94490 155706 94870
rect 156086 94490 156220 94870
rect 153220 90501 156220 94490
rect 153220 90121 153354 90501
rect 153734 90121 153746 90501
rect 154126 90121 154138 90501
rect 154518 90121 154530 90501
rect 154910 90121 154922 90501
rect 155302 90121 155314 90501
rect 155694 90121 155706 90501
rect 156086 90121 156220 90501
rect 153220 90109 156220 90121
rect 153220 89729 153354 90109
rect 153734 89729 153746 90109
rect 154126 89729 154138 90109
rect 154518 89729 154530 90109
rect 154910 89729 154922 90109
rect 155302 89729 155314 90109
rect 155694 89729 155706 90109
rect 156086 89729 156220 90109
rect 153220 89717 156220 89729
rect 153220 89337 153354 89717
rect 153734 89337 153746 89717
rect 154126 89337 154138 89717
rect 154518 89337 154530 89717
rect 154910 89337 154922 89717
rect 155302 89337 155314 89717
rect 155694 89337 155706 89717
rect 156086 89337 156220 89717
rect 153220 89325 156220 89337
rect 153220 88945 153354 89325
rect 153734 88945 153746 89325
rect 154126 88945 154138 89325
rect 154518 88945 154530 89325
rect 154910 88945 154922 89325
rect 155302 88945 155314 89325
rect 155694 88945 155706 89325
rect 156086 88945 156220 89325
rect 153220 88933 156220 88945
rect 153220 88553 153354 88933
rect 153734 88553 153746 88933
rect 154126 88553 154138 88933
rect 154518 88553 154530 88933
rect 154910 88553 154922 88933
rect 155302 88553 155314 88933
rect 155694 88553 155706 88933
rect 156086 88553 156220 88933
rect 153220 88541 156220 88553
rect 153220 88161 153354 88541
rect 153734 88161 153746 88541
rect 154126 88161 154138 88541
rect 154518 88161 154530 88541
rect 154910 88161 154922 88541
rect 155302 88161 155314 88541
rect 155694 88161 155706 88541
rect 156086 88161 156220 88541
rect 153220 79750 156220 88161
rect 160400 90501 164000 90664
rect 160400 90121 160442 90501
rect 160822 90121 160834 90501
rect 161214 90121 161226 90501
rect 161606 90121 161618 90501
rect 161998 90121 162010 90501
rect 162390 90121 162402 90501
rect 162782 90121 162794 90501
rect 163174 90121 163186 90501
rect 163566 90121 163578 90501
rect 163958 90121 164000 90501
rect 160400 90109 164000 90121
rect 160400 89729 160442 90109
rect 160822 89729 160834 90109
rect 161214 89729 161226 90109
rect 161606 89729 161618 90109
rect 161998 89729 162010 90109
rect 162390 89729 162402 90109
rect 162782 89729 162794 90109
rect 163174 89729 163186 90109
rect 163566 89729 163578 90109
rect 163958 89729 164000 90109
rect 160400 89717 164000 89729
rect 160400 89337 160442 89717
rect 160822 89337 160834 89717
rect 161214 89337 161226 89717
rect 161606 89337 161618 89717
rect 161998 89337 162010 89717
rect 162390 89337 162402 89717
rect 162782 89337 162794 89717
rect 163174 89337 163186 89717
rect 163566 89337 163578 89717
rect 163958 89337 164000 89717
rect 160400 89325 164000 89337
rect 160400 88945 160442 89325
rect 160822 88945 160834 89325
rect 161214 88945 161226 89325
rect 161606 88945 161618 89325
rect 161998 88945 162010 89325
rect 162390 88945 162402 89325
rect 162782 88945 162794 89325
rect 163174 88945 163186 89325
rect 163566 88945 163578 89325
rect 163958 88945 164000 89325
rect 160400 88933 164000 88945
rect 160400 88553 160442 88933
rect 160822 88553 160834 88933
rect 161214 88553 161226 88933
rect 161606 88553 161618 88933
rect 161998 88553 162010 88933
rect 162390 88553 162402 88933
rect 162782 88553 162794 88933
rect 163174 88553 163186 88933
rect 163566 88553 163578 88933
rect 163958 88553 164000 88933
rect 160400 88541 164000 88553
rect 160400 88161 160442 88541
rect 160822 88161 160834 88541
rect 161214 88161 161226 88541
rect 161606 88161 161618 88541
rect 161998 88161 162010 88541
rect 162390 88161 162402 88541
rect 162782 88161 162794 88541
rect 163174 88161 163186 88541
rect 163566 88161 163578 88541
rect 163958 88161 164000 88541
rect 160400 87998 164000 88161
rect 164400 85169 168000 85332
rect 164400 84789 164442 85169
rect 164822 84789 164834 85169
rect 165214 84789 165226 85169
rect 165606 84789 165618 85169
rect 165998 84789 166010 85169
rect 166390 84789 166402 85169
rect 166782 84789 166794 85169
rect 167174 84789 167186 85169
rect 167566 84789 167578 85169
rect 167958 84789 168000 85169
rect 164400 84777 168000 84789
rect 164400 84397 164442 84777
rect 164822 84397 164834 84777
rect 165214 84397 165226 84777
rect 165606 84397 165618 84777
rect 165998 84397 166010 84777
rect 166390 84397 166402 84777
rect 166782 84397 166794 84777
rect 167174 84397 167186 84777
rect 167566 84397 167578 84777
rect 167958 84397 168000 84777
rect 164400 84385 168000 84397
rect 164400 84005 164442 84385
rect 164822 84005 164834 84385
rect 165214 84005 165226 84385
rect 165606 84005 165618 84385
rect 165998 84005 166010 84385
rect 166390 84005 166402 84385
rect 166782 84005 166794 84385
rect 167174 84005 167186 84385
rect 167566 84005 167578 84385
rect 167958 84005 168000 84385
rect 164400 83993 168000 84005
rect 164400 83613 164442 83993
rect 164822 83613 164834 83993
rect 165214 83613 165226 83993
rect 165606 83613 165618 83993
rect 165998 83613 166010 83993
rect 166390 83613 166402 83993
rect 166782 83613 166794 83993
rect 167174 83613 167186 83993
rect 167566 83613 167578 83993
rect 167958 83613 168000 83993
rect 164400 83601 168000 83613
rect 164400 83221 164442 83601
rect 164822 83221 164834 83601
rect 165214 83221 165226 83601
rect 165606 83221 165618 83601
rect 165998 83221 166010 83601
rect 166390 83221 166402 83601
rect 166782 83221 166794 83601
rect 167174 83221 167186 83601
rect 167566 83221 167578 83601
rect 167958 83221 168000 83601
rect 164400 83209 168000 83221
rect 164400 82829 164442 83209
rect 164822 82829 164834 83209
rect 165214 82829 165226 83209
rect 165606 82829 165618 83209
rect 165998 82829 166010 83209
rect 166390 82829 166402 83209
rect 166782 82829 166794 83209
rect 167174 82829 167186 83209
rect 167566 82829 167578 83209
rect 167958 82829 168000 83209
rect 164400 82666 168000 82829
rect 153220 79370 153354 79750
rect 153734 79370 153746 79750
rect 154126 79370 154138 79750
rect 154518 79370 154530 79750
rect 154910 79370 154922 79750
rect 155302 79370 155314 79750
rect 155694 79370 155706 79750
rect 156086 79370 156220 79750
rect 153220 74501 156220 79370
rect 153220 74121 153354 74501
rect 153734 74121 153746 74501
rect 154126 74121 154138 74501
rect 154518 74121 154530 74501
rect 154910 74121 154922 74501
rect 155302 74121 155314 74501
rect 155694 74121 155706 74501
rect 156086 74121 156220 74501
rect 153220 74109 156220 74121
rect 153220 73729 153354 74109
rect 153734 73729 153746 74109
rect 154126 73729 154138 74109
rect 154518 73729 154530 74109
rect 154910 73729 154922 74109
rect 155302 73729 155314 74109
rect 155694 73729 155706 74109
rect 156086 73729 156220 74109
rect 153220 73717 156220 73729
rect 153220 73337 153354 73717
rect 153734 73337 153746 73717
rect 154126 73337 154138 73717
rect 154518 73337 154530 73717
rect 154910 73337 154922 73717
rect 155302 73337 155314 73717
rect 155694 73337 155706 73717
rect 156086 73337 156220 73717
rect 153220 73325 156220 73337
rect 153220 72945 153354 73325
rect 153734 72945 153746 73325
rect 154126 72945 154138 73325
rect 154518 72945 154530 73325
rect 154910 72945 154922 73325
rect 155302 72945 155314 73325
rect 155694 72945 155706 73325
rect 156086 72945 156220 73325
rect 153220 72933 156220 72945
rect 153220 72553 153354 72933
rect 153734 72553 153746 72933
rect 154126 72553 154138 72933
rect 154518 72553 154530 72933
rect 154910 72553 154922 72933
rect 155302 72553 155314 72933
rect 155694 72553 155706 72933
rect 156086 72553 156220 72933
rect 153220 72541 156220 72553
rect 153220 72161 153354 72541
rect 153734 72161 153746 72541
rect 154126 72161 154138 72541
rect 154518 72161 154530 72541
rect 154910 72161 154922 72541
rect 155302 72161 155314 72541
rect 155694 72161 155706 72541
rect 156086 72161 156220 72541
rect 139868 70186 139898 70566
rect 140278 70186 140308 70566
rect 139868 70174 140308 70186
rect 139868 69794 139898 70174
rect 140278 69794 140308 70174
rect 139868 69782 140308 69794
rect 139868 69402 139898 69782
rect 140278 69402 140308 69782
rect 139868 69390 140308 69402
rect 139868 69010 139898 69390
rect 140278 69010 140308 69390
rect 139868 68998 140308 69010
rect 139868 68618 139898 68998
rect 140278 68618 140308 68998
rect 139868 68606 140308 68618
rect 139868 68226 139898 68606
rect 140278 68226 140308 68606
rect 139868 68214 140308 68226
rect 139868 67834 139898 68214
rect 140278 67834 140308 68214
rect 139868 67700 140308 67834
rect 153220 70566 156220 72161
rect 160400 74501 164000 74664
rect 160400 74121 160442 74501
rect 160822 74121 160834 74501
rect 161214 74121 161226 74501
rect 161606 74121 161618 74501
rect 161998 74121 162010 74501
rect 162390 74121 162402 74501
rect 162782 74121 162794 74501
rect 163174 74121 163186 74501
rect 163566 74121 163578 74501
rect 163958 74121 164000 74501
rect 160400 74109 164000 74121
rect 160400 73729 160442 74109
rect 160822 73729 160834 74109
rect 161214 73729 161226 74109
rect 161606 73729 161618 74109
rect 161998 73729 162010 74109
rect 162390 73729 162402 74109
rect 162782 73729 162794 74109
rect 163174 73729 163186 74109
rect 163566 73729 163578 74109
rect 163958 73729 164000 74109
rect 160400 73717 164000 73729
rect 160400 73337 160442 73717
rect 160822 73337 160834 73717
rect 161214 73337 161226 73717
rect 161606 73337 161618 73717
rect 161998 73337 162010 73717
rect 162390 73337 162402 73717
rect 162782 73337 162794 73717
rect 163174 73337 163186 73717
rect 163566 73337 163578 73717
rect 163958 73337 164000 73717
rect 160400 73325 164000 73337
rect 160400 72945 160442 73325
rect 160822 72945 160834 73325
rect 161214 72945 161226 73325
rect 161606 72945 161618 73325
rect 161998 72945 162010 73325
rect 162390 72945 162402 73325
rect 162782 72945 162794 73325
rect 163174 72945 163186 73325
rect 163566 72945 163578 73325
rect 163958 72945 164000 73325
rect 160400 72933 164000 72945
rect 160400 72553 160442 72933
rect 160822 72553 160834 72933
rect 161214 72553 161226 72933
rect 161606 72553 161618 72933
rect 161998 72553 162010 72933
rect 162390 72553 162402 72933
rect 162782 72553 162794 72933
rect 163174 72553 163186 72933
rect 163566 72553 163578 72933
rect 163958 72553 164000 72933
rect 160400 72541 164000 72553
rect 160400 72161 160442 72541
rect 160822 72161 160834 72541
rect 161214 72161 161226 72541
rect 161606 72161 161618 72541
rect 161998 72161 162010 72541
rect 162390 72161 162402 72541
rect 162782 72161 162794 72541
rect 163174 72161 163186 72541
rect 163566 72161 163578 72541
rect 163958 72161 164000 72541
rect 160400 71998 164000 72161
rect 153220 70186 153354 70566
rect 153734 70186 153746 70566
rect 154126 70186 154138 70566
rect 154518 70186 154530 70566
rect 154910 70186 154922 70566
rect 155302 70186 155314 70566
rect 155694 70186 155706 70566
rect 156086 70186 156220 70566
rect 153220 70174 156220 70186
rect 153220 69794 153354 70174
rect 153734 69794 153746 70174
rect 154126 69794 154138 70174
rect 154518 69794 154530 70174
rect 154910 69794 154922 70174
rect 155302 69794 155314 70174
rect 155694 69794 155706 70174
rect 156086 69794 156220 70174
rect 153220 69782 156220 69794
rect 153220 69402 153354 69782
rect 153734 69402 153746 69782
rect 154126 69402 154138 69782
rect 154518 69402 154530 69782
rect 154910 69402 154922 69782
rect 155302 69402 155314 69782
rect 155694 69402 155706 69782
rect 156086 69402 156220 69782
rect 153220 69390 156220 69402
rect 153220 69010 153354 69390
rect 153734 69010 153746 69390
rect 154126 69010 154138 69390
rect 154518 69010 154530 69390
rect 154910 69010 154922 69390
rect 155302 69010 155314 69390
rect 155694 69010 155706 69390
rect 156086 69010 156220 69390
rect 153220 68998 156220 69010
rect 153220 68618 153354 68998
rect 153734 68618 153746 68998
rect 154126 68618 154138 68998
rect 154518 68618 154530 68998
rect 154910 68618 154922 68998
rect 155302 68618 155314 68998
rect 155694 68618 155706 68998
rect 156086 68618 156220 68998
rect 153220 68606 156220 68618
rect 153220 68226 153354 68606
rect 153734 68226 153746 68606
rect 154126 68226 154138 68606
rect 154518 68226 154530 68606
rect 154910 68226 154922 68606
rect 155302 68226 155314 68606
rect 155694 68226 155706 68606
rect 156086 68226 156220 68606
rect 153220 68214 156220 68226
rect 153220 67834 153354 68214
rect 153734 67834 153746 68214
rect 154126 67834 154138 68214
rect 154518 67834 154530 68214
rect 154910 67834 154922 68214
rect 155302 67834 155314 68214
rect 155694 67834 155706 68214
rect 156086 67834 156220 68214
rect 153220 67700 156220 67834
<< via6 >>
rect 67882 155562 68262 155942
rect 68274 155562 68654 155942
rect 68666 155562 69046 155942
rect 69058 155562 69438 155942
rect 69450 155562 69830 155942
rect 69842 155562 70222 155942
rect 70234 155562 70614 155942
rect 67882 155170 68262 155550
rect 68274 155170 68654 155550
rect 68666 155170 69046 155550
rect 69058 155170 69438 155550
rect 69450 155170 69830 155550
rect 69842 155170 70222 155550
rect 70234 155170 70614 155550
rect 67882 154778 68262 155158
rect 68274 154778 68654 155158
rect 68666 154778 69046 155158
rect 69058 154778 69438 155158
rect 69450 154778 69830 155158
rect 69842 154778 70222 155158
rect 70234 154778 70614 155158
rect 67882 154386 68262 154766
rect 68274 154386 68654 154766
rect 68666 154386 69046 154766
rect 69058 154386 69438 154766
rect 69450 154386 69830 154766
rect 69842 154386 70222 154766
rect 70234 154386 70614 154766
rect 67882 153994 68262 154374
rect 68274 153994 68654 154374
rect 68666 153994 69046 154374
rect 69058 153994 69438 154374
rect 69450 153994 69830 154374
rect 69842 153994 70222 154374
rect 70234 153994 70614 154374
rect 67882 153602 68262 153982
rect 68274 153602 68654 153982
rect 68666 153602 69046 153982
rect 69058 153602 69438 153982
rect 69450 153602 69830 153982
rect 69842 153602 70222 153982
rect 70234 153602 70614 153982
rect 67882 153210 68262 153590
rect 68274 153210 68654 153590
rect 68666 153210 69046 153590
rect 69058 153210 69438 153590
rect 69450 153210 69830 153590
rect 69842 153210 70222 153590
rect 70234 153210 70614 153590
rect 79418 155562 79798 155942
rect 79418 155170 79798 155550
rect 79418 154778 79798 155158
rect 79418 154386 79798 154766
rect 79418 153994 79798 154374
rect 79418 153602 79798 153982
rect 79418 153210 79798 153590
rect 67882 139850 68262 140230
rect 68274 139850 68654 140230
rect 68666 139850 69046 140230
rect 69058 139850 69438 140230
rect 69450 139850 69830 140230
rect 69842 139850 70222 140230
rect 70234 139850 70614 140230
rect 56042 132789 56422 133169
rect 56434 132789 56814 133169
rect 56826 132789 57206 133169
rect 57218 132789 57598 133169
rect 57610 132789 57990 133169
rect 58002 132789 58382 133169
rect 58394 132789 58774 133169
rect 58786 132789 59166 133169
rect 59178 132789 59558 133169
rect 56042 132397 56422 132777
rect 56434 132397 56814 132777
rect 56826 132397 57206 132777
rect 57218 132397 57598 132777
rect 57610 132397 57990 132777
rect 58002 132397 58382 132777
rect 58394 132397 58774 132777
rect 58786 132397 59166 132777
rect 59178 132397 59558 132777
rect 56042 132005 56422 132385
rect 56434 132005 56814 132385
rect 56826 132005 57206 132385
rect 57218 132005 57598 132385
rect 57610 132005 57990 132385
rect 58002 132005 58382 132385
rect 58394 132005 58774 132385
rect 58786 132005 59166 132385
rect 59178 132005 59558 132385
rect 56042 131613 56422 131993
rect 56434 131613 56814 131993
rect 56826 131613 57206 131993
rect 57218 131613 57598 131993
rect 57610 131613 57990 131993
rect 58002 131613 58382 131993
rect 58394 131613 58774 131993
rect 58786 131613 59166 131993
rect 59178 131613 59558 131993
rect 56042 131221 56422 131601
rect 56434 131221 56814 131601
rect 56826 131221 57206 131601
rect 57218 131221 57598 131601
rect 57610 131221 57990 131601
rect 58002 131221 58382 131601
rect 58394 131221 58774 131601
rect 58786 131221 59166 131601
rect 59178 131221 59558 131601
rect 56042 130829 56422 131209
rect 56434 130829 56814 131209
rect 56826 130829 57206 131209
rect 57218 130829 57598 131209
rect 57610 130829 57990 131209
rect 58002 130829 58382 131209
rect 58394 130829 58774 131209
rect 58786 130829 59166 131209
rect 59178 130829 59558 131209
rect 67882 124730 68262 125110
rect 68274 124730 68654 125110
rect 68666 124730 69046 125110
rect 69058 124730 69438 125110
rect 69450 124730 69830 125110
rect 69842 124730 70222 125110
rect 70234 124730 70614 125110
rect 56042 116789 56422 117169
rect 56434 116789 56814 117169
rect 56826 116789 57206 117169
rect 57218 116789 57598 117169
rect 57610 116789 57990 117169
rect 58002 116789 58382 117169
rect 58394 116789 58774 117169
rect 58786 116789 59166 117169
rect 59178 116789 59558 117169
rect 56042 116397 56422 116777
rect 56434 116397 56814 116777
rect 56826 116397 57206 116777
rect 57218 116397 57598 116777
rect 57610 116397 57990 116777
rect 58002 116397 58382 116777
rect 58394 116397 58774 116777
rect 58786 116397 59166 116777
rect 59178 116397 59558 116777
rect 56042 116005 56422 116385
rect 56434 116005 56814 116385
rect 56826 116005 57206 116385
rect 57218 116005 57598 116385
rect 57610 116005 57990 116385
rect 58002 116005 58382 116385
rect 58394 116005 58774 116385
rect 58786 116005 59166 116385
rect 59178 116005 59558 116385
rect 56042 115613 56422 115993
rect 56434 115613 56814 115993
rect 56826 115613 57206 115993
rect 57218 115613 57598 115993
rect 57610 115613 57990 115993
rect 58002 115613 58382 115993
rect 58394 115613 58774 115993
rect 58786 115613 59166 115993
rect 59178 115613 59558 115993
rect 56042 115221 56422 115601
rect 56434 115221 56814 115601
rect 56826 115221 57206 115601
rect 57218 115221 57598 115601
rect 57610 115221 57990 115601
rect 58002 115221 58382 115601
rect 58394 115221 58774 115601
rect 58786 115221 59166 115601
rect 59178 115221 59558 115601
rect 56042 114829 56422 115209
rect 56434 114829 56814 115209
rect 56826 114829 57206 115209
rect 57218 114829 57598 115209
rect 57610 114829 57990 115209
rect 58002 114829 58382 115209
rect 58394 114829 58774 115209
rect 58786 114829 59166 115209
rect 59178 114829 59558 115209
rect 67882 109610 68262 109990
rect 68274 109610 68654 109990
rect 68666 109610 69046 109990
rect 69058 109610 69438 109990
rect 69450 109610 69830 109990
rect 69842 109610 70222 109990
rect 70234 109610 70614 109990
rect 60042 106121 60422 106501
rect 60434 106121 60814 106501
rect 60826 106121 61206 106501
rect 61218 106121 61598 106501
rect 61610 106121 61990 106501
rect 62002 106121 62382 106501
rect 62394 106121 62774 106501
rect 62786 106121 63166 106501
rect 63178 106121 63558 106501
rect 60042 105729 60422 106109
rect 60434 105729 60814 106109
rect 60826 105729 61206 106109
rect 61218 105729 61598 106109
rect 61610 105729 61990 106109
rect 62002 105729 62382 106109
rect 62394 105729 62774 106109
rect 62786 105729 63166 106109
rect 63178 105729 63558 106109
rect 60042 105337 60422 105717
rect 60434 105337 60814 105717
rect 60826 105337 61206 105717
rect 61218 105337 61598 105717
rect 61610 105337 61990 105717
rect 62002 105337 62382 105717
rect 62394 105337 62774 105717
rect 62786 105337 63166 105717
rect 63178 105337 63558 105717
rect 60042 104945 60422 105325
rect 60434 104945 60814 105325
rect 60826 104945 61206 105325
rect 61218 104945 61598 105325
rect 61610 104945 61990 105325
rect 62002 104945 62382 105325
rect 62394 104945 62774 105325
rect 62786 104945 63166 105325
rect 63178 104945 63558 105325
rect 60042 104553 60422 104933
rect 60434 104553 60814 104933
rect 60826 104553 61206 104933
rect 61218 104553 61598 104933
rect 61610 104553 61990 104933
rect 62002 104553 62382 104933
rect 62394 104553 62774 104933
rect 62786 104553 63166 104933
rect 63178 104553 63558 104933
rect 60042 104161 60422 104541
rect 60434 104161 60814 104541
rect 60826 104161 61206 104541
rect 61218 104161 61598 104541
rect 61610 104161 61990 104541
rect 62002 104161 62382 104541
rect 62394 104161 62774 104541
rect 62786 104161 63166 104541
rect 63178 104161 63558 104541
rect 67882 106121 68262 106501
rect 68274 106121 68654 106501
rect 68666 106121 69046 106501
rect 69058 106121 69438 106501
rect 69450 106121 69830 106501
rect 69842 106121 70222 106501
rect 70234 106121 70614 106501
rect 67882 105729 68262 106109
rect 68274 105729 68654 106109
rect 68666 105729 69046 106109
rect 69058 105729 69438 106109
rect 69450 105729 69830 106109
rect 69842 105729 70222 106109
rect 70234 105729 70614 106109
rect 67882 105337 68262 105717
rect 68274 105337 68654 105717
rect 68666 105337 69046 105717
rect 69058 105337 69438 105717
rect 69450 105337 69830 105717
rect 69842 105337 70222 105717
rect 70234 105337 70614 105717
rect 67882 104945 68262 105325
rect 68274 104945 68654 105325
rect 68666 104945 69046 105325
rect 69058 104945 69438 105325
rect 69450 104945 69830 105325
rect 69842 104945 70222 105325
rect 70234 104945 70614 105325
rect 67882 104553 68262 104933
rect 68274 104553 68654 104933
rect 68666 104553 69046 104933
rect 69058 104553 69438 104933
rect 69450 104553 69830 104933
rect 69842 104553 70222 104933
rect 70234 104553 70614 104933
rect 67882 104161 68262 104541
rect 68274 104161 68654 104541
rect 68666 104161 69046 104541
rect 69058 104161 69438 104541
rect 69450 104161 69830 104541
rect 69842 104161 70222 104541
rect 70234 104161 70614 104541
rect 56042 100789 56422 101169
rect 56434 100789 56814 101169
rect 56826 100789 57206 101169
rect 57218 100789 57598 101169
rect 57610 100789 57990 101169
rect 58002 100789 58382 101169
rect 58394 100789 58774 101169
rect 58786 100789 59166 101169
rect 59178 100789 59558 101169
rect 56042 100397 56422 100777
rect 56434 100397 56814 100777
rect 56826 100397 57206 100777
rect 57218 100397 57598 100777
rect 57610 100397 57990 100777
rect 58002 100397 58382 100777
rect 58394 100397 58774 100777
rect 58786 100397 59166 100777
rect 59178 100397 59558 100777
rect 56042 100005 56422 100385
rect 56434 100005 56814 100385
rect 56826 100005 57206 100385
rect 57218 100005 57598 100385
rect 57610 100005 57990 100385
rect 58002 100005 58382 100385
rect 58394 100005 58774 100385
rect 58786 100005 59166 100385
rect 59178 100005 59558 100385
rect 56042 99613 56422 99993
rect 56434 99613 56814 99993
rect 56826 99613 57206 99993
rect 57218 99613 57598 99993
rect 57610 99613 57990 99993
rect 58002 99613 58382 99993
rect 58394 99613 58774 99993
rect 58786 99613 59166 99993
rect 59178 99613 59558 99993
rect 56042 99221 56422 99601
rect 56434 99221 56814 99601
rect 56826 99221 57206 99601
rect 57218 99221 57598 99601
rect 57610 99221 57990 99601
rect 58002 99221 58382 99601
rect 58394 99221 58774 99601
rect 58786 99221 59166 99601
rect 59178 99221 59558 99601
rect 56042 98829 56422 99209
rect 56434 98829 56814 99209
rect 56826 98829 57206 99209
rect 57218 98829 57598 99209
rect 57610 98829 57990 99209
rect 58002 98829 58382 99209
rect 58394 98829 58774 99209
rect 58786 98829 59166 99209
rect 59178 98829 59558 99209
rect 67882 94490 68262 94870
rect 68274 94490 68654 94870
rect 68666 94490 69046 94870
rect 69058 94490 69438 94870
rect 69450 94490 69830 94870
rect 69842 94490 70222 94870
rect 70234 94490 70614 94870
rect 60042 90121 60422 90501
rect 60434 90121 60814 90501
rect 60826 90121 61206 90501
rect 61218 90121 61598 90501
rect 61610 90121 61990 90501
rect 62002 90121 62382 90501
rect 62394 90121 62774 90501
rect 62786 90121 63166 90501
rect 63178 90121 63558 90501
rect 60042 89729 60422 90109
rect 60434 89729 60814 90109
rect 60826 89729 61206 90109
rect 61218 89729 61598 90109
rect 61610 89729 61990 90109
rect 62002 89729 62382 90109
rect 62394 89729 62774 90109
rect 62786 89729 63166 90109
rect 63178 89729 63558 90109
rect 60042 89337 60422 89717
rect 60434 89337 60814 89717
rect 60826 89337 61206 89717
rect 61218 89337 61598 89717
rect 61610 89337 61990 89717
rect 62002 89337 62382 89717
rect 62394 89337 62774 89717
rect 62786 89337 63166 89717
rect 63178 89337 63558 89717
rect 60042 88945 60422 89325
rect 60434 88945 60814 89325
rect 60826 88945 61206 89325
rect 61218 88945 61598 89325
rect 61610 88945 61990 89325
rect 62002 88945 62382 89325
rect 62394 88945 62774 89325
rect 62786 88945 63166 89325
rect 63178 88945 63558 89325
rect 60042 88553 60422 88933
rect 60434 88553 60814 88933
rect 60826 88553 61206 88933
rect 61218 88553 61598 88933
rect 61610 88553 61990 88933
rect 62002 88553 62382 88933
rect 62394 88553 62774 88933
rect 62786 88553 63166 88933
rect 63178 88553 63558 88933
rect 60042 88161 60422 88541
rect 60434 88161 60814 88541
rect 60826 88161 61206 88541
rect 61218 88161 61598 88541
rect 61610 88161 61990 88541
rect 62002 88161 62382 88541
rect 62394 88161 62774 88541
rect 62786 88161 63166 88541
rect 63178 88161 63558 88541
rect 67882 90121 68262 90501
rect 68274 90121 68654 90501
rect 68666 90121 69046 90501
rect 69058 90121 69438 90501
rect 69450 90121 69830 90501
rect 69842 90121 70222 90501
rect 70234 90121 70614 90501
rect 67882 89729 68262 90109
rect 68274 89729 68654 90109
rect 68666 89729 69046 90109
rect 69058 89729 69438 90109
rect 69450 89729 69830 90109
rect 69842 89729 70222 90109
rect 70234 89729 70614 90109
rect 67882 89337 68262 89717
rect 68274 89337 68654 89717
rect 68666 89337 69046 89717
rect 69058 89337 69438 89717
rect 69450 89337 69830 89717
rect 69842 89337 70222 89717
rect 70234 89337 70614 89717
rect 67882 88945 68262 89325
rect 68274 88945 68654 89325
rect 68666 88945 69046 89325
rect 69058 88945 69438 89325
rect 69450 88945 69830 89325
rect 69842 88945 70222 89325
rect 70234 88945 70614 89325
rect 67882 88553 68262 88933
rect 68274 88553 68654 88933
rect 68666 88553 69046 88933
rect 69058 88553 69438 88933
rect 69450 88553 69830 88933
rect 69842 88553 70222 88933
rect 70234 88553 70614 88933
rect 67882 88161 68262 88541
rect 68274 88161 68654 88541
rect 68666 88161 69046 88541
rect 69058 88161 69438 88541
rect 69450 88161 69830 88541
rect 69842 88161 70222 88541
rect 70234 88161 70614 88541
rect 56042 84789 56422 85169
rect 56434 84789 56814 85169
rect 56826 84789 57206 85169
rect 57218 84789 57598 85169
rect 57610 84789 57990 85169
rect 58002 84789 58382 85169
rect 58394 84789 58774 85169
rect 58786 84789 59166 85169
rect 59178 84789 59558 85169
rect 56042 84397 56422 84777
rect 56434 84397 56814 84777
rect 56826 84397 57206 84777
rect 57218 84397 57598 84777
rect 57610 84397 57990 84777
rect 58002 84397 58382 84777
rect 58394 84397 58774 84777
rect 58786 84397 59166 84777
rect 59178 84397 59558 84777
rect 56042 84005 56422 84385
rect 56434 84005 56814 84385
rect 56826 84005 57206 84385
rect 57218 84005 57598 84385
rect 57610 84005 57990 84385
rect 58002 84005 58382 84385
rect 58394 84005 58774 84385
rect 58786 84005 59166 84385
rect 59178 84005 59558 84385
rect 56042 83613 56422 83993
rect 56434 83613 56814 83993
rect 56826 83613 57206 83993
rect 57218 83613 57598 83993
rect 57610 83613 57990 83993
rect 58002 83613 58382 83993
rect 58394 83613 58774 83993
rect 58786 83613 59166 83993
rect 59178 83613 59558 83993
rect 56042 83221 56422 83601
rect 56434 83221 56814 83601
rect 56826 83221 57206 83601
rect 57218 83221 57598 83601
rect 57610 83221 57990 83601
rect 58002 83221 58382 83601
rect 58394 83221 58774 83601
rect 58786 83221 59166 83601
rect 59178 83221 59558 83601
rect 56042 82829 56422 83209
rect 56434 82829 56814 83209
rect 56826 82829 57206 83209
rect 57218 82829 57598 83209
rect 57610 82829 57990 83209
rect 58002 82829 58382 83209
rect 58394 82829 58774 83209
rect 58786 82829 59166 83209
rect 59178 82829 59558 83209
rect 67882 79370 68262 79750
rect 68274 79370 68654 79750
rect 68666 79370 69046 79750
rect 69058 79370 69438 79750
rect 69450 79370 69830 79750
rect 69842 79370 70222 79750
rect 70234 79370 70614 79750
rect 60042 74121 60422 74501
rect 60434 74121 60814 74501
rect 60826 74121 61206 74501
rect 61218 74121 61598 74501
rect 61610 74121 61990 74501
rect 62002 74121 62382 74501
rect 62394 74121 62774 74501
rect 62786 74121 63166 74501
rect 63178 74121 63558 74501
rect 60042 73729 60422 74109
rect 60434 73729 60814 74109
rect 60826 73729 61206 74109
rect 61218 73729 61598 74109
rect 61610 73729 61990 74109
rect 62002 73729 62382 74109
rect 62394 73729 62774 74109
rect 62786 73729 63166 74109
rect 63178 73729 63558 74109
rect 60042 73337 60422 73717
rect 60434 73337 60814 73717
rect 60826 73337 61206 73717
rect 61218 73337 61598 73717
rect 61610 73337 61990 73717
rect 62002 73337 62382 73717
rect 62394 73337 62774 73717
rect 62786 73337 63166 73717
rect 63178 73337 63558 73717
rect 60042 72945 60422 73325
rect 60434 72945 60814 73325
rect 60826 72945 61206 73325
rect 61218 72945 61598 73325
rect 61610 72945 61990 73325
rect 62002 72945 62382 73325
rect 62394 72945 62774 73325
rect 62786 72945 63166 73325
rect 63178 72945 63558 73325
rect 60042 72553 60422 72933
rect 60434 72553 60814 72933
rect 60826 72553 61206 72933
rect 61218 72553 61598 72933
rect 61610 72553 61990 72933
rect 62002 72553 62382 72933
rect 62394 72553 62774 72933
rect 62786 72553 63166 72933
rect 63178 72553 63558 72933
rect 60042 72161 60422 72541
rect 60434 72161 60814 72541
rect 60826 72161 61206 72541
rect 61218 72161 61598 72541
rect 61610 72161 61990 72541
rect 62002 72161 62382 72541
rect 62394 72161 62774 72541
rect 62786 72161 63166 72541
rect 63178 72161 63558 72541
rect 67882 74121 68262 74501
rect 68274 74121 68654 74501
rect 68666 74121 69046 74501
rect 69058 74121 69438 74501
rect 69450 74121 69830 74501
rect 69842 74121 70222 74501
rect 70234 74121 70614 74501
rect 67882 73729 68262 74109
rect 68274 73729 68654 74109
rect 68666 73729 69046 74109
rect 69058 73729 69438 74109
rect 69450 73729 69830 74109
rect 69842 73729 70222 74109
rect 70234 73729 70614 74109
rect 67882 73337 68262 73717
rect 68274 73337 68654 73717
rect 68666 73337 69046 73717
rect 69058 73337 69438 73717
rect 69450 73337 69830 73717
rect 69842 73337 70222 73717
rect 70234 73337 70614 73717
rect 67882 72945 68262 73325
rect 68274 72945 68654 73325
rect 68666 72945 69046 73325
rect 69058 72945 69438 73325
rect 69450 72945 69830 73325
rect 69842 72945 70222 73325
rect 70234 72945 70614 73325
rect 67882 72553 68262 72933
rect 68274 72553 68654 72933
rect 68666 72553 69046 72933
rect 69058 72553 69438 72933
rect 69450 72553 69830 72933
rect 69842 72553 70222 72933
rect 70234 72553 70614 72933
rect 67882 72161 68262 72541
rect 68274 72161 68654 72541
rect 68666 72161 69046 72541
rect 69058 72161 69438 72541
rect 69450 72161 69830 72541
rect 69842 72161 70222 72541
rect 70234 72161 70614 72541
rect 71882 151562 72262 151942
rect 72274 151562 72654 151942
rect 72666 151562 73046 151942
rect 73058 151562 73438 151942
rect 73450 151562 73830 151942
rect 73842 151562 74222 151942
rect 74234 151562 74614 151942
rect 71882 151170 72262 151550
rect 72274 151170 72654 151550
rect 72666 151170 73046 151550
rect 73058 151170 73438 151550
rect 73450 151170 73830 151550
rect 73842 151170 74222 151550
rect 74234 151170 74614 151550
rect 71882 150778 72262 151158
rect 72274 150778 72654 151158
rect 72666 150778 73046 151158
rect 73058 150778 73438 151158
rect 73450 150778 73830 151158
rect 73842 150778 74222 151158
rect 74234 150778 74614 151158
rect 71882 150386 72262 150766
rect 72274 150386 72654 150766
rect 72666 150386 73046 150766
rect 73058 150386 73438 150766
rect 73450 150386 73830 150766
rect 73842 150386 74222 150766
rect 74234 150386 74614 150766
rect 71882 149994 72262 150374
rect 72274 149994 72654 150374
rect 72666 149994 73046 150374
rect 73058 149994 73438 150374
rect 73450 149994 73830 150374
rect 73842 149994 74222 150374
rect 74234 149994 74614 150374
rect 71882 149602 72262 149982
rect 72274 149602 72654 149982
rect 72666 149602 73046 149982
rect 73058 149602 73438 149982
rect 73450 149602 73830 149982
rect 73842 149602 74222 149982
rect 74234 149602 74614 149982
rect 71882 149210 72262 149590
rect 72274 149210 72654 149590
rect 72666 149210 73046 149590
rect 73058 149210 73438 149590
rect 73450 149210 73830 149590
rect 73842 149210 74222 149590
rect 74234 149210 74614 149590
rect 71882 138610 72262 138990
rect 72274 138610 72654 138990
rect 72666 138610 73046 138990
rect 73058 138610 73438 138990
rect 73450 138610 73830 138990
rect 73842 138610 74222 138990
rect 74234 138610 74614 138990
rect 71882 132789 72262 133169
rect 72274 132789 72654 133169
rect 72666 132789 73046 133169
rect 73058 132789 73438 133169
rect 73450 132789 73830 133169
rect 73842 132789 74222 133169
rect 74234 132789 74614 133169
rect 71882 132397 72262 132777
rect 72274 132397 72654 132777
rect 72666 132397 73046 132777
rect 73058 132397 73438 132777
rect 73450 132397 73830 132777
rect 73842 132397 74222 132777
rect 74234 132397 74614 132777
rect 71882 132005 72262 132385
rect 72274 132005 72654 132385
rect 72666 132005 73046 132385
rect 73058 132005 73438 132385
rect 73450 132005 73830 132385
rect 73842 132005 74222 132385
rect 74234 132005 74614 132385
rect 71882 131613 72262 131993
rect 72274 131613 72654 131993
rect 72666 131613 73046 131993
rect 73058 131613 73438 131993
rect 73450 131613 73830 131993
rect 73842 131613 74222 131993
rect 74234 131613 74614 131993
rect 71882 131221 72262 131601
rect 72274 131221 72654 131601
rect 72666 131221 73046 131601
rect 73058 131221 73438 131601
rect 73450 131221 73830 131601
rect 73842 131221 74222 131601
rect 74234 131221 74614 131601
rect 71882 130829 72262 131209
rect 72274 130829 72654 131209
rect 72666 130829 73046 131209
rect 73058 130829 73438 131209
rect 73450 130829 73830 131209
rect 73842 130829 74222 131209
rect 74234 130829 74614 131209
rect 71882 123490 72262 123870
rect 72274 123490 72654 123870
rect 72666 123490 73046 123870
rect 73058 123490 73438 123870
rect 73450 123490 73830 123870
rect 73842 123490 74222 123870
rect 74234 123490 74614 123870
rect 71882 116789 72262 117169
rect 72274 116789 72654 117169
rect 72666 116789 73046 117169
rect 73058 116789 73438 117169
rect 73450 116789 73830 117169
rect 73842 116789 74222 117169
rect 74234 116789 74614 117169
rect 71882 116397 72262 116777
rect 72274 116397 72654 116777
rect 72666 116397 73046 116777
rect 73058 116397 73438 116777
rect 73450 116397 73830 116777
rect 73842 116397 74222 116777
rect 74234 116397 74614 116777
rect 71882 116005 72262 116385
rect 72274 116005 72654 116385
rect 72666 116005 73046 116385
rect 73058 116005 73438 116385
rect 73450 116005 73830 116385
rect 73842 116005 74222 116385
rect 74234 116005 74614 116385
rect 71882 115613 72262 115993
rect 72274 115613 72654 115993
rect 72666 115613 73046 115993
rect 73058 115613 73438 115993
rect 73450 115613 73830 115993
rect 73842 115613 74222 115993
rect 74234 115613 74614 115993
rect 71882 115221 72262 115601
rect 72274 115221 72654 115601
rect 72666 115221 73046 115601
rect 73058 115221 73438 115601
rect 73450 115221 73830 115601
rect 73842 115221 74222 115601
rect 74234 115221 74614 115601
rect 71882 114829 72262 115209
rect 72274 114829 72654 115209
rect 72666 114829 73046 115209
rect 73058 114829 73438 115209
rect 73450 114829 73830 115209
rect 73842 114829 74222 115209
rect 74234 114829 74614 115209
rect 71882 108370 72262 108750
rect 72274 108370 72654 108750
rect 72666 108370 73046 108750
rect 73058 108370 73438 108750
rect 73450 108370 73830 108750
rect 73842 108370 74222 108750
rect 74234 108370 74614 108750
rect 71882 100789 72262 101169
rect 72274 100789 72654 101169
rect 72666 100789 73046 101169
rect 73058 100789 73438 101169
rect 73450 100789 73830 101169
rect 73842 100789 74222 101169
rect 74234 100789 74614 101169
rect 71882 100397 72262 100777
rect 72274 100397 72654 100777
rect 72666 100397 73046 100777
rect 73058 100397 73438 100777
rect 73450 100397 73830 100777
rect 73842 100397 74222 100777
rect 74234 100397 74614 100777
rect 71882 100005 72262 100385
rect 72274 100005 72654 100385
rect 72666 100005 73046 100385
rect 73058 100005 73438 100385
rect 73450 100005 73830 100385
rect 73842 100005 74222 100385
rect 74234 100005 74614 100385
rect 71882 99613 72262 99993
rect 72274 99613 72654 99993
rect 72666 99613 73046 99993
rect 73058 99613 73438 99993
rect 73450 99613 73830 99993
rect 73842 99613 74222 99993
rect 74234 99613 74614 99993
rect 71882 99221 72262 99601
rect 72274 99221 72654 99601
rect 72666 99221 73046 99601
rect 73058 99221 73438 99601
rect 73450 99221 73830 99601
rect 73842 99221 74222 99601
rect 74234 99221 74614 99601
rect 71882 98829 72262 99209
rect 72274 98829 72654 99209
rect 72666 98829 73046 99209
rect 73058 98829 73438 99209
rect 73450 98829 73830 99209
rect 73842 98829 74222 99209
rect 74234 98829 74614 99209
rect 71882 93250 72262 93630
rect 72274 93250 72654 93630
rect 72666 93250 73046 93630
rect 73058 93250 73438 93630
rect 73450 93250 73830 93630
rect 73842 93250 74222 93630
rect 74234 93250 74614 93630
rect 71882 84789 72262 85169
rect 72274 84789 72654 85169
rect 72666 84789 73046 85169
rect 73058 84789 73438 85169
rect 73450 84789 73830 85169
rect 73842 84789 74222 85169
rect 74234 84789 74614 85169
rect 71882 84397 72262 84777
rect 72274 84397 72654 84777
rect 72666 84397 73046 84777
rect 73058 84397 73438 84777
rect 73450 84397 73830 84777
rect 73842 84397 74222 84777
rect 74234 84397 74614 84777
rect 71882 84005 72262 84385
rect 72274 84005 72654 84385
rect 72666 84005 73046 84385
rect 73058 84005 73438 84385
rect 73450 84005 73830 84385
rect 73842 84005 74222 84385
rect 74234 84005 74614 84385
rect 71882 83613 72262 83993
rect 72274 83613 72654 83993
rect 72666 83613 73046 83993
rect 73058 83613 73438 83993
rect 73450 83613 73830 83993
rect 73842 83613 74222 83993
rect 74234 83613 74614 83993
rect 71882 83221 72262 83601
rect 72274 83221 72654 83601
rect 72666 83221 73046 83601
rect 73058 83221 73438 83601
rect 73450 83221 73830 83601
rect 73842 83221 74222 83601
rect 74234 83221 74614 83601
rect 71882 82829 72262 83209
rect 72274 82829 72654 83209
rect 72666 82829 73046 83209
rect 73058 82829 73438 83209
rect 73450 82829 73830 83209
rect 73842 82829 74222 83209
rect 74234 82829 74614 83209
rect 71882 78130 72262 78510
rect 72274 78130 72654 78510
rect 72666 78130 73046 78510
rect 73058 78130 73438 78510
rect 73450 78130 73830 78510
rect 73842 78130 74222 78510
rect 74234 78130 74614 78510
rect 71882 74186 72262 74566
rect 72274 74186 72654 74566
rect 72666 74186 73046 74566
rect 73058 74186 73438 74566
rect 73450 74186 73830 74566
rect 73842 74186 74222 74566
rect 74234 74186 74614 74566
rect 71882 73794 72262 74174
rect 72274 73794 72654 74174
rect 72666 73794 73046 74174
rect 73058 73794 73438 74174
rect 73450 73794 73830 74174
rect 73842 73794 74222 74174
rect 74234 73794 74614 74174
rect 71882 73402 72262 73782
rect 72274 73402 72654 73782
rect 72666 73402 73046 73782
rect 73058 73402 73438 73782
rect 73450 73402 73830 73782
rect 73842 73402 74222 73782
rect 74234 73402 74614 73782
rect 71882 73010 72262 73390
rect 72274 73010 72654 73390
rect 72666 73010 73046 73390
rect 73058 73010 73438 73390
rect 73450 73010 73830 73390
rect 73842 73010 74222 73390
rect 74234 73010 74614 73390
rect 71882 72618 72262 72998
rect 72274 72618 72654 72998
rect 72666 72618 73046 72998
rect 73058 72618 73438 72998
rect 73450 72618 73830 72998
rect 73842 72618 74222 72998
rect 74234 72618 74614 72998
rect 71882 72226 72262 72606
rect 72274 72226 72654 72606
rect 72666 72226 73046 72606
rect 73058 72226 73438 72606
rect 73450 72226 73830 72606
rect 73842 72226 74222 72606
rect 74234 72226 74614 72606
rect 71882 71834 72262 72214
rect 72274 71834 72654 72214
rect 72666 71834 73046 72214
rect 73058 71834 73438 72214
rect 73450 71834 73830 72214
rect 73842 71834 74222 72214
rect 74234 71834 74614 72214
rect 78178 151562 78558 151942
rect 78178 151170 78558 151550
rect 78178 150778 78558 151158
rect 78178 150386 78558 150766
rect 78178 149994 78558 150374
rect 78178 149602 78558 149982
rect 78178 149210 78558 149590
rect 78178 138610 78558 138990
rect 78178 123490 78558 123870
rect 78178 108370 78558 108750
rect 78178 93250 78558 93630
rect 78178 78130 78558 78510
rect 78178 74186 78558 74566
rect 78178 73794 78558 74174
rect 78178 73402 78558 73782
rect 78178 73010 78558 73390
rect 78178 72618 78558 72998
rect 78178 72226 78558 72606
rect 78178 71834 78558 72214
rect 94538 155562 94918 155942
rect 94538 155170 94918 155550
rect 94538 154778 94918 155158
rect 94538 154386 94918 154766
rect 94538 153994 94918 154374
rect 94538 153602 94918 153982
rect 94538 153210 94918 153590
rect 79418 139850 79798 140230
rect 79418 124730 79798 125110
rect 79418 109610 79798 109990
rect 79418 94490 79798 94870
rect 79418 79370 79798 79750
rect 67882 70186 68262 70566
rect 68274 70186 68654 70566
rect 68666 70186 69046 70566
rect 69058 70186 69438 70566
rect 69450 70186 69830 70566
rect 69842 70186 70222 70566
rect 70234 70186 70614 70566
rect 67882 69794 68262 70174
rect 68274 69794 68654 70174
rect 68666 69794 69046 70174
rect 69058 69794 69438 70174
rect 69450 69794 69830 70174
rect 69842 69794 70222 70174
rect 70234 69794 70614 70174
rect 67882 69402 68262 69782
rect 68274 69402 68654 69782
rect 68666 69402 69046 69782
rect 69058 69402 69438 69782
rect 69450 69402 69830 69782
rect 69842 69402 70222 69782
rect 70234 69402 70614 69782
rect 67882 69010 68262 69390
rect 68274 69010 68654 69390
rect 68666 69010 69046 69390
rect 69058 69010 69438 69390
rect 69450 69010 69830 69390
rect 69842 69010 70222 69390
rect 70234 69010 70614 69390
rect 67882 68618 68262 68998
rect 68274 68618 68654 68998
rect 68666 68618 69046 68998
rect 69058 68618 69438 68998
rect 69450 68618 69830 68998
rect 69842 68618 70222 68998
rect 70234 68618 70614 68998
rect 67882 68226 68262 68606
rect 68274 68226 68654 68606
rect 68666 68226 69046 68606
rect 69058 68226 69438 68606
rect 69450 68226 69830 68606
rect 69842 68226 70222 68606
rect 70234 68226 70614 68606
rect 67882 67834 68262 68214
rect 68274 67834 68654 68214
rect 68666 67834 69046 68214
rect 69058 67834 69438 68214
rect 69450 67834 69830 68214
rect 69842 67834 70222 68214
rect 70234 67834 70614 68214
rect 93298 151562 93678 151942
rect 93298 151170 93678 151550
rect 93298 150778 93678 151158
rect 93298 150386 93678 150766
rect 93298 149994 93678 150374
rect 93298 149602 93678 149982
rect 93298 149210 93678 149590
rect 93298 138610 93678 138990
rect 93298 123490 93678 123870
rect 93298 108370 93678 108750
rect 93298 93250 93678 93630
rect 93298 78130 93678 78510
rect 93298 74186 93678 74566
rect 93298 73794 93678 74174
rect 93298 73402 93678 73782
rect 93298 73010 93678 73390
rect 93298 72618 93678 72998
rect 93298 72226 93678 72606
rect 93298 71834 93678 72214
rect 109658 155562 110038 155942
rect 109658 155170 110038 155550
rect 109658 154778 110038 155158
rect 109658 154386 110038 154766
rect 109658 153994 110038 154374
rect 109658 153602 110038 153982
rect 109658 153210 110038 153590
rect 94538 139850 94918 140230
rect 94538 124730 94918 125110
rect 94538 109610 94918 109990
rect 94538 94490 94918 94870
rect 94538 79370 94918 79750
rect 79418 70186 79798 70566
rect 79418 69794 79798 70174
rect 79418 69402 79798 69782
rect 79418 69010 79798 69390
rect 79418 68618 79798 68998
rect 79418 68226 79798 68606
rect 79418 67834 79798 68214
rect 108418 151562 108798 151942
rect 108418 151170 108798 151550
rect 108418 150778 108798 151158
rect 108418 150386 108798 150766
rect 108418 149994 108798 150374
rect 108418 149602 108798 149982
rect 108418 149210 108798 149590
rect 108418 138610 108798 138990
rect 108418 123490 108798 123870
rect 108418 108370 108798 108750
rect 108418 93250 108798 93630
rect 108418 78130 108798 78510
rect 108418 74186 108798 74566
rect 108418 73794 108798 74174
rect 108418 73402 108798 73782
rect 108418 73010 108798 73390
rect 108418 72618 108798 72998
rect 108418 72226 108798 72606
rect 108418 71834 108798 72214
rect 124778 155562 125158 155942
rect 124778 155170 125158 155550
rect 124778 154778 125158 155158
rect 124778 154386 125158 154766
rect 124778 153994 125158 154374
rect 124778 153602 125158 153982
rect 124778 153210 125158 153590
rect 109658 139850 110038 140230
rect 109658 124730 110038 125110
rect 109658 109610 110038 109990
rect 109658 94490 110038 94870
rect 109658 79370 110038 79750
rect 94538 70186 94918 70566
rect 94538 69794 94918 70174
rect 94538 69402 94918 69782
rect 94538 69010 94918 69390
rect 94538 68618 94918 68998
rect 94538 68226 94918 68606
rect 94538 67834 94918 68214
rect 123538 151562 123918 151942
rect 123538 151170 123918 151550
rect 123538 150778 123918 151158
rect 123538 150386 123918 150766
rect 123538 149994 123918 150374
rect 123538 149602 123918 149982
rect 123538 149210 123918 149590
rect 123538 138610 123918 138990
rect 123538 123490 123918 123870
rect 123538 108370 123918 108750
rect 123538 93250 123918 93630
rect 123538 78130 123918 78510
rect 123538 74186 123918 74566
rect 123538 73794 123918 74174
rect 123538 73402 123918 73782
rect 123538 73010 123918 73390
rect 123538 72618 123918 72998
rect 123538 72226 123918 72606
rect 123538 71834 123918 72214
rect 139898 155562 140278 155942
rect 139898 155170 140278 155550
rect 139898 154778 140278 155158
rect 139898 154386 140278 154766
rect 139898 153994 140278 154374
rect 139898 153602 140278 153982
rect 139898 153210 140278 153590
rect 124778 139850 125158 140230
rect 124778 124730 125158 125110
rect 124778 109610 125158 109990
rect 124778 94490 125158 94870
rect 124778 79370 125158 79750
rect 109658 70186 110038 70566
rect 109658 69794 110038 70174
rect 109658 69402 110038 69782
rect 109658 69010 110038 69390
rect 109658 68618 110038 68998
rect 109658 68226 110038 68606
rect 109658 67834 110038 68214
rect 138658 151562 139038 151942
rect 138658 151170 139038 151550
rect 138658 150778 139038 151158
rect 138658 150386 139038 150766
rect 138658 149994 139038 150374
rect 138658 149602 139038 149982
rect 138658 149210 139038 149590
rect 138658 138610 139038 138990
rect 138658 123490 139038 123870
rect 138658 108370 139038 108750
rect 138658 93250 139038 93630
rect 138658 78130 139038 78510
rect 138658 74186 139038 74566
rect 138658 73794 139038 74174
rect 138658 73402 139038 73782
rect 138658 73010 139038 73390
rect 138658 72618 139038 72998
rect 138658 72226 139038 72606
rect 138658 71834 139038 72214
rect 153354 155562 153734 155942
rect 153746 155562 154126 155942
rect 154138 155562 154518 155942
rect 154530 155562 154910 155942
rect 154922 155562 155302 155942
rect 155314 155562 155694 155942
rect 155706 155562 156086 155942
rect 153354 155170 153734 155550
rect 153746 155170 154126 155550
rect 154138 155170 154518 155550
rect 154530 155170 154910 155550
rect 154922 155170 155302 155550
rect 155314 155170 155694 155550
rect 155706 155170 156086 155550
rect 153354 154778 153734 155158
rect 153746 154778 154126 155158
rect 154138 154778 154518 155158
rect 154530 154778 154910 155158
rect 154922 154778 155302 155158
rect 155314 154778 155694 155158
rect 155706 154778 156086 155158
rect 153354 154386 153734 154766
rect 153746 154386 154126 154766
rect 154138 154386 154518 154766
rect 154530 154386 154910 154766
rect 154922 154386 155302 154766
rect 155314 154386 155694 154766
rect 155706 154386 156086 154766
rect 153354 153994 153734 154374
rect 153746 153994 154126 154374
rect 154138 153994 154518 154374
rect 154530 153994 154910 154374
rect 154922 153994 155302 154374
rect 155314 153994 155694 154374
rect 155706 153994 156086 154374
rect 153354 153602 153734 153982
rect 153746 153602 154126 153982
rect 154138 153602 154518 153982
rect 154530 153602 154910 153982
rect 154922 153602 155302 153982
rect 155314 153602 155694 153982
rect 155706 153602 156086 153982
rect 153354 153210 153734 153590
rect 153746 153210 154126 153590
rect 154138 153210 154518 153590
rect 154530 153210 154910 153590
rect 154922 153210 155302 153590
rect 155314 153210 155694 153590
rect 155706 153210 156086 153590
rect 139898 139850 140278 140230
rect 139898 124730 140278 125110
rect 139898 109610 140278 109990
rect 139898 94490 140278 94870
rect 139898 79370 140278 79750
rect 124778 70186 125158 70566
rect 124778 69794 125158 70174
rect 124778 69402 125158 69782
rect 124778 69010 125158 69390
rect 124778 68618 125158 68998
rect 124778 68226 125158 68606
rect 124778 67834 125158 68214
rect 149354 151562 149734 151942
rect 149746 151562 150126 151942
rect 150138 151562 150518 151942
rect 150530 151562 150910 151942
rect 150922 151562 151302 151942
rect 151314 151562 151694 151942
rect 151706 151562 152086 151942
rect 149354 151170 149734 151550
rect 149746 151170 150126 151550
rect 150138 151170 150518 151550
rect 150530 151170 150910 151550
rect 150922 151170 151302 151550
rect 151314 151170 151694 151550
rect 151706 151170 152086 151550
rect 149354 150778 149734 151158
rect 149746 150778 150126 151158
rect 150138 150778 150518 151158
rect 150530 150778 150910 151158
rect 150922 150778 151302 151158
rect 151314 150778 151694 151158
rect 151706 150778 152086 151158
rect 149354 150386 149734 150766
rect 149746 150386 150126 150766
rect 150138 150386 150518 150766
rect 150530 150386 150910 150766
rect 150922 150386 151302 150766
rect 151314 150386 151694 150766
rect 151706 150386 152086 150766
rect 149354 149994 149734 150374
rect 149746 149994 150126 150374
rect 150138 149994 150518 150374
rect 150530 149994 150910 150374
rect 150922 149994 151302 150374
rect 151314 149994 151694 150374
rect 151706 149994 152086 150374
rect 149354 149602 149734 149982
rect 149746 149602 150126 149982
rect 150138 149602 150518 149982
rect 150530 149602 150910 149982
rect 150922 149602 151302 149982
rect 151314 149602 151694 149982
rect 151706 149602 152086 149982
rect 149354 149210 149734 149590
rect 149746 149210 150126 149590
rect 150138 149210 150518 149590
rect 150530 149210 150910 149590
rect 150922 149210 151302 149590
rect 151314 149210 151694 149590
rect 151706 149210 152086 149590
rect 149354 138610 149734 138990
rect 149746 138610 150126 138990
rect 150138 138610 150518 138990
rect 150530 138610 150910 138990
rect 150922 138610 151302 138990
rect 151314 138610 151694 138990
rect 151706 138610 152086 138990
rect 149354 132789 149734 133169
rect 149746 132789 150126 133169
rect 150138 132789 150518 133169
rect 150530 132789 150910 133169
rect 150922 132789 151302 133169
rect 151314 132789 151694 133169
rect 151706 132789 152086 133169
rect 149354 132397 149734 132777
rect 149746 132397 150126 132777
rect 150138 132397 150518 132777
rect 150530 132397 150910 132777
rect 150922 132397 151302 132777
rect 151314 132397 151694 132777
rect 151706 132397 152086 132777
rect 149354 132005 149734 132385
rect 149746 132005 150126 132385
rect 150138 132005 150518 132385
rect 150530 132005 150910 132385
rect 150922 132005 151302 132385
rect 151314 132005 151694 132385
rect 151706 132005 152086 132385
rect 149354 131613 149734 131993
rect 149746 131613 150126 131993
rect 150138 131613 150518 131993
rect 150530 131613 150910 131993
rect 150922 131613 151302 131993
rect 151314 131613 151694 131993
rect 151706 131613 152086 131993
rect 149354 131221 149734 131601
rect 149746 131221 150126 131601
rect 150138 131221 150518 131601
rect 150530 131221 150910 131601
rect 150922 131221 151302 131601
rect 151314 131221 151694 131601
rect 151706 131221 152086 131601
rect 149354 130829 149734 131209
rect 149746 130829 150126 131209
rect 150138 130829 150518 131209
rect 150530 130829 150910 131209
rect 150922 130829 151302 131209
rect 151314 130829 151694 131209
rect 151706 130829 152086 131209
rect 149354 123490 149734 123870
rect 149746 123490 150126 123870
rect 150138 123490 150518 123870
rect 150530 123490 150910 123870
rect 150922 123490 151302 123870
rect 151314 123490 151694 123870
rect 151706 123490 152086 123870
rect 149354 116789 149734 117169
rect 149746 116789 150126 117169
rect 150138 116789 150518 117169
rect 150530 116789 150910 117169
rect 150922 116789 151302 117169
rect 151314 116789 151694 117169
rect 151706 116789 152086 117169
rect 149354 116397 149734 116777
rect 149746 116397 150126 116777
rect 150138 116397 150518 116777
rect 150530 116397 150910 116777
rect 150922 116397 151302 116777
rect 151314 116397 151694 116777
rect 151706 116397 152086 116777
rect 149354 116005 149734 116385
rect 149746 116005 150126 116385
rect 150138 116005 150518 116385
rect 150530 116005 150910 116385
rect 150922 116005 151302 116385
rect 151314 116005 151694 116385
rect 151706 116005 152086 116385
rect 149354 115613 149734 115993
rect 149746 115613 150126 115993
rect 150138 115613 150518 115993
rect 150530 115613 150910 115993
rect 150922 115613 151302 115993
rect 151314 115613 151694 115993
rect 151706 115613 152086 115993
rect 149354 115221 149734 115601
rect 149746 115221 150126 115601
rect 150138 115221 150518 115601
rect 150530 115221 150910 115601
rect 150922 115221 151302 115601
rect 151314 115221 151694 115601
rect 151706 115221 152086 115601
rect 149354 114829 149734 115209
rect 149746 114829 150126 115209
rect 150138 114829 150518 115209
rect 150530 114829 150910 115209
rect 150922 114829 151302 115209
rect 151314 114829 151694 115209
rect 151706 114829 152086 115209
rect 149354 108370 149734 108750
rect 149746 108370 150126 108750
rect 150138 108370 150518 108750
rect 150530 108370 150910 108750
rect 150922 108370 151302 108750
rect 151314 108370 151694 108750
rect 151706 108370 152086 108750
rect 149354 100789 149734 101169
rect 149746 100789 150126 101169
rect 150138 100789 150518 101169
rect 150530 100789 150910 101169
rect 150922 100789 151302 101169
rect 151314 100789 151694 101169
rect 151706 100789 152086 101169
rect 149354 100397 149734 100777
rect 149746 100397 150126 100777
rect 150138 100397 150518 100777
rect 150530 100397 150910 100777
rect 150922 100397 151302 100777
rect 151314 100397 151694 100777
rect 151706 100397 152086 100777
rect 149354 100005 149734 100385
rect 149746 100005 150126 100385
rect 150138 100005 150518 100385
rect 150530 100005 150910 100385
rect 150922 100005 151302 100385
rect 151314 100005 151694 100385
rect 151706 100005 152086 100385
rect 149354 99613 149734 99993
rect 149746 99613 150126 99993
rect 150138 99613 150518 99993
rect 150530 99613 150910 99993
rect 150922 99613 151302 99993
rect 151314 99613 151694 99993
rect 151706 99613 152086 99993
rect 149354 99221 149734 99601
rect 149746 99221 150126 99601
rect 150138 99221 150518 99601
rect 150530 99221 150910 99601
rect 150922 99221 151302 99601
rect 151314 99221 151694 99601
rect 151706 99221 152086 99601
rect 149354 98829 149734 99209
rect 149746 98829 150126 99209
rect 150138 98829 150518 99209
rect 150530 98829 150910 99209
rect 150922 98829 151302 99209
rect 151314 98829 151694 99209
rect 151706 98829 152086 99209
rect 149354 93250 149734 93630
rect 149746 93250 150126 93630
rect 150138 93250 150518 93630
rect 150530 93250 150910 93630
rect 150922 93250 151302 93630
rect 151314 93250 151694 93630
rect 151706 93250 152086 93630
rect 149354 84789 149734 85169
rect 149746 84789 150126 85169
rect 150138 84789 150518 85169
rect 150530 84789 150910 85169
rect 150922 84789 151302 85169
rect 151314 84789 151694 85169
rect 151706 84789 152086 85169
rect 149354 84397 149734 84777
rect 149746 84397 150126 84777
rect 150138 84397 150518 84777
rect 150530 84397 150910 84777
rect 150922 84397 151302 84777
rect 151314 84397 151694 84777
rect 151706 84397 152086 84777
rect 149354 84005 149734 84385
rect 149746 84005 150126 84385
rect 150138 84005 150518 84385
rect 150530 84005 150910 84385
rect 150922 84005 151302 84385
rect 151314 84005 151694 84385
rect 151706 84005 152086 84385
rect 149354 83613 149734 83993
rect 149746 83613 150126 83993
rect 150138 83613 150518 83993
rect 150530 83613 150910 83993
rect 150922 83613 151302 83993
rect 151314 83613 151694 83993
rect 151706 83613 152086 83993
rect 149354 83221 149734 83601
rect 149746 83221 150126 83601
rect 150138 83221 150518 83601
rect 150530 83221 150910 83601
rect 150922 83221 151302 83601
rect 151314 83221 151694 83601
rect 151706 83221 152086 83601
rect 149354 82829 149734 83209
rect 149746 82829 150126 83209
rect 150138 82829 150518 83209
rect 150530 82829 150910 83209
rect 150922 82829 151302 83209
rect 151314 82829 151694 83209
rect 151706 82829 152086 83209
rect 149354 78130 149734 78510
rect 149746 78130 150126 78510
rect 150138 78130 150518 78510
rect 150530 78130 150910 78510
rect 150922 78130 151302 78510
rect 151314 78130 151694 78510
rect 151706 78130 152086 78510
rect 149354 74186 149734 74566
rect 149746 74186 150126 74566
rect 150138 74186 150518 74566
rect 150530 74186 150910 74566
rect 150922 74186 151302 74566
rect 151314 74186 151694 74566
rect 151706 74186 152086 74566
rect 149354 73794 149734 74174
rect 149746 73794 150126 74174
rect 150138 73794 150518 74174
rect 150530 73794 150910 74174
rect 150922 73794 151302 74174
rect 151314 73794 151694 74174
rect 151706 73794 152086 74174
rect 149354 73402 149734 73782
rect 149746 73402 150126 73782
rect 150138 73402 150518 73782
rect 150530 73402 150910 73782
rect 150922 73402 151302 73782
rect 151314 73402 151694 73782
rect 151706 73402 152086 73782
rect 149354 73010 149734 73390
rect 149746 73010 150126 73390
rect 150138 73010 150518 73390
rect 150530 73010 150910 73390
rect 150922 73010 151302 73390
rect 151314 73010 151694 73390
rect 151706 73010 152086 73390
rect 149354 72618 149734 72998
rect 149746 72618 150126 72998
rect 150138 72618 150518 72998
rect 150530 72618 150910 72998
rect 150922 72618 151302 72998
rect 151314 72618 151694 72998
rect 151706 72618 152086 72998
rect 149354 72226 149734 72606
rect 149746 72226 150126 72606
rect 150138 72226 150518 72606
rect 150530 72226 150910 72606
rect 150922 72226 151302 72606
rect 151314 72226 151694 72606
rect 151706 72226 152086 72606
rect 149354 71834 149734 72214
rect 149746 71834 150126 72214
rect 150138 71834 150518 72214
rect 150530 71834 150910 72214
rect 150922 71834 151302 72214
rect 151314 71834 151694 72214
rect 151706 71834 152086 72214
rect 153354 139850 153734 140230
rect 153746 139850 154126 140230
rect 154138 139850 154518 140230
rect 154530 139850 154910 140230
rect 154922 139850 155302 140230
rect 155314 139850 155694 140230
rect 155706 139850 156086 140230
rect 164442 132789 164822 133169
rect 164834 132789 165214 133169
rect 165226 132789 165606 133169
rect 165618 132789 165998 133169
rect 166010 132789 166390 133169
rect 166402 132789 166782 133169
rect 166794 132789 167174 133169
rect 167186 132789 167566 133169
rect 167578 132789 167958 133169
rect 164442 132397 164822 132777
rect 164834 132397 165214 132777
rect 165226 132397 165606 132777
rect 165618 132397 165998 132777
rect 166010 132397 166390 132777
rect 166402 132397 166782 132777
rect 166794 132397 167174 132777
rect 167186 132397 167566 132777
rect 167578 132397 167958 132777
rect 164442 132005 164822 132385
rect 164834 132005 165214 132385
rect 165226 132005 165606 132385
rect 165618 132005 165998 132385
rect 166010 132005 166390 132385
rect 166402 132005 166782 132385
rect 166794 132005 167174 132385
rect 167186 132005 167566 132385
rect 167578 132005 167958 132385
rect 164442 131613 164822 131993
rect 164834 131613 165214 131993
rect 165226 131613 165606 131993
rect 165618 131613 165998 131993
rect 166010 131613 166390 131993
rect 166402 131613 166782 131993
rect 166794 131613 167174 131993
rect 167186 131613 167566 131993
rect 167578 131613 167958 131993
rect 164442 131221 164822 131601
rect 164834 131221 165214 131601
rect 165226 131221 165606 131601
rect 165618 131221 165998 131601
rect 166010 131221 166390 131601
rect 166402 131221 166782 131601
rect 166794 131221 167174 131601
rect 167186 131221 167566 131601
rect 167578 131221 167958 131601
rect 164442 130829 164822 131209
rect 164834 130829 165214 131209
rect 165226 130829 165606 131209
rect 165618 130829 165998 131209
rect 166010 130829 166390 131209
rect 166402 130829 166782 131209
rect 166794 130829 167174 131209
rect 167186 130829 167566 131209
rect 167578 130829 167958 131209
rect 153354 124730 153734 125110
rect 153746 124730 154126 125110
rect 154138 124730 154518 125110
rect 154530 124730 154910 125110
rect 154922 124730 155302 125110
rect 155314 124730 155694 125110
rect 155706 124730 156086 125110
rect 164442 116789 164822 117169
rect 164834 116789 165214 117169
rect 165226 116789 165606 117169
rect 165618 116789 165998 117169
rect 166010 116789 166390 117169
rect 166402 116789 166782 117169
rect 166794 116789 167174 117169
rect 167186 116789 167566 117169
rect 167578 116789 167958 117169
rect 164442 116397 164822 116777
rect 164834 116397 165214 116777
rect 165226 116397 165606 116777
rect 165618 116397 165998 116777
rect 166010 116397 166390 116777
rect 166402 116397 166782 116777
rect 166794 116397 167174 116777
rect 167186 116397 167566 116777
rect 167578 116397 167958 116777
rect 164442 116005 164822 116385
rect 164834 116005 165214 116385
rect 165226 116005 165606 116385
rect 165618 116005 165998 116385
rect 166010 116005 166390 116385
rect 166402 116005 166782 116385
rect 166794 116005 167174 116385
rect 167186 116005 167566 116385
rect 167578 116005 167958 116385
rect 164442 115613 164822 115993
rect 164834 115613 165214 115993
rect 165226 115613 165606 115993
rect 165618 115613 165998 115993
rect 166010 115613 166390 115993
rect 166402 115613 166782 115993
rect 166794 115613 167174 115993
rect 167186 115613 167566 115993
rect 167578 115613 167958 115993
rect 164442 115221 164822 115601
rect 164834 115221 165214 115601
rect 165226 115221 165606 115601
rect 165618 115221 165998 115601
rect 166010 115221 166390 115601
rect 166402 115221 166782 115601
rect 166794 115221 167174 115601
rect 167186 115221 167566 115601
rect 167578 115221 167958 115601
rect 164442 114829 164822 115209
rect 164834 114829 165214 115209
rect 165226 114829 165606 115209
rect 165618 114829 165998 115209
rect 166010 114829 166390 115209
rect 166402 114829 166782 115209
rect 166794 114829 167174 115209
rect 167186 114829 167566 115209
rect 167578 114829 167958 115209
rect 153354 109610 153734 109990
rect 153746 109610 154126 109990
rect 154138 109610 154518 109990
rect 154530 109610 154910 109990
rect 154922 109610 155302 109990
rect 155314 109610 155694 109990
rect 155706 109610 156086 109990
rect 153354 106121 153734 106501
rect 153746 106121 154126 106501
rect 154138 106121 154518 106501
rect 154530 106121 154910 106501
rect 154922 106121 155302 106501
rect 155314 106121 155694 106501
rect 155706 106121 156086 106501
rect 153354 105729 153734 106109
rect 153746 105729 154126 106109
rect 154138 105729 154518 106109
rect 154530 105729 154910 106109
rect 154922 105729 155302 106109
rect 155314 105729 155694 106109
rect 155706 105729 156086 106109
rect 153354 105337 153734 105717
rect 153746 105337 154126 105717
rect 154138 105337 154518 105717
rect 154530 105337 154910 105717
rect 154922 105337 155302 105717
rect 155314 105337 155694 105717
rect 155706 105337 156086 105717
rect 153354 104945 153734 105325
rect 153746 104945 154126 105325
rect 154138 104945 154518 105325
rect 154530 104945 154910 105325
rect 154922 104945 155302 105325
rect 155314 104945 155694 105325
rect 155706 104945 156086 105325
rect 153354 104553 153734 104933
rect 153746 104553 154126 104933
rect 154138 104553 154518 104933
rect 154530 104553 154910 104933
rect 154922 104553 155302 104933
rect 155314 104553 155694 104933
rect 155706 104553 156086 104933
rect 153354 104161 153734 104541
rect 153746 104161 154126 104541
rect 154138 104161 154518 104541
rect 154530 104161 154910 104541
rect 154922 104161 155302 104541
rect 155314 104161 155694 104541
rect 155706 104161 156086 104541
rect 160442 106121 160822 106501
rect 160834 106121 161214 106501
rect 161226 106121 161606 106501
rect 161618 106121 161998 106501
rect 162010 106121 162390 106501
rect 162402 106121 162782 106501
rect 162794 106121 163174 106501
rect 163186 106121 163566 106501
rect 163578 106121 163958 106501
rect 160442 105729 160822 106109
rect 160834 105729 161214 106109
rect 161226 105729 161606 106109
rect 161618 105729 161998 106109
rect 162010 105729 162390 106109
rect 162402 105729 162782 106109
rect 162794 105729 163174 106109
rect 163186 105729 163566 106109
rect 163578 105729 163958 106109
rect 160442 105337 160822 105717
rect 160834 105337 161214 105717
rect 161226 105337 161606 105717
rect 161618 105337 161998 105717
rect 162010 105337 162390 105717
rect 162402 105337 162782 105717
rect 162794 105337 163174 105717
rect 163186 105337 163566 105717
rect 163578 105337 163958 105717
rect 160442 104945 160822 105325
rect 160834 104945 161214 105325
rect 161226 104945 161606 105325
rect 161618 104945 161998 105325
rect 162010 104945 162390 105325
rect 162402 104945 162782 105325
rect 162794 104945 163174 105325
rect 163186 104945 163566 105325
rect 163578 104945 163958 105325
rect 160442 104553 160822 104933
rect 160834 104553 161214 104933
rect 161226 104553 161606 104933
rect 161618 104553 161998 104933
rect 162010 104553 162390 104933
rect 162402 104553 162782 104933
rect 162794 104553 163174 104933
rect 163186 104553 163566 104933
rect 163578 104553 163958 104933
rect 160442 104161 160822 104541
rect 160834 104161 161214 104541
rect 161226 104161 161606 104541
rect 161618 104161 161998 104541
rect 162010 104161 162390 104541
rect 162402 104161 162782 104541
rect 162794 104161 163174 104541
rect 163186 104161 163566 104541
rect 163578 104161 163958 104541
rect 164442 100789 164822 101169
rect 164834 100789 165214 101169
rect 165226 100789 165606 101169
rect 165618 100789 165998 101169
rect 166010 100789 166390 101169
rect 166402 100789 166782 101169
rect 166794 100789 167174 101169
rect 167186 100789 167566 101169
rect 167578 100789 167958 101169
rect 164442 100397 164822 100777
rect 164834 100397 165214 100777
rect 165226 100397 165606 100777
rect 165618 100397 165998 100777
rect 166010 100397 166390 100777
rect 166402 100397 166782 100777
rect 166794 100397 167174 100777
rect 167186 100397 167566 100777
rect 167578 100397 167958 100777
rect 164442 100005 164822 100385
rect 164834 100005 165214 100385
rect 165226 100005 165606 100385
rect 165618 100005 165998 100385
rect 166010 100005 166390 100385
rect 166402 100005 166782 100385
rect 166794 100005 167174 100385
rect 167186 100005 167566 100385
rect 167578 100005 167958 100385
rect 164442 99613 164822 99993
rect 164834 99613 165214 99993
rect 165226 99613 165606 99993
rect 165618 99613 165998 99993
rect 166010 99613 166390 99993
rect 166402 99613 166782 99993
rect 166794 99613 167174 99993
rect 167186 99613 167566 99993
rect 167578 99613 167958 99993
rect 164442 99221 164822 99601
rect 164834 99221 165214 99601
rect 165226 99221 165606 99601
rect 165618 99221 165998 99601
rect 166010 99221 166390 99601
rect 166402 99221 166782 99601
rect 166794 99221 167174 99601
rect 167186 99221 167566 99601
rect 167578 99221 167958 99601
rect 164442 98829 164822 99209
rect 164834 98829 165214 99209
rect 165226 98829 165606 99209
rect 165618 98829 165998 99209
rect 166010 98829 166390 99209
rect 166402 98829 166782 99209
rect 166794 98829 167174 99209
rect 167186 98829 167566 99209
rect 167578 98829 167958 99209
rect 153354 94490 153734 94870
rect 153746 94490 154126 94870
rect 154138 94490 154518 94870
rect 154530 94490 154910 94870
rect 154922 94490 155302 94870
rect 155314 94490 155694 94870
rect 155706 94490 156086 94870
rect 153354 90121 153734 90501
rect 153746 90121 154126 90501
rect 154138 90121 154518 90501
rect 154530 90121 154910 90501
rect 154922 90121 155302 90501
rect 155314 90121 155694 90501
rect 155706 90121 156086 90501
rect 153354 89729 153734 90109
rect 153746 89729 154126 90109
rect 154138 89729 154518 90109
rect 154530 89729 154910 90109
rect 154922 89729 155302 90109
rect 155314 89729 155694 90109
rect 155706 89729 156086 90109
rect 153354 89337 153734 89717
rect 153746 89337 154126 89717
rect 154138 89337 154518 89717
rect 154530 89337 154910 89717
rect 154922 89337 155302 89717
rect 155314 89337 155694 89717
rect 155706 89337 156086 89717
rect 153354 88945 153734 89325
rect 153746 88945 154126 89325
rect 154138 88945 154518 89325
rect 154530 88945 154910 89325
rect 154922 88945 155302 89325
rect 155314 88945 155694 89325
rect 155706 88945 156086 89325
rect 153354 88553 153734 88933
rect 153746 88553 154126 88933
rect 154138 88553 154518 88933
rect 154530 88553 154910 88933
rect 154922 88553 155302 88933
rect 155314 88553 155694 88933
rect 155706 88553 156086 88933
rect 153354 88161 153734 88541
rect 153746 88161 154126 88541
rect 154138 88161 154518 88541
rect 154530 88161 154910 88541
rect 154922 88161 155302 88541
rect 155314 88161 155694 88541
rect 155706 88161 156086 88541
rect 160442 90121 160822 90501
rect 160834 90121 161214 90501
rect 161226 90121 161606 90501
rect 161618 90121 161998 90501
rect 162010 90121 162390 90501
rect 162402 90121 162782 90501
rect 162794 90121 163174 90501
rect 163186 90121 163566 90501
rect 163578 90121 163958 90501
rect 160442 89729 160822 90109
rect 160834 89729 161214 90109
rect 161226 89729 161606 90109
rect 161618 89729 161998 90109
rect 162010 89729 162390 90109
rect 162402 89729 162782 90109
rect 162794 89729 163174 90109
rect 163186 89729 163566 90109
rect 163578 89729 163958 90109
rect 160442 89337 160822 89717
rect 160834 89337 161214 89717
rect 161226 89337 161606 89717
rect 161618 89337 161998 89717
rect 162010 89337 162390 89717
rect 162402 89337 162782 89717
rect 162794 89337 163174 89717
rect 163186 89337 163566 89717
rect 163578 89337 163958 89717
rect 160442 88945 160822 89325
rect 160834 88945 161214 89325
rect 161226 88945 161606 89325
rect 161618 88945 161998 89325
rect 162010 88945 162390 89325
rect 162402 88945 162782 89325
rect 162794 88945 163174 89325
rect 163186 88945 163566 89325
rect 163578 88945 163958 89325
rect 160442 88553 160822 88933
rect 160834 88553 161214 88933
rect 161226 88553 161606 88933
rect 161618 88553 161998 88933
rect 162010 88553 162390 88933
rect 162402 88553 162782 88933
rect 162794 88553 163174 88933
rect 163186 88553 163566 88933
rect 163578 88553 163958 88933
rect 160442 88161 160822 88541
rect 160834 88161 161214 88541
rect 161226 88161 161606 88541
rect 161618 88161 161998 88541
rect 162010 88161 162390 88541
rect 162402 88161 162782 88541
rect 162794 88161 163174 88541
rect 163186 88161 163566 88541
rect 163578 88161 163958 88541
rect 164442 84789 164822 85169
rect 164834 84789 165214 85169
rect 165226 84789 165606 85169
rect 165618 84789 165998 85169
rect 166010 84789 166390 85169
rect 166402 84789 166782 85169
rect 166794 84789 167174 85169
rect 167186 84789 167566 85169
rect 167578 84789 167958 85169
rect 164442 84397 164822 84777
rect 164834 84397 165214 84777
rect 165226 84397 165606 84777
rect 165618 84397 165998 84777
rect 166010 84397 166390 84777
rect 166402 84397 166782 84777
rect 166794 84397 167174 84777
rect 167186 84397 167566 84777
rect 167578 84397 167958 84777
rect 164442 84005 164822 84385
rect 164834 84005 165214 84385
rect 165226 84005 165606 84385
rect 165618 84005 165998 84385
rect 166010 84005 166390 84385
rect 166402 84005 166782 84385
rect 166794 84005 167174 84385
rect 167186 84005 167566 84385
rect 167578 84005 167958 84385
rect 164442 83613 164822 83993
rect 164834 83613 165214 83993
rect 165226 83613 165606 83993
rect 165618 83613 165998 83993
rect 166010 83613 166390 83993
rect 166402 83613 166782 83993
rect 166794 83613 167174 83993
rect 167186 83613 167566 83993
rect 167578 83613 167958 83993
rect 164442 83221 164822 83601
rect 164834 83221 165214 83601
rect 165226 83221 165606 83601
rect 165618 83221 165998 83601
rect 166010 83221 166390 83601
rect 166402 83221 166782 83601
rect 166794 83221 167174 83601
rect 167186 83221 167566 83601
rect 167578 83221 167958 83601
rect 164442 82829 164822 83209
rect 164834 82829 165214 83209
rect 165226 82829 165606 83209
rect 165618 82829 165998 83209
rect 166010 82829 166390 83209
rect 166402 82829 166782 83209
rect 166794 82829 167174 83209
rect 167186 82829 167566 83209
rect 167578 82829 167958 83209
rect 153354 79370 153734 79750
rect 153746 79370 154126 79750
rect 154138 79370 154518 79750
rect 154530 79370 154910 79750
rect 154922 79370 155302 79750
rect 155314 79370 155694 79750
rect 155706 79370 156086 79750
rect 153354 74121 153734 74501
rect 153746 74121 154126 74501
rect 154138 74121 154518 74501
rect 154530 74121 154910 74501
rect 154922 74121 155302 74501
rect 155314 74121 155694 74501
rect 155706 74121 156086 74501
rect 153354 73729 153734 74109
rect 153746 73729 154126 74109
rect 154138 73729 154518 74109
rect 154530 73729 154910 74109
rect 154922 73729 155302 74109
rect 155314 73729 155694 74109
rect 155706 73729 156086 74109
rect 153354 73337 153734 73717
rect 153746 73337 154126 73717
rect 154138 73337 154518 73717
rect 154530 73337 154910 73717
rect 154922 73337 155302 73717
rect 155314 73337 155694 73717
rect 155706 73337 156086 73717
rect 153354 72945 153734 73325
rect 153746 72945 154126 73325
rect 154138 72945 154518 73325
rect 154530 72945 154910 73325
rect 154922 72945 155302 73325
rect 155314 72945 155694 73325
rect 155706 72945 156086 73325
rect 153354 72553 153734 72933
rect 153746 72553 154126 72933
rect 154138 72553 154518 72933
rect 154530 72553 154910 72933
rect 154922 72553 155302 72933
rect 155314 72553 155694 72933
rect 155706 72553 156086 72933
rect 153354 72161 153734 72541
rect 153746 72161 154126 72541
rect 154138 72161 154518 72541
rect 154530 72161 154910 72541
rect 154922 72161 155302 72541
rect 155314 72161 155694 72541
rect 155706 72161 156086 72541
rect 139898 70186 140278 70566
rect 139898 69794 140278 70174
rect 139898 69402 140278 69782
rect 139898 69010 140278 69390
rect 139898 68618 140278 68998
rect 139898 68226 140278 68606
rect 139898 67834 140278 68214
rect 160442 74121 160822 74501
rect 160834 74121 161214 74501
rect 161226 74121 161606 74501
rect 161618 74121 161998 74501
rect 162010 74121 162390 74501
rect 162402 74121 162782 74501
rect 162794 74121 163174 74501
rect 163186 74121 163566 74501
rect 163578 74121 163958 74501
rect 160442 73729 160822 74109
rect 160834 73729 161214 74109
rect 161226 73729 161606 74109
rect 161618 73729 161998 74109
rect 162010 73729 162390 74109
rect 162402 73729 162782 74109
rect 162794 73729 163174 74109
rect 163186 73729 163566 74109
rect 163578 73729 163958 74109
rect 160442 73337 160822 73717
rect 160834 73337 161214 73717
rect 161226 73337 161606 73717
rect 161618 73337 161998 73717
rect 162010 73337 162390 73717
rect 162402 73337 162782 73717
rect 162794 73337 163174 73717
rect 163186 73337 163566 73717
rect 163578 73337 163958 73717
rect 160442 72945 160822 73325
rect 160834 72945 161214 73325
rect 161226 72945 161606 73325
rect 161618 72945 161998 73325
rect 162010 72945 162390 73325
rect 162402 72945 162782 73325
rect 162794 72945 163174 73325
rect 163186 72945 163566 73325
rect 163578 72945 163958 73325
rect 160442 72553 160822 72933
rect 160834 72553 161214 72933
rect 161226 72553 161606 72933
rect 161618 72553 161998 72933
rect 162010 72553 162390 72933
rect 162402 72553 162782 72933
rect 162794 72553 163174 72933
rect 163186 72553 163566 72933
rect 163578 72553 163958 72933
rect 160442 72161 160822 72541
rect 160834 72161 161214 72541
rect 161226 72161 161606 72541
rect 161618 72161 161998 72541
rect 162010 72161 162390 72541
rect 162402 72161 162782 72541
rect 162794 72161 163174 72541
rect 163186 72161 163566 72541
rect 163578 72161 163958 72541
rect 153354 70186 153734 70566
rect 153746 70186 154126 70566
rect 154138 70186 154518 70566
rect 154530 70186 154910 70566
rect 154922 70186 155302 70566
rect 155314 70186 155694 70566
rect 155706 70186 156086 70566
rect 153354 69794 153734 70174
rect 153746 69794 154126 70174
rect 154138 69794 154518 70174
rect 154530 69794 154910 70174
rect 154922 69794 155302 70174
rect 155314 69794 155694 70174
rect 155706 69794 156086 70174
rect 153354 69402 153734 69782
rect 153746 69402 154126 69782
rect 154138 69402 154518 69782
rect 154530 69402 154910 69782
rect 154922 69402 155302 69782
rect 155314 69402 155694 69782
rect 155706 69402 156086 69782
rect 153354 69010 153734 69390
rect 153746 69010 154126 69390
rect 154138 69010 154518 69390
rect 154530 69010 154910 69390
rect 154922 69010 155302 69390
rect 155314 69010 155694 69390
rect 155706 69010 156086 69390
rect 153354 68618 153734 68998
rect 153746 68618 154126 68998
rect 154138 68618 154518 68998
rect 154530 68618 154910 68998
rect 154922 68618 155302 68998
rect 155314 68618 155694 68998
rect 155706 68618 156086 68998
rect 153354 68226 153734 68606
rect 153746 68226 154126 68606
rect 154138 68226 154518 68606
rect 154530 68226 154910 68606
rect 154922 68226 155302 68606
rect 155314 68226 155694 68606
rect 155706 68226 156086 68606
rect 153354 67834 153734 68214
rect 153746 67834 154126 68214
rect 154138 67834 154518 68214
rect 154530 67834 154910 68214
rect 154922 67834 155302 68214
rect 155314 67834 155694 68214
rect 155706 67834 156086 68214
<< metal7 >>
rect 65000 196000 79000 210000
rect 81000 196000 95000 210000
rect 97000 196000 111000 210000
rect 113000 196000 127000 210000
rect 129000 196000 143000 210000
rect 145000 196000 159000 210000
rect 14000 145000 28000 159000
rect 67748 155942 156220 156076
rect 67748 155562 67882 155942
rect 68262 155562 68274 155942
rect 68654 155562 68666 155942
rect 69046 155562 69058 155942
rect 69438 155562 69450 155942
rect 69830 155562 69842 155942
rect 70222 155562 70234 155942
rect 70614 155562 79418 155942
rect 79798 155562 94538 155942
rect 94918 155562 109658 155942
rect 110038 155562 124778 155942
rect 125158 155562 139898 155942
rect 140278 155562 153354 155942
rect 153734 155562 153746 155942
rect 154126 155562 154138 155942
rect 154518 155562 154530 155942
rect 154910 155562 154922 155942
rect 155302 155562 155314 155942
rect 155694 155562 155706 155942
rect 156086 155562 156220 155942
rect 67748 155550 156220 155562
rect 67748 155170 67882 155550
rect 68262 155170 68274 155550
rect 68654 155170 68666 155550
rect 69046 155170 69058 155550
rect 69438 155170 69450 155550
rect 69830 155170 69842 155550
rect 70222 155170 70234 155550
rect 70614 155170 79418 155550
rect 79798 155170 94538 155550
rect 94918 155170 109658 155550
rect 110038 155170 124778 155550
rect 125158 155170 139898 155550
rect 140278 155170 153354 155550
rect 153734 155170 153746 155550
rect 154126 155170 154138 155550
rect 154518 155170 154530 155550
rect 154910 155170 154922 155550
rect 155302 155170 155314 155550
rect 155694 155170 155706 155550
rect 156086 155170 156220 155550
rect 67748 155158 156220 155170
rect 67748 154778 67882 155158
rect 68262 154778 68274 155158
rect 68654 154778 68666 155158
rect 69046 154778 69058 155158
rect 69438 154778 69450 155158
rect 69830 154778 69842 155158
rect 70222 154778 70234 155158
rect 70614 154778 79418 155158
rect 79798 154778 94538 155158
rect 94918 154778 109658 155158
rect 110038 154778 124778 155158
rect 125158 154778 139898 155158
rect 140278 154778 153354 155158
rect 153734 154778 153746 155158
rect 154126 154778 154138 155158
rect 154518 154778 154530 155158
rect 154910 154778 154922 155158
rect 155302 154778 155314 155158
rect 155694 154778 155706 155158
rect 156086 154778 156220 155158
rect 67748 154766 156220 154778
rect 67748 154386 67882 154766
rect 68262 154386 68274 154766
rect 68654 154386 68666 154766
rect 69046 154386 69058 154766
rect 69438 154386 69450 154766
rect 69830 154386 69842 154766
rect 70222 154386 70234 154766
rect 70614 154386 79418 154766
rect 79798 154386 94538 154766
rect 94918 154386 109658 154766
rect 110038 154386 124778 154766
rect 125158 154386 139898 154766
rect 140278 154386 153354 154766
rect 153734 154386 153746 154766
rect 154126 154386 154138 154766
rect 154518 154386 154530 154766
rect 154910 154386 154922 154766
rect 155302 154386 155314 154766
rect 155694 154386 155706 154766
rect 156086 154386 156220 154766
rect 67748 154374 156220 154386
rect 67748 153994 67882 154374
rect 68262 153994 68274 154374
rect 68654 153994 68666 154374
rect 69046 153994 69058 154374
rect 69438 153994 69450 154374
rect 69830 153994 69842 154374
rect 70222 153994 70234 154374
rect 70614 153994 79418 154374
rect 79798 153994 94538 154374
rect 94918 153994 109658 154374
rect 110038 153994 124778 154374
rect 125158 153994 139898 154374
rect 140278 153994 153354 154374
rect 153734 153994 153746 154374
rect 154126 153994 154138 154374
rect 154518 153994 154530 154374
rect 154910 153994 154922 154374
rect 155302 153994 155314 154374
rect 155694 153994 155706 154374
rect 156086 153994 156220 154374
rect 67748 153982 156220 153994
rect 67748 153602 67882 153982
rect 68262 153602 68274 153982
rect 68654 153602 68666 153982
rect 69046 153602 69058 153982
rect 69438 153602 69450 153982
rect 69830 153602 69842 153982
rect 70222 153602 70234 153982
rect 70614 153602 79418 153982
rect 79798 153602 94538 153982
rect 94918 153602 109658 153982
rect 110038 153602 124778 153982
rect 125158 153602 139898 153982
rect 140278 153602 153354 153982
rect 153734 153602 153746 153982
rect 154126 153602 154138 153982
rect 154518 153602 154530 153982
rect 154910 153602 154922 153982
rect 155302 153602 155314 153982
rect 155694 153602 155706 153982
rect 156086 153602 156220 153982
rect 67748 153590 156220 153602
rect 67748 153210 67882 153590
rect 68262 153210 68274 153590
rect 68654 153210 68666 153590
rect 69046 153210 69058 153590
rect 69438 153210 69450 153590
rect 69830 153210 69842 153590
rect 70222 153210 70234 153590
rect 70614 153210 79418 153590
rect 79798 153210 94538 153590
rect 94918 153210 109658 153590
rect 110038 153210 124778 153590
rect 125158 153210 139898 153590
rect 140278 153210 153354 153590
rect 153734 153210 153746 153590
rect 154126 153210 154138 153590
rect 154518 153210 154530 153590
rect 154910 153210 154922 153590
rect 155302 153210 155314 153590
rect 155694 153210 155706 153590
rect 156086 153210 156220 153590
rect 67748 153076 156220 153210
rect 71748 151942 152220 152076
rect 71748 151562 71882 151942
rect 72262 151562 72274 151942
rect 72654 151562 72666 151942
rect 73046 151562 73058 151942
rect 73438 151562 73450 151942
rect 73830 151562 73842 151942
rect 74222 151562 74234 151942
rect 74614 151562 78178 151942
rect 78558 151562 93298 151942
rect 93678 151562 108418 151942
rect 108798 151562 123538 151942
rect 123918 151562 138658 151942
rect 139038 151562 149354 151942
rect 149734 151562 149746 151942
rect 150126 151562 150138 151942
rect 150518 151562 150530 151942
rect 150910 151562 150922 151942
rect 151302 151562 151314 151942
rect 151694 151562 151706 151942
rect 152086 151562 152220 151942
rect 71748 151550 152220 151562
rect 71748 151170 71882 151550
rect 72262 151170 72274 151550
rect 72654 151170 72666 151550
rect 73046 151170 73058 151550
rect 73438 151170 73450 151550
rect 73830 151170 73842 151550
rect 74222 151170 74234 151550
rect 74614 151170 78178 151550
rect 78558 151170 93298 151550
rect 93678 151170 108418 151550
rect 108798 151170 123538 151550
rect 123918 151170 138658 151550
rect 139038 151170 149354 151550
rect 149734 151170 149746 151550
rect 150126 151170 150138 151550
rect 150518 151170 150530 151550
rect 150910 151170 150922 151550
rect 151302 151170 151314 151550
rect 151694 151170 151706 151550
rect 152086 151170 152220 151550
rect 71748 151158 152220 151170
rect 71748 150778 71882 151158
rect 72262 150778 72274 151158
rect 72654 150778 72666 151158
rect 73046 150778 73058 151158
rect 73438 150778 73450 151158
rect 73830 150778 73842 151158
rect 74222 150778 74234 151158
rect 74614 150778 78178 151158
rect 78558 150778 93298 151158
rect 93678 150778 108418 151158
rect 108798 150778 123538 151158
rect 123918 150778 138658 151158
rect 139038 150778 149354 151158
rect 149734 150778 149746 151158
rect 150126 150778 150138 151158
rect 150518 150778 150530 151158
rect 150910 150778 150922 151158
rect 151302 150778 151314 151158
rect 151694 150778 151706 151158
rect 152086 150778 152220 151158
rect 71748 150766 152220 150778
rect 71748 150386 71882 150766
rect 72262 150386 72274 150766
rect 72654 150386 72666 150766
rect 73046 150386 73058 150766
rect 73438 150386 73450 150766
rect 73830 150386 73842 150766
rect 74222 150386 74234 150766
rect 74614 150386 78178 150766
rect 78558 150386 93298 150766
rect 93678 150386 108418 150766
rect 108798 150386 123538 150766
rect 123918 150386 138658 150766
rect 139038 150386 149354 150766
rect 149734 150386 149746 150766
rect 150126 150386 150138 150766
rect 150518 150386 150530 150766
rect 150910 150386 150922 150766
rect 151302 150386 151314 150766
rect 151694 150386 151706 150766
rect 152086 150386 152220 150766
rect 71748 150374 152220 150386
rect 71748 149994 71882 150374
rect 72262 149994 72274 150374
rect 72654 149994 72666 150374
rect 73046 149994 73058 150374
rect 73438 149994 73450 150374
rect 73830 149994 73842 150374
rect 74222 149994 74234 150374
rect 74614 149994 78178 150374
rect 78558 149994 93298 150374
rect 93678 149994 108418 150374
rect 108798 149994 123538 150374
rect 123918 149994 138658 150374
rect 139038 149994 149354 150374
rect 149734 149994 149746 150374
rect 150126 149994 150138 150374
rect 150518 149994 150530 150374
rect 150910 149994 150922 150374
rect 151302 149994 151314 150374
rect 151694 149994 151706 150374
rect 152086 149994 152220 150374
rect 71748 149982 152220 149994
rect 71748 149602 71882 149982
rect 72262 149602 72274 149982
rect 72654 149602 72666 149982
rect 73046 149602 73058 149982
rect 73438 149602 73450 149982
rect 73830 149602 73842 149982
rect 74222 149602 74234 149982
rect 74614 149602 78178 149982
rect 78558 149602 93298 149982
rect 93678 149602 108418 149982
rect 108798 149602 123538 149982
rect 123918 149602 138658 149982
rect 139038 149602 149354 149982
rect 149734 149602 149746 149982
rect 150126 149602 150138 149982
rect 150518 149602 150530 149982
rect 150910 149602 150922 149982
rect 151302 149602 151314 149982
rect 151694 149602 151706 149982
rect 152086 149602 152220 149982
rect 71748 149590 152220 149602
rect 71748 149210 71882 149590
rect 72262 149210 72274 149590
rect 72654 149210 72666 149590
rect 73046 149210 73058 149590
rect 73438 149210 73450 149590
rect 73830 149210 73842 149590
rect 74222 149210 74234 149590
rect 74614 149210 78178 149590
rect 78558 149210 93298 149590
rect 93678 149210 108418 149590
rect 108798 149210 123538 149590
rect 123918 149210 138658 149590
rect 139038 149210 149354 149590
rect 149734 149210 149746 149590
rect 150126 149210 150138 149590
rect 150518 149210 150530 149590
rect 150910 149210 150922 149590
rect 151302 149210 151314 149590
rect 151694 149210 151706 149590
rect 152086 149210 152220 149590
rect 71748 149076 152220 149210
rect 196000 145000 210000 159000
rect 14000 129000 28000 143000
rect 67748 140230 156220 140260
rect 67748 139850 67882 140230
rect 68262 139850 68274 140230
rect 68654 139850 68666 140230
rect 69046 139850 69058 140230
rect 69438 139850 69450 140230
rect 69830 139850 69842 140230
rect 70222 139850 70234 140230
rect 70614 139850 79418 140230
rect 79798 139850 94538 140230
rect 94918 139850 109658 140230
rect 110038 139850 124778 140230
rect 125158 139850 139898 140230
rect 140278 139850 153354 140230
rect 153734 139850 153746 140230
rect 154126 139850 154138 140230
rect 154518 139850 154530 140230
rect 154910 139850 154922 140230
rect 155302 139850 155314 140230
rect 155694 139850 155706 140230
rect 156086 139850 156220 140230
rect 67748 139820 156220 139850
rect 71748 138990 152220 139020
rect 71748 138610 71882 138990
rect 72262 138610 72274 138990
rect 72654 138610 72666 138990
rect 73046 138610 73058 138990
rect 73438 138610 73450 138990
rect 73830 138610 73842 138990
rect 74222 138610 74234 138990
rect 74614 138610 78178 138990
rect 78558 138610 93298 138990
rect 93678 138610 108418 138990
rect 108798 138610 123538 138990
rect 123918 138610 138658 138990
rect 139038 138610 149354 138990
rect 149734 138610 149746 138990
rect 150126 138610 150138 138990
rect 150518 138610 150530 138990
rect 150910 138610 150922 138990
rect 151302 138610 151314 138990
rect 151694 138610 151706 138990
rect 152086 138610 152220 138990
rect 71748 138580 152220 138610
rect 56000 133169 74748 133332
rect 56000 132789 56042 133169
rect 56422 132789 56434 133169
rect 56814 132789 56826 133169
rect 57206 132789 57218 133169
rect 57598 132789 57610 133169
rect 57990 132789 58002 133169
rect 58382 132789 58394 133169
rect 58774 132789 58786 133169
rect 59166 132789 59178 133169
rect 59558 132789 71882 133169
rect 72262 132789 72274 133169
rect 72654 132789 72666 133169
rect 73046 132789 73058 133169
rect 73438 132789 73450 133169
rect 73830 132789 73842 133169
rect 74222 132789 74234 133169
rect 74614 132789 74748 133169
rect 56000 132777 74748 132789
rect 56000 132397 56042 132777
rect 56422 132397 56434 132777
rect 56814 132397 56826 132777
rect 57206 132397 57218 132777
rect 57598 132397 57610 132777
rect 57990 132397 58002 132777
rect 58382 132397 58394 132777
rect 58774 132397 58786 132777
rect 59166 132397 59178 132777
rect 59558 132397 71882 132777
rect 72262 132397 72274 132777
rect 72654 132397 72666 132777
rect 73046 132397 73058 132777
rect 73438 132397 73450 132777
rect 73830 132397 73842 132777
rect 74222 132397 74234 132777
rect 74614 132397 74748 132777
rect 56000 132385 74748 132397
rect 56000 132005 56042 132385
rect 56422 132005 56434 132385
rect 56814 132005 56826 132385
rect 57206 132005 57218 132385
rect 57598 132005 57610 132385
rect 57990 132005 58002 132385
rect 58382 132005 58394 132385
rect 58774 132005 58786 132385
rect 59166 132005 59178 132385
rect 59558 132005 71882 132385
rect 72262 132005 72274 132385
rect 72654 132005 72666 132385
rect 73046 132005 73058 132385
rect 73438 132005 73450 132385
rect 73830 132005 73842 132385
rect 74222 132005 74234 132385
rect 74614 132005 74748 132385
rect 56000 131993 74748 132005
rect 56000 131613 56042 131993
rect 56422 131613 56434 131993
rect 56814 131613 56826 131993
rect 57206 131613 57218 131993
rect 57598 131613 57610 131993
rect 57990 131613 58002 131993
rect 58382 131613 58394 131993
rect 58774 131613 58786 131993
rect 59166 131613 59178 131993
rect 59558 131613 71882 131993
rect 72262 131613 72274 131993
rect 72654 131613 72666 131993
rect 73046 131613 73058 131993
rect 73438 131613 73450 131993
rect 73830 131613 73842 131993
rect 74222 131613 74234 131993
rect 74614 131613 74748 131993
rect 56000 131601 74748 131613
rect 56000 131221 56042 131601
rect 56422 131221 56434 131601
rect 56814 131221 56826 131601
rect 57206 131221 57218 131601
rect 57598 131221 57610 131601
rect 57990 131221 58002 131601
rect 58382 131221 58394 131601
rect 58774 131221 58786 131601
rect 59166 131221 59178 131601
rect 59558 131221 71882 131601
rect 72262 131221 72274 131601
rect 72654 131221 72666 131601
rect 73046 131221 73058 131601
rect 73438 131221 73450 131601
rect 73830 131221 73842 131601
rect 74222 131221 74234 131601
rect 74614 131221 74748 131601
rect 56000 131209 74748 131221
rect 56000 130829 56042 131209
rect 56422 130829 56434 131209
rect 56814 130829 56826 131209
rect 57206 130829 57218 131209
rect 57598 130829 57610 131209
rect 57990 130829 58002 131209
rect 58382 130829 58394 131209
rect 58774 130829 58786 131209
rect 59166 130829 59178 131209
rect 59558 130829 71882 131209
rect 72262 130829 72274 131209
rect 72654 130829 72666 131209
rect 73046 130829 73058 131209
rect 73438 130829 73450 131209
rect 73830 130829 73842 131209
rect 74222 130829 74234 131209
rect 74614 130829 74748 131209
rect 56000 130666 74748 130829
rect 149220 133169 168000 133332
rect 149220 132789 149354 133169
rect 149734 132789 149746 133169
rect 150126 132789 150138 133169
rect 150518 132789 150530 133169
rect 150910 132789 150922 133169
rect 151302 132789 151314 133169
rect 151694 132789 151706 133169
rect 152086 132789 164442 133169
rect 164822 132789 164834 133169
rect 165214 132789 165226 133169
rect 165606 132789 165618 133169
rect 165998 132789 166010 133169
rect 166390 132789 166402 133169
rect 166782 132789 166794 133169
rect 167174 132789 167186 133169
rect 167566 132789 167578 133169
rect 167958 132789 168000 133169
rect 149220 132777 168000 132789
rect 149220 132397 149354 132777
rect 149734 132397 149746 132777
rect 150126 132397 150138 132777
rect 150518 132397 150530 132777
rect 150910 132397 150922 132777
rect 151302 132397 151314 132777
rect 151694 132397 151706 132777
rect 152086 132397 164442 132777
rect 164822 132397 164834 132777
rect 165214 132397 165226 132777
rect 165606 132397 165618 132777
rect 165998 132397 166010 132777
rect 166390 132397 166402 132777
rect 166782 132397 166794 132777
rect 167174 132397 167186 132777
rect 167566 132397 167578 132777
rect 167958 132397 168000 132777
rect 149220 132385 168000 132397
rect 149220 132005 149354 132385
rect 149734 132005 149746 132385
rect 150126 132005 150138 132385
rect 150518 132005 150530 132385
rect 150910 132005 150922 132385
rect 151302 132005 151314 132385
rect 151694 132005 151706 132385
rect 152086 132005 164442 132385
rect 164822 132005 164834 132385
rect 165214 132005 165226 132385
rect 165606 132005 165618 132385
rect 165998 132005 166010 132385
rect 166390 132005 166402 132385
rect 166782 132005 166794 132385
rect 167174 132005 167186 132385
rect 167566 132005 167578 132385
rect 167958 132005 168000 132385
rect 149220 131993 168000 132005
rect 149220 131613 149354 131993
rect 149734 131613 149746 131993
rect 150126 131613 150138 131993
rect 150518 131613 150530 131993
rect 150910 131613 150922 131993
rect 151302 131613 151314 131993
rect 151694 131613 151706 131993
rect 152086 131613 164442 131993
rect 164822 131613 164834 131993
rect 165214 131613 165226 131993
rect 165606 131613 165618 131993
rect 165998 131613 166010 131993
rect 166390 131613 166402 131993
rect 166782 131613 166794 131993
rect 167174 131613 167186 131993
rect 167566 131613 167578 131993
rect 167958 131613 168000 131993
rect 149220 131601 168000 131613
rect 149220 131221 149354 131601
rect 149734 131221 149746 131601
rect 150126 131221 150138 131601
rect 150518 131221 150530 131601
rect 150910 131221 150922 131601
rect 151302 131221 151314 131601
rect 151694 131221 151706 131601
rect 152086 131221 164442 131601
rect 164822 131221 164834 131601
rect 165214 131221 165226 131601
rect 165606 131221 165618 131601
rect 165998 131221 166010 131601
rect 166390 131221 166402 131601
rect 166782 131221 166794 131601
rect 167174 131221 167186 131601
rect 167566 131221 167578 131601
rect 167958 131221 168000 131601
rect 149220 131209 168000 131221
rect 149220 130829 149354 131209
rect 149734 130829 149746 131209
rect 150126 130829 150138 131209
rect 150518 130829 150530 131209
rect 150910 130829 150922 131209
rect 151302 130829 151314 131209
rect 151694 130829 151706 131209
rect 152086 130829 164442 131209
rect 164822 130829 164834 131209
rect 165214 130829 165226 131209
rect 165606 130829 165618 131209
rect 165998 130829 166010 131209
rect 166390 130829 166402 131209
rect 166782 130829 166794 131209
rect 167174 130829 167186 131209
rect 167566 130829 167578 131209
rect 167958 130829 168000 131209
rect 149220 130666 168000 130829
rect 196000 129000 210000 143000
rect 14000 113000 28000 127000
rect 67748 125110 156220 125140
rect 67748 124730 67882 125110
rect 68262 124730 68274 125110
rect 68654 124730 68666 125110
rect 69046 124730 69058 125110
rect 69438 124730 69450 125110
rect 69830 124730 69842 125110
rect 70222 124730 70234 125110
rect 70614 124730 79418 125110
rect 79798 124730 94538 125110
rect 94918 124730 109658 125110
rect 110038 124730 124778 125110
rect 125158 124730 139898 125110
rect 140278 124730 153354 125110
rect 153734 124730 153746 125110
rect 154126 124730 154138 125110
rect 154518 124730 154530 125110
rect 154910 124730 154922 125110
rect 155302 124730 155314 125110
rect 155694 124730 155706 125110
rect 156086 124730 156220 125110
rect 67748 124700 156220 124730
rect 71748 123870 152220 123900
rect 71748 123490 71882 123870
rect 72262 123490 72274 123870
rect 72654 123490 72666 123870
rect 73046 123490 73058 123870
rect 73438 123490 73450 123870
rect 73830 123490 73842 123870
rect 74222 123490 74234 123870
rect 74614 123490 78178 123870
rect 78558 123490 93298 123870
rect 93678 123490 108418 123870
rect 108798 123490 123538 123870
rect 123918 123490 138658 123870
rect 139038 123490 149354 123870
rect 149734 123490 149746 123870
rect 150126 123490 150138 123870
rect 150518 123490 150530 123870
rect 150910 123490 150922 123870
rect 151302 123490 151314 123870
rect 151694 123490 151706 123870
rect 152086 123490 152220 123870
rect 71748 123460 152220 123490
rect 56000 117169 74748 117332
rect 56000 116789 56042 117169
rect 56422 116789 56434 117169
rect 56814 116789 56826 117169
rect 57206 116789 57218 117169
rect 57598 116789 57610 117169
rect 57990 116789 58002 117169
rect 58382 116789 58394 117169
rect 58774 116789 58786 117169
rect 59166 116789 59178 117169
rect 59558 116789 71882 117169
rect 72262 116789 72274 117169
rect 72654 116789 72666 117169
rect 73046 116789 73058 117169
rect 73438 116789 73450 117169
rect 73830 116789 73842 117169
rect 74222 116789 74234 117169
rect 74614 116789 74748 117169
rect 56000 116777 74748 116789
rect 56000 116397 56042 116777
rect 56422 116397 56434 116777
rect 56814 116397 56826 116777
rect 57206 116397 57218 116777
rect 57598 116397 57610 116777
rect 57990 116397 58002 116777
rect 58382 116397 58394 116777
rect 58774 116397 58786 116777
rect 59166 116397 59178 116777
rect 59558 116397 71882 116777
rect 72262 116397 72274 116777
rect 72654 116397 72666 116777
rect 73046 116397 73058 116777
rect 73438 116397 73450 116777
rect 73830 116397 73842 116777
rect 74222 116397 74234 116777
rect 74614 116397 74748 116777
rect 56000 116385 74748 116397
rect 56000 116005 56042 116385
rect 56422 116005 56434 116385
rect 56814 116005 56826 116385
rect 57206 116005 57218 116385
rect 57598 116005 57610 116385
rect 57990 116005 58002 116385
rect 58382 116005 58394 116385
rect 58774 116005 58786 116385
rect 59166 116005 59178 116385
rect 59558 116005 71882 116385
rect 72262 116005 72274 116385
rect 72654 116005 72666 116385
rect 73046 116005 73058 116385
rect 73438 116005 73450 116385
rect 73830 116005 73842 116385
rect 74222 116005 74234 116385
rect 74614 116005 74748 116385
rect 56000 115993 74748 116005
rect 56000 115613 56042 115993
rect 56422 115613 56434 115993
rect 56814 115613 56826 115993
rect 57206 115613 57218 115993
rect 57598 115613 57610 115993
rect 57990 115613 58002 115993
rect 58382 115613 58394 115993
rect 58774 115613 58786 115993
rect 59166 115613 59178 115993
rect 59558 115613 71882 115993
rect 72262 115613 72274 115993
rect 72654 115613 72666 115993
rect 73046 115613 73058 115993
rect 73438 115613 73450 115993
rect 73830 115613 73842 115993
rect 74222 115613 74234 115993
rect 74614 115613 74748 115993
rect 56000 115601 74748 115613
rect 56000 115221 56042 115601
rect 56422 115221 56434 115601
rect 56814 115221 56826 115601
rect 57206 115221 57218 115601
rect 57598 115221 57610 115601
rect 57990 115221 58002 115601
rect 58382 115221 58394 115601
rect 58774 115221 58786 115601
rect 59166 115221 59178 115601
rect 59558 115221 71882 115601
rect 72262 115221 72274 115601
rect 72654 115221 72666 115601
rect 73046 115221 73058 115601
rect 73438 115221 73450 115601
rect 73830 115221 73842 115601
rect 74222 115221 74234 115601
rect 74614 115221 74748 115601
rect 56000 115209 74748 115221
rect 56000 114829 56042 115209
rect 56422 114829 56434 115209
rect 56814 114829 56826 115209
rect 57206 114829 57218 115209
rect 57598 114829 57610 115209
rect 57990 114829 58002 115209
rect 58382 114829 58394 115209
rect 58774 114829 58786 115209
rect 59166 114829 59178 115209
rect 59558 114829 71882 115209
rect 72262 114829 72274 115209
rect 72654 114829 72666 115209
rect 73046 114829 73058 115209
rect 73438 114829 73450 115209
rect 73830 114829 73842 115209
rect 74222 114829 74234 115209
rect 74614 114829 74748 115209
rect 56000 114666 74748 114829
rect 149220 117169 168000 117332
rect 149220 116789 149354 117169
rect 149734 116789 149746 117169
rect 150126 116789 150138 117169
rect 150518 116789 150530 117169
rect 150910 116789 150922 117169
rect 151302 116789 151314 117169
rect 151694 116789 151706 117169
rect 152086 116789 164442 117169
rect 164822 116789 164834 117169
rect 165214 116789 165226 117169
rect 165606 116789 165618 117169
rect 165998 116789 166010 117169
rect 166390 116789 166402 117169
rect 166782 116789 166794 117169
rect 167174 116789 167186 117169
rect 167566 116789 167578 117169
rect 167958 116789 168000 117169
rect 149220 116777 168000 116789
rect 149220 116397 149354 116777
rect 149734 116397 149746 116777
rect 150126 116397 150138 116777
rect 150518 116397 150530 116777
rect 150910 116397 150922 116777
rect 151302 116397 151314 116777
rect 151694 116397 151706 116777
rect 152086 116397 164442 116777
rect 164822 116397 164834 116777
rect 165214 116397 165226 116777
rect 165606 116397 165618 116777
rect 165998 116397 166010 116777
rect 166390 116397 166402 116777
rect 166782 116397 166794 116777
rect 167174 116397 167186 116777
rect 167566 116397 167578 116777
rect 167958 116397 168000 116777
rect 149220 116385 168000 116397
rect 149220 116005 149354 116385
rect 149734 116005 149746 116385
rect 150126 116005 150138 116385
rect 150518 116005 150530 116385
rect 150910 116005 150922 116385
rect 151302 116005 151314 116385
rect 151694 116005 151706 116385
rect 152086 116005 164442 116385
rect 164822 116005 164834 116385
rect 165214 116005 165226 116385
rect 165606 116005 165618 116385
rect 165998 116005 166010 116385
rect 166390 116005 166402 116385
rect 166782 116005 166794 116385
rect 167174 116005 167186 116385
rect 167566 116005 167578 116385
rect 167958 116005 168000 116385
rect 149220 115993 168000 116005
rect 149220 115613 149354 115993
rect 149734 115613 149746 115993
rect 150126 115613 150138 115993
rect 150518 115613 150530 115993
rect 150910 115613 150922 115993
rect 151302 115613 151314 115993
rect 151694 115613 151706 115993
rect 152086 115613 164442 115993
rect 164822 115613 164834 115993
rect 165214 115613 165226 115993
rect 165606 115613 165618 115993
rect 165998 115613 166010 115993
rect 166390 115613 166402 115993
rect 166782 115613 166794 115993
rect 167174 115613 167186 115993
rect 167566 115613 167578 115993
rect 167958 115613 168000 115993
rect 149220 115601 168000 115613
rect 149220 115221 149354 115601
rect 149734 115221 149746 115601
rect 150126 115221 150138 115601
rect 150518 115221 150530 115601
rect 150910 115221 150922 115601
rect 151302 115221 151314 115601
rect 151694 115221 151706 115601
rect 152086 115221 164442 115601
rect 164822 115221 164834 115601
rect 165214 115221 165226 115601
rect 165606 115221 165618 115601
rect 165998 115221 166010 115601
rect 166390 115221 166402 115601
rect 166782 115221 166794 115601
rect 167174 115221 167186 115601
rect 167566 115221 167578 115601
rect 167958 115221 168000 115601
rect 149220 115209 168000 115221
rect 149220 114829 149354 115209
rect 149734 114829 149746 115209
rect 150126 114829 150138 115209
rect 150518 114829 150530 115209
rect 150910 114829 150922 115209
rect 151302 114829 151314 115209
rect 151694 114829 151706 115209
rect 152086 114829 164442 115209
rect 164822 114829 164834 115209
rect 165214 114829 165226 115209
rect 165606 114829 165618 115209
rect 165998 114829 166010 115209
rect 166390 114829 166402 115209
rect 166782 114829 166794 115209
rect 167174 114829 167186 115209
rect 167566 114829 167578 115209
rect 167958 114829 168000 115209
rect 149220 114666 168000 114829
rect 196000 113000 210000 127000
rect 14000 97000 28000 111000
rect 67748 109990 156220 110020
rect 67748 109610 67882 109990
rect 68262 109610 68274 109990
rect 68654 109610 68666 109990
rect 69046 109610 69058 109990
rect 69438 109610 69450 109990
rect 69830 109610 69842 109990
rect 70222 109610 70234 109990
rect 70614 109610 79418 109990
rect 79798 109610 94538 109990
rect 94918 109610 109658 109990
rect 110038 109610 124778 109990
rect 125158 109610 139898 109990
rect 140278 109610 153354 109990
rect 153734 109610 153746 109990
rect 154126 109610 154138 109990
rect 154518 109610 154530 109990
rect 154910 109610 154922 109990
rect 155302 109610 155314 109990
rect 155694 109610 155706 109990
rect 156086 109610 156220 109990
rect 67748 109580 156220 109610
rect 71748 108750 152220 108780
rect 71748 108370 71882 108750
rect 72262 108370 72274 108750
rect 72654 108370 72666 108750
rect 73046 108370 73058 108750
rect 73438 108370 73450 108750
rect 73830 108370 73842 108750
rect 74222 108370 74234 108750
rect 74614 108370 78178 108750
rect 78558 108370 93298 108750
rect 93678 108370 108418 108750
rect 108798 108370 123538 108750
rect 123918 108370 138658 108750
rect 139038 108370 149354 108750
rect 149734 108370 149746 108750
rect 150126 108370 150138 108750
rect 150518 108370 150530 108750
rect 150910 108370 150922 108750
rect 151302 108370 151314 108750
rect 151694 108370 151706 108750
rect 152086 108370 152220 108750
rect 71748 108340 152220 108370
rect 60000 106501 70748 106664
rect 60000 106121 60042 106501
rect 60422 106121 60434 106501
rect 60814 106121 60826 106501
rect 61206 106121 61218 106501
rect 61598 106121 61610 106501
rect 61990 106121 62002 106501
rect 62382 106121 62394 106501
rect 62774 106121 62786 106501
rect 63166 106121 63178 106501
rect 63558 106121 67882 106501
rect 68262 106121 68274 106501
rect 68654 106121 68666 106501
rect 69046 106121 69058 106501
rect 69438 106121 69450 106501
rect 69830 106121 69842 106501
rect 70222 106121 70234 106501
rect 70614 106121 70748 106501
rect 60000 106109 70748 106121
rect 60000 105729 60042 106109
rect 60422 105729 60434 106109
rect 60814 105729 60826 106109
rect 61206 105729 61218 106109
rect 61598 105729 61610 106109
rect 61990 105729 62002 106109
rect 62382 105729 62394 106109
rect 62774 105729 62786 106109
rect 63166 105729 63178 106109
rect 63558 105729 67882 106109
rect 68262 105729 68274 106109
rect 68654 105729 68666 106109
rect 69046 105729 69058 106109
rect 69438 105729 69450 106109
rect 69830 105729 69842 106109
rect 70222 105729 70234 106109
rect 70614 105729 70748 106109
rect 60000 105717 70748 105729
rect 60000 105337 60042 105717
rect 60422 105337 60434 105717
rect 60814 105337 60826 105717
rect 61206 105337 61218 105717
rect 61598 105337 61610 105717
rect 61990 105337 62002 105717
rect 62382 105337 62394 105717
rect 62774 105337 62786 105717
rect 63166 105337 63178 105717
rect 63558 105337 67882 105717
rect 68262 105337 68274 105717
rect 68654 105337 68666 105717
rect 69046 105337 69058 105717
rect 69438 105337 69450 105717
rect 69830 105337 69842 105717
rect 70222 105337 70234 105717
rect 70614 105337 70748 105717
rect 60000 105325 70748 105337
rect 60000 104945 60042 105325
rect 60422 104945 60434 105325
rect 60814 104945 60826 105325
rect 61206 104945 61218 105325
rect 61598 104945 61610 105325
rect 61990 104945 62002 105325
rect 62382 104945 62394 105325
rect 62774 104945 62786 105325
rect 63166 104945 63178 105325
rect 63558 104945 67882 105325
rect 68262 104945 68274 105325
rect 68654 104945 68666 105325
rect 69046 104945 69058 105325
rect 69438 104945 69450 105325
rect 69830 104945 69842 105325
rect 70222 104945 70234 105325
rect 70614 104945 70748 105325
rect 60000 104933 70748 104945
rect 60000 104553 60042 104933
rect 60422 104553 60434 104933
rect 60814 104553 60826 104933
rect 61206 104553 61218 104933
rect 61598 104553 61610 104933
rect 61990 104553 62002 104933
rect 62382 104553 62394 104933
rect 62774 104553 62786 104933
rect 63166 104553 63178 104933
rect 63558 104553 67882 104933
rect 68262 104553 68274 104933
rect 68654 104553 68666 104933
rect 69046 104553 69058 104933
rect 69438 104553 69450 104933
rect 69830 104553 69842 104933
rect 70222 104553 70234 104933
rect 70614 104553 70748 104933
rect 60000 104541 70748 104553
rect 60000 104161 60042 104541
rect 60422 104161 60434 104541
rect 60814 104161 60826 104541
rect 61206 104161 61218 104541
rect 61598 104161 61610 104541
rect 61990 104161 62002 104541
rect 62382 104161 62394 104541
rect 62774 104161 62786 104541
rect 63166 104161 63178 104541
rect 63558 104161 67882 104541
rect 68262 104161 68274 104541
rect 68654 104161 68666 104541
rect 69046 104161 69058 104541
rect 69438 104161 69450 104541
rect 69830 104161 69842 104541
rect 70222 104161 70234 104541
rect 70614 104161 70748 104541
rect 60000 103998 70748 104161
rect 153220 106501 164000 106664
rect 153220 106121 153354 106501
rect 153734 106121 153746 106501
rect 154126 106121 154138 106501
rect 154518 106121 154530 106501
rect 154910 106121 154922 106501
rect 155302 106121 155314 106501
rect 155694 106121 155706 106501
rect 156086 106121 160442 106501
rect 160822 106121 160834 106501
rect 161214 106121 161226 106501
rect 161606 106121 161618 106501
rect 161998 106121 162010 106501
rect 162390 106121 162402 106501
rect 162782 106121 162794 106501
rect 163174 106121 163186 106501
rect 163566 106121 163578 106501
rect 163958 106121 164000 106501
rect 153220 106109 164000 106121
rect 153220 105729 153354 106109
rect 153734 105729 153746 106109
rect 154126 105729 154138 106109
rect 154518 105729 154530 106109
rect 154910 105729 154922 106109
rect 155302 105729 155314 106109
rect 155694 105729 155706 106109
rect 156086 105729 160442 106109
rect 160822 105729 160834 106109
rect 161214 105729 161226 106109
rect 161606 105729 161618 106109
rect 161998 105729 162010 106109
rect 162390 105729 162402 106109
rect 162782 105729 162794 106109
rect 163174 105729 163186 106109
rect 163566 105729 163578 106109
rect 163958 105729 164000 106109
rect 153220 105717 164000 105729
rect 153220 105337 153354 105717
rect 153734 105337 153746 105717
rect 154126 105337 154138 105717
rect 154518 105337 154530 105717
rect 154910 105337 154922 105717
rect 155302 105337 155314 105717
rect 155694 105337 155706 105717
rect 156086 105337 160442 105717
rect 160822 105337 160834 105717
rect 161214 105337 161226 105717
rect 161606 105337 161618 105717
rect 161998 105337 162010 105717
rect 162390 105337 162402 105717
rect 162782 105337 162794 105717
rect 163174 105337 163186 105717
rect 163566 105337 163578 105717
rect 163958 105337 164000 105717
rect 153220 105325 164000 105337
rect 153220 104945 153354 105325
rect 153734 104945 153746 105325
rect 154126 104945 154138 105325
rect 154518 104945 154530 105325
rect 154910 104945 154922 105325
rect 155302 104945 155314 105325
rect 155694 104945 155706 105325
rect 156086 104945 160442 105325
rect 160822 104945 160834 105325
rect 161214 104945 161226 105325
rect 161606 104945 161618 105325
rect 161998 104945 162010 105325
rect 162390 104945 162402 105325
rect 162782 104945 162794 105325
rect 163174 104945 163186 105325
rect 163566 104945 163578 105325
rect 163958 104945 164000 105325
rect 153220 104933 164000 104945
rect 153220 104553 153354 104933
rect 153734 104553 153746 104933
rect 154126 104553 154138 104933
rect 154518 104553 154530 104933
rect 154910 104553 154922 104933
rect 155302 104553 155314 104933
rect 155694 104553 155706 104933
rect 156086 104553 160442 104933
rect 160822 104553 160834 104933
rect 161214 104553 161226 104933
rect 161606 104553 161618 104933
rect 161998 104553 162010 104933
rect 162390 104553 162402 104933
rect 162782 104553 162794 104933
rect 163174 104553 163186 104933
rect 163566 104553 163578 104933
rect 163958 104553 164000 104933
rect 153220 104541 164000 104553
rect 153220 104161 153354 104541
rect 153734 104161 153746 104541
rect 154126 104161 154138 104541
rect 154518 104161 154530 104541
rect 154910 104161 154922 104541
rect 155302 104161 155314 104541
rect 155694 104161 155706 104541
rect 156086 104161 160442 104541
rect 160822 104161 160834 104541
rect 161214 104161 161226 104541
rect 161606 104161 161618 104541
rect 161998 104161 162010 104541
rect 162390 104161 162402 104541
rect 162782 104161 162794 104541
rect 163174 104161 163186 104541
rect 163566 104161 163578 104541
rect 163958 104161 164000 104541
rect 153220 103998 164000 104161
rect 56000 101169 74748 101332
rect 56000 100789 56042 101169
rect 56422 100789 56434 101169
rect 56814 100789 56826 101169
rect 57206 100789 57218 101169
rect 57598 100789 57610 101169
rect 57990 100789 58002 101169
rect 58382 100789 58394 101169
rect 58774 100789 58786 101169
rect 59166 100789 59178 101169
rect 59558 100789 71882 101169
rect 72262 100789 72274 101169
rect 72654 100789 72666 101169
rect 73046 100789 73058 101169
rect 73438 100789 73450 101169
rect 73830 100789 73842 101169
rect 74222 100789 74234 101169
rect 74614 100789 74748 101169
rect 56000 100777 74748 100789
rect 56000 100397 56042 100777
rect 56422 100397 56434 100777
rect 56814 100397 56826 100777
rect 57206 100397 57218 100777
rect 57598 100397 57610 100777
rect 57990 100397 58002 100777
rect 58382 100397 58394 100777
rect 58774 100397 58786 100777
rect 59166 100397 59178 100777
rect 59558 100397 71882 100777
rect 72262 100397 72274 100777
rect 72654 100397 72666 100777
rect 73046 100397 73058 100777
rect 73438 100397 73450 100777
rect 73830 100397 73842 100777
rect 74222 100397 74234 100777
rect 74614 100397 74748 100777
rect 56000 100385 74748 100397
rect 56000 100005 56042 100385
rect 56422 100005 56434 100385
rect 56814 100005 56826 100385
rect 57206 100005 57218 100385
rect 57598 100005 57610 100385
rect 57990 100005 58002 100385
rect 58382 100005 58394 100385
rect 58774 100005 58786 100385
rect 59166 100005 59178 100385
rect 59558 100005 71882 100385
rect 72262 100005 72274 100385
rect 72654 100005 72666 100385
rect 73046 100005 73058 100385
rect 73438 100005 73450 100385
rect 73830 100005 73842 100385
rect 74222 100005 74234 100385
rect 74614 100005 74748 100385
rect 56000 99993 74748 100005
rect 56000 99613 56042 99993
rect 56422 99613 56434 99993
rect 56814 99613 56826 99993
rect 57206 99613 57218 99993
rect 57598 99613 57610 99993
rect 57990 99613 58002 99993
rect 58382 99613 58394 99993
rect 58774 99613 58786 99993
rect 59166 99613 59178 99993
rect 59558 99613 71882 99993
rect 72262 99613 72274 99993
rect 72654 99613 72666 99993
rect 73046 99613 73058 99993
rect 73438 99613 73450 99993
rect 73830 99613 73842 99993
rect 74222 99613 74234 99993
rect 74614 99613 74748 99993
rect 56000 99601 74748 99613
rect 56000 99221 56042 99601
rect 56422 99221 56434 99601
rect 56814 99221 56826 99601
rect 57206 99221 57218 99601
rect 57598 99221 57610 99601
rect 57990 99221 58002 99601
rect 58382 99221 58394 99601
rect 58774 99221 58786 99601
rect 59166 99221 59178 99601
rect 59558 99221 71882 99601
rect 72262 99221 72274 99601
rect 72654 99221 72666 99601
rect 73046 99221 73058 99601
rect 73438 99221 73450 99601
rect 73830 99221 73842 99601
rect 74222 99221 74234 99601
rect 74614 99221 74748 99601
rect 56000 99209 74748 99221
rect 56000 98829 56042 99209
rect 56422 98829 56434 99209
rect 56814 98829 56826 99209
rect 57206 98829 57218 99209
rect 57598 98829 57610 99209
rect 57990 98829 58002 99209
rect 58382 98829 58394 99209
rect 58774 98829 58786 99209
rect 59166 98829 59178 99209
rect 59558 98829 71882 99209
rect 72262 98829 72274 99209
rect 72654 98829 72666 99209
rect 73046 98829 73058 99209
rect 73438 98829 73450 99209
rect 73830 98829 73842 99209
rect 74222 98829 74234 99209
rect 74614 98829 74748 99209
rect 56000 98666 74748 98829
rect 149220 101169 168000 101332
rect 149220 100789 149354 101169
rect 149734 100789 149746 101169
rect 150126 100789 150138 101169
rect 150518 100789 150530 101169
rect 150910 100789 150922 101169
rect 151302 100789 151314 101169
rect 151694 100789 151706 101169
rect 152086 100789 164442 101169
rect 164822 100789 164834 101169
rect 165214 100789 165226 101169
rect 165606 100789 165618 101169
rect 165998 100789 166010 101169
rect 166390 100789 166402 101169
rect 166782 100789 166794 101169
rect 167174 100789 167186 101169
rect 167566 100789 167578 101169
rect 167958 100789 168000 101169
rect 149220 100777 168000 100789
rect 149220 100397 149354 100777
rect 149734 100397 149746 100777
rect 150126 100397 150138 100777
rect 150518 100397 150530 100777
rect 150910 100397 150922 100777
rect 151302 100397 151314 100777
rect 151694 100397 151706 100777
rect 152086 100397 164442 100777
rect 164822 100397 164834 100777
rect 165214 100397 165226 100777
rect 165606 100397 165618 100777
rect 165998 100397 166010 100777
rect 166390 100397 166402 100777
rect 166782 100397 166794 100777
rect 167174 100397 167186 100777
rect 167566 100397 167578 100777
rect 167958 100397 168000 100777
rect 149220 100385 168000 100397
rect 149220 100005 149354 100385
rect 149734 100005 149746 100385
rect 150126 100005 150138 100385
rect 150518 100005 150530 100385
rect 150910 100005 150922 100385
rect 151302 100005 151314 100385
rect 151694 100005 151706 100385
rect 152086 100005 164442 100385
rect 164822 100005 164834 100385
rect 165214 100005 165226 100385
rect 165606 100005 165618 100385
rect 165998 100005 166010 100385
rect 166390 100005 166402 100385
rect 166782 100005 166794 100385
rect 167174 100005 167186 100385
rect 167566 100005 167578 100385
rect 167958 100005 168000 100385
rect 149220 99993 168000 100005
rect 149220 99613 149354 99993
rect 149734 99613 149746 99993
rect 150126 99613 150138 99993
rect 150518 99613 150530 99993
rect 150910 99613 150922 99993
rect 151302 99613 151314 99993
rect 151694 99613 151706 99993
rect 152086 99613 164442 99993
rect 164822 99613 164834 99993
rect 165214 99613 165226 99993
rect 165606 99613 165618 99993
rect 165998 99613 166010 99993
rect 166390 99613 166402 99993
rect 166782 99613 166794 99993
rect 167174 99613 167186 99993
rect 167566 99613 167578 99993
rect 167958 99613 168000 99993
rect 149220 99601 168000 99613
rect 149220 99221 149354 99601
rect 149734 99221 149746 99601
rect 150126 99221 150138 99601
rect 150518 99221 150530 99601
rect 150910 99221 150922 99601
rect 151302 99221 151314 99601
rect 151694 99221 151706 99601
rect 152086 99221 164442 99601
rect 164822 99221 164834 99601
rect 165214 99221 165226 99601
rect 165606 99221 165618 99601
rect 165998 99221 166010 99601
rect 166390 99221 166402 99601
rect 166782 99221 166794 99601
rect 167174 99221 167186 99601
rect 167566 99221 167578 99601
rect 167958 99221 168000 99601
rect 149220 99209 168000 99221
rect 149220 98829 149354 99209
rect 149734 98829 149746 99209
rect 150126 98829 150138 99209
rect 150518 98829 150530 99209
rect 150910 98829 150922 99209
rect 151302 98829 151314 99209
rect 151694 98829 151706 99209
rect 152086 98829 164442 99209
rect 164822 98829 164834 99209
rect 165214 98829 165226 99209
rect 165606 98829 165618 99209
rect 165998 98829 166010 99209
rect 166390 98829 166402 99209
rect 166782 98829 166794 99209
rect 167174 98829 167186 99209
rect 167566 98829 167578 99209
rect 167958 98829 168000 99209
rect 149220 98666 168000 98829
rect 196000 97000 210000 111000
rect 14000 81000 28000 95000
rect 67748 94870 156220 94900
rect 67748 94490 67882 94870
rect 68262 94490 68274 94870
rect 68654 94490 68666 94870
rect 69046 94490 69058 94870
rect 69438 94490 69450 94870
rect 69830 94490 69842 94870
rect 70222 94490 70234 94870
rect 70614 94490 79418 94870
rect 79798 94490 94538 94870
rect 94918 94490 109658 94870
rect 110038 94490 124778 94870
rect 125158 94490 139898 94870
rect 140278 94490 153354 94870
rect 153734 94490 153746 94870
rect 154126 94490 154138 94870
rect 154518 94490 154530 94870
rect 154910 94490 154922 94870
rect 155302 94490 155314 94870
rect 155694 94490 155706 94870
rect 156086 94490 156220 94870
rect 67748 94460 156220 94490
rect 71748 93630 152220 93660
rect 71748 93250 71882 93630
rect 72262 93250 72274 93630
rect 72654 93250 72666 93630
rect 73046 93250 73058 93630
rect 73438 93250 73450 93630
rect 73830 93250 73842 93630
rect 74222 93250 74234 93630
rect 74614 93250 78178 93630
rect 78558 93250 93298 93630
rect 93678 93250 108418 93630
rect 108798 93250 123538 93630
rect 123918 93250 138658 93630
rect 139038 93250 149354 93630
rect 149734 93250 149746 93630
rect 150126 93250 150138 93630
rect 150518 93250 150530 93630
rect 150910 93250 150922 93630
rect 151302 93250 151314 93630
rect 151694 93250 151706 93630
rect 152086 93250 152220 93630
rect 71748 93220 152220 93250
rect 60000 90501 70748 90664
rect 60000 90121 60042 90501
rect 60422 90121 60434 90501
rect 60814 90121 60826 90501
rect 61206 90121 61218 90501
rect 61598 90121 61610 90501
rect 61990 90121 62002 90501
rect 62382 90121 62394 90501
rect 62774 90121 62786 90501
rect 63166 90121 63178 90501
rect 63558 90121 67882 90501
rect 68262 90121 68274 90501
rect 68654 90121 68666 90501
rect 69046 90121 69058 90501
rect 69438 90121 69450 90501
rect 69830 90121 69842 90501
rect 70222 90121 70234 90501
rect 70614 90121 70748 90501
rect 60000 90109 70748 90121
rect 60000 89729 60042 90109
rect 60422 89729 60434 90109
rect 60814 89729 60826 90109
rect 61206 89729 61218 90109
rect 61598 89729 61610 90109
rect 61990 89729 62002 90109
rect 62382 89729 62394 90109
rect 62774 89729 62786 90109
rect 63166 89729 63178 90109
rect 63558 89729 67882 90109
rect 68262 89729 68274 90109
rect 68654 89729 68666 90109
rect 69046 89729 69058 90109
rect 69438 89729 69450 90109
rect 69830 89729 69842 90109
rect 70222 89729 70234 90109
rect 70614 89729 70748 90109
rect 60000 89717 70748 89729
rect 60000 89337 60042 89717
rect 60422 89337 60434 89717
rect 60814 89337 60826 89717
rect 61206 89337 61218 89717
rect 61598 89337 61610 89717
rect 61990 89337 62002 89717
rect 62382 89337 62394 89717
rect 62774 89337 62786 89717
rect 63166 89337 63178 89717
rect 63558 89337 67882 89717
rect 68262 89337 68274 89717
rect 68654 89337 68666 89717
rect 69046 89337 69058 89717
rect 69438 89337 69450 89717
rect 69830 89337 69842 89717
rect 70222 89337 70234 89717
rect 70614 89337 70748 89717
rect 60000 89325 70748 89337
rect 60000 88945 60042 89325
rect 60422 88945 60434 89325
rect 60814 88945 60826 89325
rect 61206 88945 61218 89325
rect 61598 88945 61610 89325
rect 61990 88945 62002 89325
rect 62382 88945 62394 89325
rect 62774 88945 62786 89325
rect 63166 88945 63178 89325
rect 63558 88945 67882 89325
rect 68262 88945 68274 89325
rect 68654 88945 68666 89325
rect 69046 88945 69058 89325
rect 69438 88945 69450 89325
rect 69830 88945 69842 89325
rect 70222 88945 70234 89325
rect 70614 88945 70748 89325
rect 60000 88933 70748 88945
rect 60000 88553 60042 88933
rect 60422 88553 60434 88933
rect 60814 88553 60826 88933
rect 61206 88553 61218 88933
rect 61598 88553 61610 88933
rect 61990 88553 62002 88933
rect 62382 88553 62394 88933
rect 62774 88553 62786 88933
rect 63166 88553 63178 88933
rect 63558 88553 67882 88933
rect 68262 88553 68274 88933
rect 68654 88553 68666 88933
rect 69046 88553 69058 88933
rect 69438 88553 69450 88933
rect 69830 88553 69842 88933
rect 70222 88553 70234 88933
rect 70614 88553 70748 88933
rect 60000 88541 70748 88553
rect 60000 88161 60042 88541
rect 60422 88161 60434 88541
rect 60814 88161 60826 88541
rect 61206 88161 61218 88541
rect 61598 88161 61610 88541
rect 61990 88161 62002 88541
rect 62382 88161 62394 88541
rect 62774 88161 62786 88541
rect 63166 88161 63178 88541
rect 63558 88161 67882 88541
rect 68262 88161 68274 88541
rect 68654 88161 68666 88541
rect 69046 88161 69058 88541
rect 69438 88161 69450 88541
rect 69830 88161 69842 88541
rect 70222 88161 70234 88541
rect 70614 88161 70748 88541
rect 60000 87998 70748 88161
rect 153220 90501 164000 90664
rect 153220 90121 153354 90501
rect 153734 90121 153746 90501
rect 154126 90121 154138 90501
rect 154518 90121 154530 90501
rect 154910 90121 154922 90501
rect 155302 90121 155314 90501
rect 155694 90121 155706 90501
rect 156086 90121 160442 90501
rect 160822 90121 160834 90501
rect 161214 90121 161226 90501
rect 161606 90121 161618 90501
rect 161998 90121 162010 90501
rect 162390 90121 162402 90501
rect 162782 90121 162794 90501
rect 163174 90121 163186 90501
rect 163566 90121 163578 90501
rect 163958 90121 164000 90501
rect 153220 90109 164000 90121
rect 153220 89729 153354 90109
rect 153734 89729 153746 90109
rect 154126 89729 154138 90109
rect 154518 89729 154530 90109
rect 154910 89729 154922 90109
rect 155302 89729 155314 90109
rect 155694 89729 155706 90109
rect 156086 89729 160442 90109
rect 160822 89729 160834 90109
rect 161214 89729 161226 90109
rect 161606 89729 161618 90109
rect 161998 89729 162010 90109
rect 162390 89729 162402 90109
rect 162782 89729 162794 90109
rect 163174 89729 163186 90109
rect 163566 89729 163578 90109
rect 163958 89729 164000 90109
rect 153220 89717 164000 89729
rect 153220 89337 153354 89717
rect 153734 89337 153746 89717
rect 154126 89337 154138 89717
rect 154518 89337 154530 89717
rect 154910 89337 154922 89717
rect 155302 89337 155314 89717
rect 155694 89337 155706 89717
rect 156086 89337 160442 89717
rect 160822 89337 160834 89717
rect 161214 89337 161226 89717
rect 161606 89337 161618 89717
rect 161998 89337 162010 89717
rect 162390 89337 162402 89717
rect 162782 89337 162794 89717
rect 163174 89337 163186 89717
rect 163566 89337 163578 89717
rect 163958 89337 164000 89717
rect 153220 89325 164000 89337
rect 153220 88945 153354 89325
rect 153734 88945 153746 89325
rect 154126 88945 154138 89325
rect 154518 88945 154530 89325
rect 154910 88945 154922 89325
rect 155302 88945 155314 89325
rect 155694 88945 155706 89325
rect 156086 88945 160442 89325
rect 160822 88945 160834 89325
rect 161214 88945 161226 89325
rect 161606 88945 161618 89325
rect 161998 88945 162010 89325
rect 162390 88945 162402 89325
rect 162782 88945 162794 89325
rect 163174 88945 163186 89325
rect 163566 88945 163578 89325
rect 163958 88945 164000 89325
rect 153220 88933 164000 88945
rect 153220 88553 153354 88933
rect 153734 88553 153746 88933
rect 154126 88553 154138 88933
rect 154518 88553 154530 88933
rect 154910 88553 154922 88933
rect 155302 88553 155314 88933
rect 155694 88553 155706 88933
rect 156086 88553 160442 88933
rect 160822 88553 160834 88933
rect 161214 88553 161226 88933
rect 161606 88553 161618 88933
rect 161998 88553 162010 88933
rect 162390 88553 162402 88933
rect 162782 88553 162794 88933
rect 163174 88553 163186 88933
rect 163566 88553 163578 88933
rect 163958 88553 164000 88933
rect 153220 88541 164000 88553
rect 153220 88161 153354 88541
rect 153734 88161 153746 88541
rect 154126 88161 154138 88541
rect 154518 88161 154530 88541
rect 154910 88161 154922 88541
rect 155302 88161 155314 88541
rect 155694 88161 155706 88541
rect 156086 88161 160442 88541
rect 160822 88161 160834 88541
rect 161214 88161 161226 88541
rect 161606 88161 161618 88541
rect 161998 88161 162010 88541
rect 162390 88161 162402 88541
rect 162782 88161 162794 88541
rect 163174 88161 163186 88541
rect 163566 88161 163578 88541
rect 163958 88161 164000 88541
rect 153220 87998 164000 88161
rect 56000 85169 74748 85332
rect 56000 84789 56042 85169
rect 56422 84789 56434 85169
rect 56814 84789 56826 85169
rect 57206 84789 57218 85169
rect 57598 84789 57610 85169
rect 57990 84789 58002 85169
rect 58382 84789 58394 85169
rect 58774 84789 58786 85169
rect 59166 84789 59178 85169
rect 59558 84789 71882 85169
rect 72262 84789 72274 85169
rect 72654 84789 72666 85169
rect 73046 84789 73058 85169
rect 73438 84789 73450 85169
rect 73830 84789 73842 85169
rect 74222 84789 74234 85169
rect 74614 84789 74748 85169
rect 56000 84777 74748 84789
rect 56000 84397 56042 84777
rect 56422 84397 56434 84777
rect 56814 84397 56826 84777
rect 57206 84397 57218 84777
rect 57598 84397 57610 84777
rect 57990 84397 58002 84777
rect 58382 84397 58394 84777
rect 58774 84397 58786 84777
rect 59166 84397 59178 84777
rect 59558 84397 71882 84777
rect 72262 84397 72274 84777
rect 72654 84397 72666 84777
rect 73046 84397 73058 84777
rect 73438 84397 73450 84777
rect 73830 84397 73842 84777
rect 74222 84397 74234 84777
rect 74614 84397 74748 84777
rect 56000 84385 74748 84397
rect 56000 84005 56042 84385
rect 56422 84005 56434 84385
rect 56814 84005 56826 84385
rect 57206 84005 57218 84385
rect 57598 84005 57610 84385
rect 57990 84005 58002 84385
rect 58382 84005 58394 84385
rect 58774 84005 58786 84385
rect 59166 84005 59178 84385
rect 59558 84005 71882 84385
rect 72262 84005 72274 84385
rect 72654 84005 72666 84385
rect 73046 84005 73058 84385
rect 73438 84005 73450 84385
rect 73830 84005 73842 84385
rect 74222 84005 74234 84385
rect 74614 84005 74748 84385
rect 56000 83993 74748 84005
rect 56000 83613 56042 83993
rect 56422 83613 56434 83993
rect 56814 83613 56826 83993
rect 57206 83613 57218 83993
rect 57598 83613 57610 83993
rect 57990 83613 58002 83993
rect 58382 83613 58394 83993
rect 58774 83613 58786 83993
rect 59166 83613 59178 83993
rect 59558 83613 71882 83993
rect 72262 83613 72274 83993
rect 72654 83613 72666 83993
rect 73046 83613 73058 83993
rect 73438 83613 73450 83993
rect 73830 83613 73842 83993
rect 74222 83613 74234 83993
rect 74614 83613 74748 83993
rect 56000 83601 74748 83613
rect 56000 83221 56042 83601
rect 56422 83221 56434 83601
rect 56814 83221 56826 83601
rect 57206 83221 57218 83601
rect 57598 83221 57610 83601
rect 57990 83221 58002 83601
rect 58382 83221 58394 83601
rect 58774 83221 58786 83601
rect 59166 83221 59178 83601
rect 59558 83221 71882 83601
rect 72262 83221 72274 83601
rect 72654 83221 72666 83601
rect 73046 83221 73058 83601
rect 73438 83221 73450 83601
rect 73830 83221 73842 83601
rect 74222 83221 74234 83601
rect 74614 83221 74748 83601
rect 56000 83209 74748 83221
rect 56000 82829 56042 83209
rect 56422 82829 56434 83209
rect 56814 82829 56826 83209
rect 57206 82829 57218 83209
rect 57598 82829 57610 83209
rect 57990 82829 58002 83209
rect 58382 82829 58394 83209
rect 58774 82829 58786 83209
rect 59166 82829 59178 83209
rect 59558 82829 71882 83209
rect 72262 82829 72274 83209
rect 72654 82829 72666 83209
rect 73046 82829 73058 83209
rect 73438 82829 73450 83209
rect 73830 82829 73842 83209
rect 74222 82829 74234 83209
rect 74614 82829 74748 83209
rect 56000 82666 74748 82829
rect 149220 85169 168000 85332
rect 149220 84789 149354 85169
rect 149734 84789 149746 85169
rect 150126 84789 150138 85169
rect 150518 84789 150530 85169
rect 150910 84789 150922 85169
rect 151302 84789 151314 85169
rect 151694 84789 151706 85169
rect 152086 84789 164442 85169
rect 164822 84789 164834 85169
rect 165214 84789 165226 85169
rect 165606 84789 165618 85169
rect 165998 84789 166010 85169
rect 166390 84789 166402 85169
rect 166782 84789 166794 85169
rect 167174 84789 167186 85169
rect 167566 84789 167578 85169
rect 167958 84789 168000 85169
rect 149220 84777 168000 84789
rect 149220 84397 149354 84777
rect 149734 84397 149746 84777
rect 150126 84397 150138 84777
rect 150518 84397 150530 84777
rect 150910 84397 150922 84777
rect 151302 84397 151314 84777
rect 151694 84397 151706 84777
rect 152086 84397 164442 84777
rect 164822 84397 164834 84777
rect 165214 84397 165226 84777
rect 165606 84397 165618 84777
rect 165998 84397 166010 84777
rect 166390 84397 166402 84777
rect 166782 84397 166794 84777
rect 167174 84397 167186 84777
rect 167566 84397 167578 84777
rect 167958 84397 168000 84777
rect 149220 84385 168000 84397
rect 149220 84005 149354 84385
rect 149734 84005 149746 84385
rect 150126 84005 150138 84385
rect 150518 84005 150530 84385
rect 150910 84005 150922 84385
rect 151302 84005 151314 84385
rect 151694 84005 151706 84385
rect 152086 84005 164442 84385
rect 164822 84005 164834 84385
rect 165214 84005 165226 84385
rect 165606 84005 165618 84385
rect 165998 84005 166010 84385
rect 166390 84005 166402 84385
rect 166782 84005 166794 84385
rect 167174 84005 167186 84385
rect 167566 84005 167578 84385
rect 167958 84005 168000 84385
rect 149220 83993 168000 84005
rect 149220 83613 149354 83993
rect 149734 83613 149746 83993
rect 150126 83613 150138 83993
rect 150518 83613 150530 83993
rect 150910 83613 150922 83993
rect 151302 83613 151314 83993
rect 151694 83613 151706 83993
rect 152086 83613 164442 83993
rect 164822 83613 164834 83993
rect 165214 83613 165226 83993
rect 165606 83613 165618 83993
rect 165998 83613 166010 83993
rect 166390 83613 166402 83993
rect 166782 83613 166794 83993
rect 167174 83613 167186 83993
rect 167566 83613 167578 83993
rect 167958 83613 168000 83993
rect 149220 83601 168000 83613
rect 149220 83221 149354 83601
rect 149734 83221 149746 83601
rect 150126 83221 150138 83601
rect 150518 83221 150530 83601
rect 150910 83221 150922 83601
rect 151302 83221 151314 83601
rect 151694 83221 151706 83601
rect 152086 83221 164442 83601
rect 164822 83221 164834 83601
rect 165214 83221 165226 83601
rect 165606 83221 165618 83601
rect 165998 83221 166010 83601
rect 166390 83221 166402 83601
rect 166782 83221 166794 83601
rect 167174 83221 167186 83601
rect 167566 83221 167578 83601
rect 167958 83221 168000 83601
rect 149220 83209 168000 83221
rect 149220 82829 149354 83209
rect 149734 82829 149746 83209
rect 150126 82829 150138 83209
rect 150518 82829 150530 83209
rect 150910 82829 150922 83209
rect 151302 82829 151314 83209
rect 151694 82829 151706 83209
rect 152086 82829 164442 83209
rect 164822 82829 164834 83209
rect 165214 82829 165226 83209
rect 165606 82829 165618 83209
rect 165998 82829 166010 83209
rect 166390 82829 166402 83209
rect 166782 82829 166794 83209
rect 167174 82829 167186 83209
rect 167566 82829 167578 83209
rect 167958 82829 168000 83209
rect 149220 82666 168000 82829
rect 196000 81000 210000 95000
rect 67748 79750 156220 79780
rect 67748 79370 67882 79750
rect 68262 79370 68274 79750
rect 68654 79370 68666 79750
rect 69046 79370 69058 79750
rect 69438 79370 69450 79750
rect 69830 79370 69842 79750
rect 70222 79370 70234 79750
rect 70614 79370 79418 79750
rect 79798 79370 94538 79750
rect 94918 79370 109658 79750
rect 110038 79370 124778 79750
rect 125158 79370 139898 79750
rect 140278 79370 153354 79750
rect 153734 79370 153746 79750
rect 154126 79370 154138 79750
rect 154518 79370 154530 79750
rect 154910 79370 154922 79750
rect 155302 79370 155314 79750
rect 155694 79370 155706 79750
rect 156086 79370 156220 79750
rect 67748 79340 156220 79370
rect 14000 65000 28000 79000
rect 71748 78510 152220 78540
rect 71748 78130 71882 78510
rect 72262 78130 72274 78510
rect 72654 78130 72666 78510
rect 73046 78130 73058 78510
rect 73438 78130 73450 78510
rect 73830 78130 73842 78510
rect 74222 78130 74234 78510
rect 74614 78130 78178 78510
rect 78558 78130 93298 78510
rect 93678 78130 108418 78510
rect 108798 78130 123538 78510
rect 123918 78130 138658 78510
rect 139038 78130 149354 78510
rect 149734 78130 149746 78510
rect 150126 78130 150138 78510
rect 150518 78130 150530 78510
rect 150910 78130 150922 78510
rect 151302 78130 151314 78510
rect 151694 78130 151706 78510
rect 152086 78130 152220 78510
rect 71748 78100 152220 78130
rect 60000 74501 70748 74664
rect 60000 74121 60042 74501
rect 60422 74121 60434 74501
rect 60814 74121 60826 74501
rect 61206 74121 61218 74501
rect 61598 74121 61610 74501
rect 61990 74121 62002 74501
rect 62382 74121 62394 74501
rect 62774 74121 62786 74501
rect 63166 74121 63178 74501
rect 63558 74121 67882 74501
rect 68262 74121 68274 74501
rect 68654 74121 68666 74501
rect 69046 74121 69058 74501
rect 69438 74121 69450 74501
rect 69830 74121 69842 74501
rect 70222 74121 70234 74501
rect 70614 74121 70748 74501
rect 60000 74109 70748 74121
rect 60000 73729 60042 74109
rect 60422 73729 60434 74109
rect 60814 73729 60826 74109
rect 61206 73729 61218 74109
rect 61598 73729 61610 74109
rect 61990 73729 62002 74109
rect 62382 73729 62394 74109
rect 62774 73729 62786 74109
rect 63166 73729 63178 74109
rect 63558 73729 67882 74109
rect 68262 73729 68274 74109
rect 68654 73729 68666 74109
rect 69046 73729 69058 74109
rect 69438 73729 69450 74109
rect 69830 73729 69842 74109
rect 70222 73729 70234 74109
rect 70614 73729 70748 74109
rect 60000 73717 70748 73729
rect 60000 73337 60042 73717
rect 60422 73337 60434 73717
rect 60814 73337 60826 73717
rect 61206 73337 61218 73717
rect 61598 73337 61610 73717
rect 61990 73337 62002 73717
rect 62382 73337 62394 73717
rect 62774 73337 62786 73717
rect 63166 73337 63178 73717
rect 63558 73337 67882 73717
rect 68262 73337 68274 73717
rect 68654 73337 68666 73717
rect 69046 73337 69058 73717
rect 69438 73337 69450 73717
rect 69830 73337 69842 73717
rect 70222 73337 70234 73717
rect 70614 73337 70748 73717
rect 60000 73325 70748 73337
rect 60000 72945 60042 73325
rect 60422 72945 60434 73325
rect 60814 72945 60826 73325
rect 61206 72945 61218 73325
rect 61598 72945 61610 73325
rect 61990 72945 62002 73325
rect 62382 72945 62394 73325
rect 62774 72945 62786 73325
rect 63166 72945 63178 73325
rect 63558 72945 67882 73325
rect 68262 72945 68274 73325
rect 68654 72945 68666 73325
rect 69046 72945 69058 73325
rect 69438 72945 69450 73325
rect 69830 72945 69842 73325
rect 70222 72945 70234 73325
rect 70614 72945 70748 73325
rect 60000 72933 70748 72945
rect 60000 72553 60042 72933
rect 60422 72553 60434 72933
rect 60814 72553 60826 72933
rect 61206 72553 61218 72933
rect 61598 72553 61610 72933
rect 61990 72553 62002 72933
rect 62382 72553 62394 72933
rect 62774 72553 62786 72933
rect 63166 72553 63178 72933
rect 63558 72553 67882 72933
rect 68262 72553 68274 72933
rect 68654 72553 68666 72933
rect 69046 72553 69058 72933
rect 69438 72553 69450 72933
rect 69830 72553 69842 72933
rect 70222 72553 70234 72933
rect 70614 72553 70748 72933
rect 60000 72541 70748 72553
rect 60000 72161 60042 72541
rect 60422 72161 60434 72541
rect 60814 72161 60826 72541
rect 61206 72161 61218 72541
rect 61598 72161 61610 72541
rect 61990 72161 62002 72541
rect 62382 72161 62394 72541
rect 62774 72161 62786 72541
rect 63166 72161 63178 72541
rect 63558 72161 67882 72541
rect 68262 72161 68274 72541
rect 68654 72161 68666 72541
rect 69046 72161 69058 72541
rect 69438 72161 69450 72541
rect 69830 72161 69842 72541
rect 70222 72161 70234 72541
rect 70614 72161 70748 72541
rect 60000 71998 70748 72161
rect 71748 74566 152220 74700
rect 71748 74186 71882 74566
rect 72262 74186 72274 74566
rect 72654 74186 72666 74566
rect 73046 74186 73058 74566
rect 73438 74186 73450 74566
rect 73830 74186 73842 74566
rect 74222 74186 74234 74566
rect 74614 74186 78178 74566
rect 78558 74186 93298 74566
rect 93678 74186 108418 74566
rect 108798 74186 123538 74566
rect 123918 74186 138658 74566
rect 139038 74186 149354 74566
rect 149734 74186 149746 74566
rect 150126 74186 150138 74566
rect 150518 74186 150530 74566
rect 150910 74186 150922 74566
rect 151302 74186 151314 74566
rect 151694 74186 151706 74566
rect 152086 74186 152220 74566
rect 71748 74174 152220 74186
rect 71748 73794 71882 74174
rect 72262 73794 72274 74174
rect 72654 73794 72666 74174
rect 73046 73794 73058 74174
rect 73438 73794 73450 74174
rect 73830 73794 73842 74174
rect 74222 73794 74234 74174
rect 74614 73794 78178 74174
rect 78558 73794 93298 74174
rect 93678 73794 108418 74174
rect 108798 73794 123538 74174
rect 123918 73794 138658 74174
rect 139038 73794 149354 74174
rect 149734 73794 149746 74174
rect 150126 73794 150138 74174
rect 150518 73794 150530 74174
rect 150910 73794 150922 74174
rect 151302 73794 151314 74174
rect 151694 73794 151706 74174
rect 152086 73794 152220 74174
rect 71748 73782 152220 73794
rect 71748 73402 71882 73782
rect 72262 73402 72274 73782
rect 72654 73402 72666 73782
rect 73046 73402 73058 73782
rect 73438 73402 73450 73782
rect 73830 73402 73842 73782
rect 74222 73402 74234 73782
rect 74614 73402 78178 73782
rect 78558 73402 93298 73782
rect 93678 73402 108418 73782
rect 108798 73402 123538 73782
rect 123918 73402 138658 73782
rect 139038 73402 149354 73782
rect 149734 73402 149746 73782
rect 150126 73402 150138 73782
rect 150518 73402 150530 73782
rect 150910 73402 150922 73782
rect 151302 73402 151314 73782
rect 151694 73402 151706 73782
rect 152086 73402 152220 73782
rect 71748 73390 152220 73402
rect 71748 73010 71882 73390
rect 72262 73010 72274 73390
rect 72654 73010 72666 73390
rect 73046 73010 73058 73390
rect 73438 73010 73450 73390
rect 73830 73010 73842 73390
rect 74222 73010 74234 73390
rect 74614 73010 78178 73390
rect 78558 73010 93298 73390
rect 93678 73010 108418 73390
rect 108798 73010 123538 73390
rect 123918 73010 138658 73390
rect 139038 73010 149354 73390
rect 149734 73010 149746 73390
rect 150126 73010 150138 73390
rect 150518 73010 150530 73390
rect 150910 73010 150922 73390
rect 151302 73010 151314 73390
rect 151694 73010 151706 73390
rect 152086 73010 152220 73390
rect 71748 72998 152220 73010
rect 71748 72618 71882 72998
rect 72262 72618 72274 72998
rect 72654 72618 72666 72998
rect 73046 72618 73058 72998
rect 73438 72618 73450 72998
rect 73830 72618 73842 72998
rect 74222 72618 74234 72998
rect 74614 72618 78178 72998
rect 78558 72618 93298 72998
rect 93678 72618 108418 72998
rect 108798 72618 123538 72998
rect 123918 72618 138658 72998
rect 139038 72618 149354 72998
rect 149734 72618 149746 72998
rect 150126 72618 150138 72998
rect 150518 72618 150530 72998
rect 150910 72618 150922 72998
rect 151302 72618 151314 72998
rect 151694 72618 151706 72998
rect 152086 72618 152220 72998
rect 71748 72606 152220 72618
rect 71748 72226 71882 72606
rect 72262 72226 72274 72606
rect 72654 72226 72666 72606
rect 73046 72226 73058 72606
rect 73438 72226 73450 72606
rect 73830 72226 73842 72606
rect 74222 72226 74234 72606
rect 74614 72226 78178 72606
rect 78558 72226 93298 72606
rect 93678 72226 108418 72606
rect 108798 72226 123538 72606
rect 123918 72226 138658 72606
rect 139038 72226 149354 72606
rect 149734 72226 149746 72606
rect 150126 72226 150138 72606
rect 150518 72226 150530 72606
rect 150910 72226 150922 72606
rect 151302 72226 151314 72606
rect 151694 72226 151706 72606
rect 152086 72226 152220 72606
rect 71748 72214 152220 72226
rect 71748 71834 71882 72214
rect 72262 71834 72274 72214
rect 72654 71834 72666 72214
rect 73046 71834 73058 72214
rect 73438 71834 73450 72214
rect 73830 71834 73842 72214
rect 74222 71834 74234 72214
rect 74614 71834 78178 72214
rect 78558 71834 93298 72214
rect 93678 71834 108418 72214
rect 108798 71834 123538 72214
rect 123918 71834 138658 72214
rect 139038 71834 149354 72214
rect 149734 71834 149746 72214
rect 150126 71834 150138 72214
rect 150518 71834 150530 72214
rect 150910 71834 150922 72214
rect 151302 71834 151314 72214
rect 151694 71834 151706 72214
rect 152086 71834 152220 72214
rect 153220 74501 164000 74664
rect 153220 74121 153354 74501
rect 153734 74121 153746 74501
rect 154126 74121 154138 74501
rect 154518 74121 154530 74501
rect 154910 74121 154922 74501
rect 155302 74121 155314 74501
rect 155694 74121 155706 74501
rect 156086 74121 160442 74501
rect 160822 74121 160834 74501
rect 161214 74121 161226 74501
rect 161606 74121 161618 74501
rect 161998 74121 162010 74501
rect 162390 74121 162402 74501
rect 162782 74121 162794 74501
rect 163174 74121 163186 74501
rect 163566 74121 163578 74501
rect 163958 74121 164000 74501
rect 153220 74109 164000 74121
rect 153220 73729 153354 74109
rect 153734 73729 153746 74109
rect 154126 73729 154138 74109
rect 154518 73729 154530 74109
rect 154910 73729 154922 74109
rect 155302 73729 155314 74109
rect 155694 73729 155706 74109
rect 156086 73729 160442 74109
rect 160822 73729 160834 74109
rect 161214 73729 161226 74109
rect 161606 73729 161618 74109
rect 161998 73729 162010 74109
rect 162390 73729 162402 74109
rect 162782 73729 162794 74109
rect 163174 73729 163186 74109
rect 163566 73729 163578 74109
rect 163958 73729 164000 74109
rect 153220 73717 164000 73729
rect 153220 73337 153354 73717
rect 153734 73337 153746 73717
rect 154126 73337 154138 73717
rect 154518 73337 154530 73717
rect 154910 73337 154922 73717
rect 155302 73337 155314 73717
rect 155694 73337 155706 73717
rect 156086 73337 160442 73717
rect 160822 73337 160834 73717
rect 161214 73337 161226 73717
rect 161606 73337 161618 73717
rect 161998 73337 162010 73717
rect 162390 73337 162402 73717
rect 162782 73337 162794 73717
rect 163174 73337 163186 73717
rect 163566 73337 163578 73717
rect 163958 73337 164000 73717
rect 153220 73325 164000 73337
rect 153220 72945 153354 73325
rect 153734 72945 153746 73325
rect 154126 72945 154138 73325
rect 154518 72945 154530 73325
rect 154910 72945 154922 73325
rect 155302 72945 155314 73325
rect 155694 72945 155706 73325
rect 156086 72945 160442 73325
rect 160822 72945 160834 73325
rect 161214 72945 161226 73325
rect 161606 72945 161618 73325
rect 161998 72945 162010 73325
rect 162390 72945 162402 73325
rect 162782 72945 162794 73325
rect 163174 72945 163186 73325
rect 163566 72945 163578 73325
rect 163958 72945 164000 73325
rect 153220 72933 164000 72945
rect 153220 72553 153354 72933
rect 153734 72553 153746 72933
rect 154126 72553 154138 72933
rect 154518 72553 154530 72933
rect 154910 72553 154922 72933
rect 155302 72553 155314 72933
rect 155694 72553 155706 72933
rect 156086 72553 160442 72933
rect 160822 72553 160834 72933
rect 161214 72553 161226 72933
rect 161606 72553 161618 72933
rect 161998 72553 162010 72933
rect 162390 72553 162402 72933
rect 162782 72553 162794 72933
rect 163174 72553 163186 72933
rect 163566 72553 163578 72933
rect 163958 72553 164000 72933
rect 153220 72541 164000 72553
rect 153220 72161 153354 72541
rect 153734 72161 153746 72541
rect 154126 72161 154138 72541
rect 154518 72161 154530 72541
rect 154910 72161 154922 72541
rect 155302 72161 155314 72541
rect 155694 72161 155706 72541
rect 156086 72161 160442 72541
rect 160822 72161 160834 72541
rect 161214 72161 161226 72541
rect 161606 72161 161618 72541
rect 161998 72161 162010 72541
rect 162390 72161 162402 72541
rect 162782 72161 162794 72541
rect 163174 72161 163186 72541
rect 163566 72161 163578 72541
rect 163958 72161 164000 72541
rect 153220 71998 164000 72161
rect 71748 71700 152220 71834
rect 67748 70566 156220 70700
rect 67748 70186 67882 70566
rect 68262 70186 68274 70566
rect 68654 70186 68666 70566
rect 69046 70186 69058 70566
rect 69438 70186 69450 70566
rect 69830 70186 69842 70566
rect 70222 70186 70234 70566
rect 70614 70186 79418 70566
rect 79798 70186 94538 70566
rect 94918 70186 109658 70566
rect 110038 70186 124778 70566
rect 125158 70186 139898 70566
rect 140278 70186 153354 70566
rect 153734 70186 153746 70566
rect 154126 70186 154138 70566
rect 154518 70186 154530 70566
rect 154910 70186 154922 70566
rect 155302 70186 155314 70566
rect 155694 70186 155706 70566
rect 156086 70186 156220 70566
rect 67748 70174 156220 70186
rect 67748 69794 67882 70174
rect 68262 69794 68274 70174
rect 68654 69794 68666 70174
rect 69046 69794 69058 70174
rect 69438 69794 69450 70174
rect 69830 69794 69842 70174
rect 70222 69794 70234 70174
rect 70614 69794 79418 70174
rect 79798 69794 94538 70174
rect 94918 69794 109658 70174
rect 110038 69794 124778 70174
rect 125158 69794 139898 70174
rect 140278 69794 153354 70174
rect 153734 69794 153746 70174
rect 154126 69794 154138 70174
rect 154518 69794 154530 70174
rect 154910 69794 154922 70174
rect 155302 69794 155314 70174
rect 155694 69794 155706 70174
rect 156086 69794 156220 70174
rect 67748 69782 156220 69794
rect 67748 69402 67882 69782
rect 68262 69402 68274 69782
rect 68654 69402 68666 69782
rect 69046 69402 69058 69782
rect 69438 69402 69450 69782
rect 69830 69402 69842 69782
rect 70222 69402 70234 69782
rect 70614 69402 79418 69782
rect 79798 69402 94538 69782
rect 94918 69402 109658 69782
rect 110038 69402 124778 69782
rect 125158 69402 139898 69782
rect 140278 69402 153354 69782
rect 153734 69402 153746 69782
rect 154126 69402 154138 69782
rect 154518 69402 154530 69782
rect 154910 69402 154922 69782
rect 155302 69402 155314 69782
rect 155694 69402 155706 69782
rect 156086 69402 156220 69782
rect 67748 69390 156220 69402
rect 67748 69010 67882 69390
rect 68262 69010 68274 69390
rect 68654 69010 68666 69390
rect 69046 69010 69058 69390
rect 69438 69010 69450 69390
rect 69830 69010 69842 69390
rect 70222 69010 70234 69390
rect 70614 69010 79418 69390
rect 79798 69010 94538 69390
rect 94918 69010 109658 69390
rect 110038 69010 124778 69390
rect 125158 69010 139898 69390
rect 140278 69010 153354 69390
rect 153734 69010 153746 69390
rect 154126 69010 154138 69390
rect 154518 69010 154530 69390
rect 154910 69010 154922 69390
rect 155302 69010 155314 69390
rect 155694 69010 155706 69390
rect 156086 69010 156220 69390
rect 67748 68998 156220 69010
rect 67748 68618 67882 68998
rect 68262 68618 68274 68998
rect 68654 68618 68666 68998
rect 69046 68618 69058 68998
rect 69438 68618 69450 68998
rect 69830 68618 69842 68998
rect 70222 68618 70234 68998
rect 70614 68618 79418 68998
rect 79798 68618 94538 68998
rect 94918 68618 109658 68998
rect 110038 68618 124778 68998
rect 125158 68618 139898 68998
rect 140278 68618 153354 68998
rect 153734 68618 153746 68998
rect 154126 68618 154138 68998
rect 154518 68618 154530 68998
rect 154910 68618 154922 68998
rect 155302 68618 155314 68998
rect 155694 68618 155706 68998
rect 156086 68618 156220 68998
rect 67748 68606 156220 68618
rect 67748 68226 67882 68606
rect 68262 68226 68274 68606
rect 68654 68226 68666 68606
rect 69046 68226 69058 68606
rect 69438 68226 69450 68606
rect 69830 68226 69842 68606
rect 70222 68226 70234 68606
rect 70614 68226 79418 68606
rect 79798 68226 94538 68606
rect 94918 68226 109658 68606
rect 110038 68226 124778 68606
rect 125158 68226 139898 68606
rect 140278 68226 153354 68606
rect 153734 68226 153746 68606
rect 154126 68226 154138 68606
rect 154518 68226 154530 68606
rect 154910 68226 154922 68606
rect 155302 68226 155314 68606
rect 155694 68226 155706 68606
rect 156086 68226 156220 68606
rect 67748 68214 156220 68226
rect 67748 67834 67882 68214
rect 68262 67834 68274 68214
rect 68654 67834 68666 68214
rect 69046 67834 69058 68214
rect 69438 67834 69450 68214
rect 69830 67834 69842 68214
rect 70222 67834 70234 68214
rect 70614 67834 79418 68214
rect 79798 67834 94538 68214
rect 94918 67834 109658 68214
rect 110038 67834 124778 68214
rect 125158 67834 139898 68214
rect 140278 67834 153354 68214
rect 153734 67834 153746 68214
rect 154126 67834 154138 68214
rect 154518 67834 154530 68214
rect 154910 67834 154922 68214
rect 155302 67834 155314 68214
rect 155694 67834 155706 68214
rect 156086 67834 156220 68214
rect 67748 67700 156220 67834
rect 196000 65000 210000 79000
rect 65000 14000 79000 28000
rect 81000 14000 95000 28000
rect 97000 14000 111000 28000
rect 113000 14000 127000 28000
rect 129000 14000 143000 28000
rect 145000 14000 159000 28000
use sg13g2_inv_1  _43_
timestamp 1676386529
transform -1 0 121248 0 -1 125496
box -48 -56 336 834
use sg13g2_inv_1  _44_
timestamp 1676386529
transform -1 0 122112 0 1 128520
box -48 -56 336 834
use sg13g2_inv_1  _45_
timestamp 1676386529
transform -1 0 118656 0 1 131544
box -48 -56 336 834
use sg13g2_inv_1  _46_
timestamp 1676386529
transform -1 0 101760 0 1 131544
box -48 -56 336 834
use sg13g2_inv_1  _47_
timestamp 1676386529
transform 1 0 102432 0 1 130032
box -48 -56 336 834
use sg13g2_nand4_1  _48_
timestamp 1685209130
transform -1 0 96000 0 -1 127008
box -48 -56 624 834
use sg13g2_nand4_1  _49_
timestamp 1685209130
transform 1 0 93792 0 1 128520
box -48 -56 624 834
use sg13g2_nor2_1  _50_
timestamp 1676630787
transform 1 0 97824 0 1 130032
box -48 -56 432 834
use sg13g2_nand4_1  _51_
timestamp 1685209130
transform -1 0 95040 0 -1 127008
box -48 -56 624 834
use sg13g2_nand4_1  _52_
timestamp 1685209130
transform -1 0 95040 0 1 127008
box -48 -56 624 834
use sg13g2_o21ai_1  _53_
timestamp 1685182643
transform -1 0 99648 0 1 131544
box -48 -56 538 834
use sg13g2_a21oi_1  _54_
timestamp 1683980220
transform 1 0 98496 0 -1 133056
box -48 -56 528 834
use sg13g2_a21oi_1  _55_
timestamp 1683980220
transform -1 0 101472 0 1 131544
box -48 -56 528 834
use sg13g2_nand2_1  _56_
timestamp 1676560849
transform 1 0 99936 0 1 131544
box -48 -56 432 834
use sg13g2_nor3_1  _57_
timestamp 1676643042
transform 1 0 97056 0 -1 130032
box -48 -56 528 834
use sg13g2_nor3_1  _58_
timestamp 1676643042
transform -1 0 102432 0 -1 131544
box -48 -56 528 834
use sg13g2_nor2_1  _59_
timestamp 1676630787
transform -1 0 103392 0 -1 130032
box -48 -56 432 834
use sg13g2_nor4_1  _60_
timestamp 1676646725
transform -1 0 99360 0 -1 128520
box -48 -56 624 834
use sg13g2_nor3_1  _61_
timestamp 1676643042
transform 1 0 102720 0 1 130032
box -48 -56 528 834
use sg13g2_nand3_1  _62_
timestamp 1683995554
transform -1 0 110880 0 1 130032
box -48 -56 528 834
use sg13g2_o21ai_1  _63_
timestamp 1685182643
transform -1 0 109248 0 -1 131544
box -48 -56 538 834
use sg13g2_nor2b_1  _64_
timestamp 1685188586
transform -1 0 109728 0 -1 131544
box -54 -56 528 834
use sg13g2_nand2b_1  _65_
timestamp 1676570795
transform -1 0 112704 0 -1 131544
box -48 -56 528 834
use sg13g2_nand4_1  _66_
timestamp 1685209130
transform 1 0 112128 0 1 131544
box -48 -56 624 834
use sg13g2_and3_1  _67_
timestamp 1676975269
transform 1 0 112800 0 -1 131544
box -48 -56 720 834
use sg13g2_nand4_1  _68_
timestamp 1685209130
transform 1 0 114816 0 -1 131544
box -48 -56 624 834
use sg13g2_nand2_1  _69_
timestamp 1676560849
transform 1 0 117408 0 1 130032
box -48 -56 432 834
use sg13g2_a21oi_1  _70_
timestamp 1683980220
transform -1 0 119520 0 -1 131544
box -48 -56 528 834
use sg13g2_o21ai_1  _71_
timestamp 1685182643
transform 1 0 118944 0 -1 128520
box -48 -56 538 834
use sg13g2_a21oi_1  _72_
timestamp 1683980220
transform -1 0 120000 0 -1 128520
box -48 -56 528 834
use sg13g2_o21ai_1  _73_
timestamp 1685182643
transform 1 0 118752 0 1 127008
box -48 -56 538 834
use sg13g2_or4_1  _74_
timestamp 1677158204
transform 1 0 118176 0 -1 128520
box -48 -56 816 834
use sg13g2_and3_1  _75_
timestamp 1676975269
transform 1 0 118848 0 1 125496
box -48 -56 720 834
use sg13g2_dfrbpq_1  _76_
timestamp 1746542328
transform 1 0 97344 0 -1 134568
box -48 -56 2640 834
use sg13g2_tiehi  _76__3
timestamp 1680007851
transform -1 0 98112 0 1 133056
box -48 -56 432 834
use sg13g2_dfrbpq_1  _77_
timestamp 1746542328
transform 1 0 103776 0 -1 133056
box -48 -56 2640 834
use sg13g2_tiehi  _77__10
timestamp 1680007851
transform -1 0 104640 0 1 131544
box -48 -56 432 834
use sg13g2_dfrbpq_1  _78_
timestamp 1746542328
transform 1 0 103488 0 -1 130032
box -48 -56 2640 834
use sg13g2_tiehi  _78__8
timestamp 1680007851
transform -1 0 104352 0 1 128520
box -48 -56 432 834
use sg13g2_tiehi  _79__6
timestamp 1680007851
transform -1 0 110208 0 -1 133056
box -48 -56 432 834
use sg13g2_dfrbpq_1  _79_
timestamp 1746542328
transform 1 0 109344 0 1 131544
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _80_
timestamp 1746542328
transform 1 0 113472 0 -1 134568
box -48 -56 2640 834
use sg13g2_tiehi  _80__4
timestamp 1680007851
transform -1 0 114336 0 1 133056
box -48 -56 432 834
use sg13g2_tiehi  _81__9
timestamp 1680007851
transform -1 0 120192 0 -1 134568
box -48 -56 432 834
use sg13g2_dfrbpq_1  _81_
timestamp 1746542328
transform 1 0 119328 0 1 133056
box -48 -56 2640 834
use sg13g2_tiehi  _82__5
timestamp 1680007851
transform -1 0 121536 0 1 128520
box -48 -56 432 834
use sg13g2_dfrbpq_1  _82_
timestamp 1746542328
transform 1 0 120672 0 -1 128520
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _83_
timestamp 1746542328
transform 1 0 119136 0 -1 123984
box -48 -56 2640 834
use sg13g2_tiehi  _83__7
timestamp 1680007851
transform -1 0 120000 0 1 122472
box -48 -56 432 834
use sg13g2_IOPadIn  clk_pad
timestamp 1716382777
transform 1 0 64000 0 1 28000
box -124 0 16124 36000
use sg13g2_buf_16  clkbuf_0_clk_PAD2CORE
timestamp 1676557096
transform -1 0 112800 0 -1 130032
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_0__f_clk_PAD2CORE
timestamp 1676557096
transform 1 0 108000 0 1 130032
box -48 -56 2448 834
use sg13g2_buf_16  clkbuf_1_1__f_clk_PAD2CORE
timestamp 1676557096
transform -1 0 116160 0 -1 130032
box -48 -56 2448 834
use sg13g2_decap_8  FILLER_0_0
timestamp 1679585382
transform 1 0 75648 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_7
timestamp 1679585382
transform 1 0 76320 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_14
timestamp 1679585382
transform 1 0 76992 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_21
timestamp 1679585382
transform 1 0 77664 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_28
timestamp 1679585382
transform 1 0 78336 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_35
timestamp 1679585382
transform 1 0 79008 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_42
timestamp 1679585382
transform 1 0 79680 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_49
timestamp 1679585382
transform 1 0 80352 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_56
timestamp 1679585382
transform 1 0 81024 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_63
timestamp 1679585382
transform 1 0 81696 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_70
timestamp 1679585382
transform 1 0 82368 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_77
timestamp 1679585382
transform 1 0 83040 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_84
timestamp 1679585382
transform 1 0 83712 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_91
timestamp 1679585382
transform 1 0 84384 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_98
timestamp 1679585382
transform 1 0 85056 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_105
timestamp 1679585382
transform 1 0 85728 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_112
timestamp 1679585382
transform 1 0 86400 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_119
timestamp 1679585382
transform 1 0 87072 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_126
timestamp 1679585382
transform 1 0 87744 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_133
timestamp 1679585382
transform 1 0 88416 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_140
timestamp 1679585382
transform 1 0 89088 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_147
timestamp 1679585382
transform 1 0 89760 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_154
timestamp 1679585382
transform 1 0 90432 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_161
timestamp 1679585382
transform 1 0 91104 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_168
timestamp 1679585382
transform 1 0 91776 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_175
timestamp 1679585382
transform 1 0 92448 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_182
timestamp 1679585382
transform 1 0 93120 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_189
timestamp 1679585382
transform 1 0 93792 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_196
timestamp 1679585382
transform 1 0 94464 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_203
timestamp 1679585382
transform 1 0 95136 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_210
timestamp 1679585382
transform 1 0 95808 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_217
timestamp 1679585382
transform 1 0 96480 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_224
timestamp 1679585382
transform 1 0 97152 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_231
timestamp 1679585382
transform 1 0 97824 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_238
timestamp 1679585382
transform 1 0 98496 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_245
timestamp 1679585382
transform 1 0 99168 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_252
timestamp 1679585382
transform 1 0 99840 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_259
timestamp 1679585382
transform 1 0 100512 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_266
timestamp 1679585382
transform 1 0 101184 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_273
timestamp 1679585382
transform 1 0 101856 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_280
timestamp 1679585382
transform 1 0 102528 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_287
timestamp 1679585382
transform 1 0 103200 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_294
timestamp 1679585382
transform 1 0 103872 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_301
timestamp 1679585382
transform 1 0 104544 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_308
timestamp 1679585382
transform 1 0 105216 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_315
timestamp 1679585382
transform 1 0 105888 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_322
timestamp 1679585382
transform 1 0 106560 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_329
timestamp 1679585382
transform 1 0 107232 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_336
timestamp 1679585382
transform 1 0 107904 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_343
timestamp 1679585382
transform 1 0 108576 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_350
timestamp 1679585382
transform 1 0 109248 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_357
timestamp 1679585382
transform 1 0 109920 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_364
timestamp 1679585382
transform 1 0 110592 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_371
timestamp 1679585382
transform 1 0 111264 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_378
timestamp 1679585382
transform 1 0 111936 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_385
timestamp 1679585382
transform 1 0 112608 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_392
timestamp 1679585382
transform 1 0 113280 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_399
timestamp 1679585382
transform 1 0 113952 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_406
timestamp 1679585382
transform 1 0 114624 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_413
timestamp 1679585382
transform 1 0 115296 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_420
timestamp 1679585382
transform 1 0 115968 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_427
timestamp 1679585382
transform 1 0 116640 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_434
timestamp 1679585382
transform 1 0 117312 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_441
timestamp 1679585382
transform 1 0 117984 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_448
timestamp 1679585382
transform 1 0 118656 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_455
timestamp 1679585382
transform 1 0 119328 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_462
timestamp 1679585382
transform 1 0 120000 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_469
timestamp 1679585382
transform 1 0 120672 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_476
timestamp 1679585382
transform 1 0 121344 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_483
timestamp 1679585382
transform 1 0 122016 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_490
timestamp 1679585382
transform 1 0 122688 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_497
timestamp 1679585382
transform 1 0 123360 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_504
timestamp 1679585382
transform 1 0 124032 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_511
timestamp 1679585382
transform 1 0 124704 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_518
timestamp 1679585382
transform 1 0 125376 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_525
timestamp 1679585382
transform 1 0 126048 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_532
timestamp 1679585382
transform 1 0 126720 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_539
timestamp 1679585382
transform 1 0 127392 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_546
timestamp 1679585382
transform 1 0 128064 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_553
timestamp 1679585382
transform 1 0 128736 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_560
timestamp 1679585382
transform 1 0 129408 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_567
timestamp 1679585382
transform 1 0 130080 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_574
timestamp 1679585382
transform 1 0 130752 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_581
timestamp 1679585382
transform 1 0 131424 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_588
timestamp 1679585382
transform 1 0 132096 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_595
timestamp 1679585382
transform 1 0 132768 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_602
timestamp 1679585382
transform 1 0 133440 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_609
timestamp 1679585382
transform 1 0 134112 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_616
timestamp 1679585382
transform 1 0 134784 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_623
timestamp 1679585382
transform 1 0 135456 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_630
timestamp 1679585382
transform 1 0 136128 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_637
timestamp 1679585382
transform 1 0 136800 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_644
timestamp 1679585382
transform 1 0 137472 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_651
timestamp 1679585382
transform 1 0 138144 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_658
timestamp 1679585382
transform 1 0 138816 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_665
timestamp 1679585382
transform 1 0 139488 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_672
timestamp 1679585382
transform 1 0 140160 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_679
timestamp 1679585382
transform 1 0 140832 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_686
timestamp 1679585382
transform 1 0 141504 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_693
timestamp 1679585382
transform 1 0 142176 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_700
timestamp 1679585382
transform 1 0 142848 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_707
timestamp 1679585382
transform 1 0 143520 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_714
timestamp 1679585382
transform 1 0 144192 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_721
timestamp 1679585382
transform 1 0 144864 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_728
timestamp 1679585382
transform 1 0 145536 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_735
timestamp 1679585382
transform 1 0 146208 0 1 75600
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_742
timestamp 1679585382
transform 1 0 146880 0 1 75600
box -48 -56 720 834
use sg13g2_decap_4  FILLER_0_749
timestamp 1679581501
transform 1 0 147552 0 1 75600
box -48 -56 432 834
use sg13g2_decap_8  FILLER_1_0
timestamp 1679585382
transform 1 0 75648 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_7
timestamp 1679585382
transform 1 0 76320 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_14
timestamp 1679585382
transform 1 0 76992 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_21
timestamp 1679585382
transform 1 0 77664 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_28
timestamp 1679585382
transform 1 0 78336 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_35
timestamp 1679585382
transform 1 0 79008 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_42
timestamp 1679585382
transform 1 0 79680 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_49
timestamp 1679585382
transform 1 0 80352 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_56
timestamp 1679585382
transform 1 0 81024 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_63
timestamp 1679585382
transform 1 0 81696 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_70
timestamp 1679585382
transform 1 0 82368 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_77
timestamp 1679585382
transform 1 0 83040 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_84
timestamp 1679585382
transform 1 0 83712 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_91
timestamp 1679585382
transform 1 0 84384 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_98
timestamp 1679585382
transform 1 0 85056 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_105
timestamp 1679585382
transform 1 0 85728 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_112
timestamp 1679585382
transform 1 0 86400 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_119
timestamp 1679585382
transform 1 0 87072 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_126
timestamp 1679585382
transform 1 0 87744 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_133
timestamp 1679585382
transform 1 0 88416 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_140
timestamp 1679585382
transform 1 0 89088 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_147
timestamp 1679585382
transform 1 0 89760 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_154
timestamp 1679585382
transform 1 0 90432 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_161
timestamp 1679585382
transform 1 0 91104 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_168
timestamp 1679585382
transform 1 0 91776 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_175
timestamp 1679585382
transform 1 0 92448 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_182
timestamp 1679585382
transform 1 0 93120 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_189
timestamp 1679585382
transform 1 0 93792 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679585382
transform 1 0 94464 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_203
timestamp 1679585382
transform 1 0 95136 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_210
timestamp 1679585382
transform 1 0 95808 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_217
timestamp 1679585382
transform 1 0 96480 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_224
timestamp 1679585382
transform 1 0 97152 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_231
timestamp 1679585382
transform 1 0 97824 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_238
timestamp 1679585382
transform 1 0 98496 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_245
timestamp 1679585382
transform 1 0 99168 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_252
timestamp 1679585382
transform 1 0 99840 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_259
timestamp 1679585382
transform 1 0 100512 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_266
timestamp 1679585382
transform 1 0 101184 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_273
timestamp 1679585382
transform 1 0 101856 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_280
timestamp 1679585382
transform 1 0 102528 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_287
timestamp 1679585382
transform 1 0 103200 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_294
timestamp 1679585382
transform 1 0 103872 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_301
timestamp 1679585382
transform 1 0 104544 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_308
timestamp 1679585382
transform 1 0 105216 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_315
timestamp 1679585382
transform 1 0 105888 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_322
timestamp 1679585382
transform 1 0 106560 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_329
timestamp 1679585382
transform 1 0 107232 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_336
timestamp 1679585382
transform 1 0 107904 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_343
timestamp 1679585382
transform 1 0 108576 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_350
timestamp 1679585382
transform 1 0 109248 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_357
timestamp 1679585382
transform 1 0 109920 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_364
timestamp 1679585382
transform 1 0 110592 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_371
timestamp 1679585382
transform 1 0 111264 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_378
timestamp 1679585382
transform 1 0 111936 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_385
timestamp 1679585382
transform 1 0 112608 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_392
timestamp 1679585382
transform 1 0 113280 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_399
timestamp 1679585382
transform 1 0 113952 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_406
timestamp 1679585382
transform 1 0 114624 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_413
timestamp 1679585382
transform 1 0 115296 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_420
timestamp 1679585382
transform 1 0 115968 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_427
timestamp 1679585382
transform 1 0 116640 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_434
timestamp 1679585382
transform 1 0 117312 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_441
timestamp 1679585382
transform 1 0 117984 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_448
timestamp 1679585382
transform 1 0 118656 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_455
timestamp 1679585382
transform 1 0 119328 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_462
timestamp 1679585382
transform 1 0 120000 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_469
timestamp 1679585382
transform 1 0 120672 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_476
timestamp 1679585382
transform 1 0 121344 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_483
timestamp 1679585382
transform 1 0 122016 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_490
timestamp 1679585382
transform 1 0 122688 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_497
timestamp 1679585382
transform 1 0 123360 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_504
timestamp 1679585382
transform 1 0 124032 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_511
timestamp 1679585382
transform 1 0 124704 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_518
timestamp 1679585382
transform 1 0 125376 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_525
timestamp 1679585382
transform 1 0 126048 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_532
timestamp 1679585382
transform 1 0 126720 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_539
timestamp 1679585382
transform 1 0 127392 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_546
timestamp 1679585382
transform 1 0 128064 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_553
timestamp 1679585382
transform 1 0 128736 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_560
timestamp 1679585382
transform 1 0 129408 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_567
timestamp 1679585382
transform 1 0 130080 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_574
timestamp 1679585382
transform 1 0 130752 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_581
timestamp 1679585382
transform 1 0 131424 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_588
timestamp 1679585382
transform 1 0 132096 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_595
timestamp 1679585382
transform 1 0 132768 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_602
timestamp 1679585382
transform 1 0 133440 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_609
timestamp 1679585382
transform 1 0 134112 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_616
timestamp 1679585382
transform 1 0 134784 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_623
timestamp 1679585382
transform 1 0 135456 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_630
timestamp 1679585382
transform 1 0 136128 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_637
timestamp 1679585382
transform 1 0 136800 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_644
timestamp 1679585382
transform 1 0 137472 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_651
timestamp 1679585382
transform 1 0 138144 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_658
timestamp 1679585382
transform 1 0 138816 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_665
timestamp 1679585382
transform 1 0 139488 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_672
timestamp 1679585382
transform 1 0 140160 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_679
timestamp 1679585382
transform 1 0 140832 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_686
timestamp 1679585382
transform 1 0 141504 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_693
timestamp 1679585382
transform 1 0 142176 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_700
timestamp 1679585382
transform 1 0 142848 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_707
timestamp 1679585382
transform 1 0 143520 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_714
timestamp 1679585382
transform 1 0 144192 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_721
timestamp 1679585382
transform 1 0 144864 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_728
timestamp 1679585382
transform 1 0 145536 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_735
timestamp 1679585382
transform 1 0 146208 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_742
timestamp 1679585382
transform 1 0 146880 0 -1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_1_749
timestamp 1679585382
transform 1 0 147552 0 -1 77112
box -48 -56 720 834
use sg13g2_fill_1  FILLER_1_756
timestamp 1677583258
transform 1 0 148224 0 -1 77112
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_0
timestamp 1679585382
transform 1 0 75648 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_7
timestamp 1679585382
transform 1 0 76320 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_14
timestamp 1679585382
transform 1 0 76992 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_21
timestamp 1679585382
transform 1 0 77664 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_28
timestamp 1679585382
transform 1 0 78336 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_35
timestamp 1679585382
transform 1 0 79008 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_42
timestamp 1679585382
transform 1 0 79680 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_49
timestamp 1679585382
transform 1 0 80352 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_56
timestamp 1679585382
transform 1 0 81024 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_63
timestamp 1679585382
transform 1 0 81696 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_70
timestamp 1679585382
transform 1 0 82368 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_77
timestamp 1679585382
transform 1 0 83040 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_84
timestamp 1679585382
transform 1 0 83712 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_91
timestamp 1679585382
transform 1 0 84384 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_98
timestamp 1679585382
transform 1 0 85056 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_105
timestamp 1679585382
transform 1 0 85728 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_112
timestamp 1679585382
transform 1 0 86400 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_119
timestamp 1679585382
transform 1 0 87072 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_126
timestamp 1679585382
transform 1 0 87744 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_133
timestamp 1679585382
transform 1 0 88416 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_140
timestamp 1679585382
transform 1 0 89088 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_147
timestamp 1679585382
transform 1 0 89760 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_154
timestamp 1679585382
transform 1 0 90432 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_161
timestamp 1679585382
transform 1 0 91104 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_168
timestamp 1679585382
transform 1 0 91776 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_175
timestamp 1679585382
transform 1 0 92448 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_182
timestamp 1679585382
transform 1 0 93120 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_189
timestamp 1679585382
transform 1 0 93792 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_196
timestamp 1679585382
transform 1 0 94464 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_203
timestamp 1679585382
transform 1 0 95136 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_210
timestamp 1679585382
transform 1 0 95808 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_217
timestamp 1679585382
transform 1 0 96480 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_224
timestamp 1679585382
transform 1 0 97152 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_231
timestamp 1679585382
transform 1 0 97824 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_238
timestamp 1679585382
transform 1 0 98496 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_245
timestamp 1679585382
transform 1 0 99168 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_252
timestamp 1679585382
transform 1 0 99840 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_259
timestamp 1679585382
transform 1 0 100512 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_266
timestamp 1679585382
transform 1 0 101184 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_273
timestamp 1679585382
transform 1 0 101856 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_280
timestamp 1679585382
transform 1 0 102528 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_287
timestamp 1679585382
transform 1 0 103200 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_294
timestamp 1679585382
transform 1 0 103872 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_301
timestamp 1679585382
transform 1 0 104544 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_308
timestamp 1679585382
transform 1 0 105216 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_315
timestamp 1679585382
transform 1 0 105888 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_322
timestamp 1679585382
transform 1 0 106560 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_329
timestamp 1679585382
transform 1 0 107232 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_336
timestamp 1679585382
transform 1 0 107904 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_343
timestamp 1679585382
transform 1 0 108576 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_350
timestamp 1679585382
transform 1 0 109248 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_357
timestamp 1679585382
transform 1 0 109920 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_364
timestamp 1679585382
transform 1 0 110592 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_371
timestamp 1679585382
transform 1 0 111264 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_378
timestamp 1679585382
transform 1 0 111936 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_385
timestamp 1679585382
transform 1 0 112608 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_392
timestamp 1679585382
transform 1 0 113280 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_399
timestamp 1679585382
transform 1 0 113952 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_406
timestamp 1679585382
transform 1 0 114624 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_413
timestamp 1679585382
transform 1 0 115296 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_420
timestamp 1679585382
transform 1 0 115968 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_427
timestamp 1679585382
transform 1 0 116640 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_434
timestamp 1679585382
transform 1 0 117312 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_441
timestamp 1679585382
transform 1 0 117984 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_448
timestamp 1679585382
transform 1 0 118656 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_455
timestamp 1679585382
transform 1 0 119328 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_462
timestamp 1679585382
transform 1 0 120000 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_469
timestamp 1679585382
transform 1 0 120672 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_476
timestamp 1679585382
transform 1 0 121344 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_483
timestamp 1679585382
transform 1 0 122016 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_490
timestamp 1679585382
transform 1 0 122688 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_497
timestamp 1679585382
transform 1 0 123360 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_504
timestamp 1679585382
transform 1 0 124032 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_511
timestamp 1679585382
transform 1 0 124704 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_518
timestamp 1679585382
transform 1 0 125376 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_525
timestamp 1679585382
transform 1 0 126048 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_532
timestamp 1679585382
transform 1 0 126720 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_539
timestamp 1679585382
transform 1 0 127392 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_546
timestamp 1679585382
transform 1 0 128064 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_553
timestamp 1679585382
transform 1 0 128736 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_560
timestamp 1679585382
transform 1 0 129408 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_567
timestamp 1679585382
transform 1 0 130080 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_574
timestamp 1679585382
transform 1 0 130752 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_581
timestamp 1679585382
transform 1 0 131424 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_588
timestamp 1679585382
transform 1 0 132096 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_595
timestamp 1679585382
transform 1 0 132768 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_602
timestamp 1679585382
transform 1 0 133440 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_609
timestamp 1679585382
transform 1 0 134112 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_616
timestamp 1679585382
transform 1 0 134784 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_623
timestamp 1679585382
transform 1 0 135456 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_630
timestamp 1679585382
transform 1 0 136128 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_637
timestamp 1679585382
transform 1 0 136800 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_644
timestamp 1679585382
transform 1 0 137472 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_651
timestamp 1679585382
transform 1 0 138144 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_658
timestamp 1679585382
transform 1 0 138816 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_665
timestamp 1679585382
transform 1 0 139488 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_672
timestamp 1679585382
transform 1 0 140160 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_679
timestamp 1679585382
transform 1 0 140832 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_686
timestamp 1679585382
transform 1 0 141504 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_693
timestamp 1679585382
transform 1 0 142176 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_700
timestamp 1679585382
transform 1 0 142848 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_707
timestamp 1679585382
transform 1 0 143520 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_714
timestamp 1679585382
transform 1 0 144192 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_721
timestamp 1679585382
transform 1 0 144864 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_728
timestamp 1679585382
transform 1 0 145536 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_735
timestamp 1679585382
transform 1 0 146208 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_742
timestamp 1679585382
transform 1 0 146880 0 1 77112
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_749
timestamp 1679585382
transform 1 0 147552 0 1 77112
box -48 -56 720 834
use sg13g2_fill_1  FILLER_2_756
timestamp 1677583258
transform 1 0 148224 0 1 77112
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_0
timestamp 1679585382
transform 1 0 75648 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_7
timestamp 1679585382
transform 1 0 76320 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_14
timestamp 1679585382
transform 1 0 76992 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_21
timestamp 1679585382
transform 1 0 77664 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_28
timestamp 1679585382
transform 1 0 78336 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_35
timestamp 1679585382
transform 1 0 79008 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_42
timestamp 1679585382
transform 1 0 79680 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_49
timestamp 1679585382
transform 1 0 80352 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_56
timestamp 1679585382
transform 1 0 81024 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_63
timestamp 1679585382
transform 1 0 81696 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_70
timestamp 1679585382
transform 1 0 82368 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_77
timestamp 1679585382
transform 1 0 83040 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_84
timestamp 1679585382
transform 1 0 83712 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_91
timestamp 1679585382
transform 1 0 84384 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_98
timestamp 1679585382
transform 1 0 85056 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_105
timestamp 1679585382
transform 1 0 85728 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_112
timestamp 1679585382
transform 1 0 86400 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_119
timestamp 1679585382
transform 1 0 87072 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_126
timestamp 1679585382
transform 1 0 87744 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_133
timestamp 1679585382
transform 1 0 88416 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_140
timestamp 1679585382
transform 1 0 89088 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_147
timestamp 1679585382
transform 1 0 89760 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_154
timestamp 1679585382
transform 1 0 90432 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_161
timestamp 1679585382
transform 1 0 91104 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_168
timestamp 1679585382
transform 1 0 91776 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_175
timestamp 1679585382
transform 1 0 92448 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_182
timestamp 1679585382
transform 1 0 93120 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_189
timestamp 1679585382
transform 1 0 93792 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_196
timestamp 1679585382
transform 1 0 94464 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_203
timestamp 1679585382
transform 1 0 95136 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_210
timestamp 1679585382
transform 1 0 95808 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_217
timestamp 1679585382
transform 1 0 96480 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_224
timestamp 1679585382
transform 1 0 97152 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_231
timestamp 1679585382
transform 1 0 97824 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_238
timestamp 1679585382
transform 1 0 98496 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_245
timestamp 1679585382
transform 1 0 99168 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_252
timestamp 1679585382
transform 1 0 99840 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_259
timestamp 1679585382
transform 1 0 100512 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_266
timestamp 1679585382
transform 1 0 101184 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_273
timestamp 1679585382
transform 1 0 101856 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_280
timestamp 1679585382
transform 1 0 102528 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_287
timestamp 1679585382
transform 1 0 103200 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_294
timestamp 1679585382
transform 1 0 103872 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_301
timestamp 1679585382
transform 1 0 104544 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_308
timestamp 1679585382
transform 1 0 105216 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_315
timestamp 1679585382
transform 1 0 105888 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_322
timestamp 1679585382
transform 1 0 106560 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_329
timestamp 1679585382
transform 1 0 107232 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_336
timestamp 1679585382
transform 1 0 107904 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_343
timestamp 1679585382
transform 1 0 108576 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_350
timestamp 1679585382
transform 1 0 109248 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_357
timestamp 1679585382
transform 1 0 109920 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_364
timestamp 1679585382
transform 1 0 110592 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_371
timestamp 1679585382
transform 1 0 111264 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_378
timestamp 1679585382
transform 1 0 111936 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_385
timestamp 1679585382
transform 1 0 112608 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_392
timestamp 1679585382
transform 1 0 113280 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_399
timestamp 1679585382
transform 1 0 113952 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_406
timestamp 1679585382
transform 1 0 114624 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_413
timestamp 1679585382
transform 1 0 115296 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_420
timestamp 1679585382
transform 1 0 115968 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_427
timestamp 1679585382
transform 1 0 116640 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_434
timestamp 1679585382
transform 1 0 117312 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_441
timestamp 1679585382
transform 1 0 117984 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_448
timestamp 1679585382
transform 1 0 118656 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_455
timestamp 1679585382
transform 1 0 119328 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_462
timestamp 1679585382
transform 1 0 120000 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_469
timestamp 1679585382
transform 1 0 120672 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_476
timestamp 1679585382
transform 1 0 121344 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_483
timestamp 1679585382
transform 1 0 122016 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_490
timestamp 1679585382
transform 1 0 122688 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_497
timestamp 1679585382
transform 1 0 123360 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_504
timestamp 1679585382
transform 1 0 124032 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_511
timestamp 1679585382
transform 1 0 124704 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_518
timestamp 1679585382
transform 1 0 125376 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_525
timestamp 1679585382
transform 1 0 126048 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_532
timestamp 1679585382
transform 1 0 126720 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_539
timestamp 1679585382
transform 1 0 127392 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_546
timestamp 1679585382
transform 1 0 128064 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_553
timestamp 1679585382
transform 1 0 128736 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_560
timestamp 1679585382
transform 1 0 129408 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_567
timestamp 1679585382
transform 1 0 130080 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_574
timestamp 1679585382
transform 1 0 130752 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_581
timestamp 1679585382
transform 1 0 131424 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_588
timestamp 1679585382
transform 1 0 132096 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_595
timestamp 1679585382
transform 1 0 132768 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_602
timestamp 1679585382
transform 1 0 133440 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_609
timestamp 1679585382
transform 1 0 134112 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_616
timestamp 1679585382
transform 1 0 134784 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_623
timestamp 1679585382
transform 1 0 135456 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_630
timestamp 1679585382
transform 1 0 136128 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_637
timestamp 1679585382
transform 1 0 136800 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_644
timestamp 1679585382
transform 1 0 137472 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_651
timestamp 1679585382
transform 1 0 138144 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_658
timestamp 1679585382
transform 1 0 138816 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_665
timestamp 1679585382
transform 1 0 139488 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_672
timestamp 1679585382
transform 1 0 140160 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_679
timestamp 1679585382
transform 1 0 140832 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_686
timestamp 1679585382
transform 1 0 141504 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_693
timestamp 1679585382
transform 1 0 142176 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_700
timestamp 1679585382
transform 1 0 142848 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_707
timestamp 1679585382
transform 1 0 143520 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_714
timestamp 1679585382
transform 1 0 144192 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_721
timestamp 1679585382
transform 1 0 144864 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_728
timestamp 1679585382
transform 1 0 145536 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_735
timestamp 1679585382
transform 1 0 146208 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_742
timestamp 1679585382
transform 1 0 146880 0 -1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_3_749
timestamp 1679585382
transform 1 0 147552 0 -1 78624
box -48 -56 720 834
use sg13g2_fill_1  FILLER_3_756
timestamp 1677583258
transform 1 0 148224 0 -1 78624
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_0
timestamp 1679585382
transform 1 0 75648 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_7
timestamp 1679585382
transform 1 0 76320 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_14
timestamp 1679585382
transform 1 0 76992 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_21
timestamp 1679585382
transform 1 0 77664 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_28
timestamp 1679585382
transform 1 0 78336 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_35
timestamp 1679585382
transform 1 0 79008 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_42
timestamp 1679585382
transform 1 0 79680 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_49
timestamp 1679585382
transform 1 0 80352 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_56
timestamp 1679585382
transform 1 0 81024 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_63
timestamp 1679585382
transform 1 0 81696 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_70
timestamp 1679585382
transform 1 0 82368 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_77
timestamp 1679585382
transform 1 0 83040 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_84
timestamp 1679585382
transform 1 0 83712 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_91
timestamp 1679585382
transform 1 0 84384 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_98
timestamp 1679585382
transform 1 0 85056 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_105
timestamp 1679585382
transform 1 0 85728 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_112
timestamp 1679585382
transform 1 0 86400 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_119
timestamp 1679585382
transform 1 0 87072 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_126
timestamp 1679585382
transform 1 0 87744 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_133
timestamp 1679585382
transform 1 0 88416 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_140
timestamp 1679585382
transform 1 0 89088 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_147
timestamp 1679585382
transform 1 0 89760 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_154
timestamp 1679585382
transform 1 0 90432 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_161
timestamp 1679585382
transform 1 0 91104 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_168
timestamp 1679585382
transform 1 0 91776 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_175
timestamp 1679585382
transform 1 0 92448 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_182
timestamp 1679585382
transform 1 0 93120 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_189
timestamp 1679585382
transform 1 0 93792 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_196
timestamp 1679585382
transform 1 0 94464 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_203
timestamp 1679585382
transform 1 0 95136 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_210
timestamp 1679585382
transform 1 0 95808 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_217
timestamp 1679585382
transform 1 0 96480 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_224
timestamp 1679585382
transform 1 0 97152 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_231
timestamp 1679585382
transform 1 0 97824 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_238
timestamp 1679585382
transform 1 0 98496 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_245
timestamp 1679585382
transform 1 0 99168 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_252
timestamp 1679585382
transform 1 0 99840 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_259
timestamp 1679585382
transform 1 0 100512 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_266
timestamp 1679585382
transform 1 0 101184 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_273
timestamp 1679585382
transform 1 0 101856 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_280
timestamp 1679585382
transform 1 0 102528 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_287
timestamp 1679585382
transform 1 0 103200 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_294
timestamp 1679585382
transform 1 0 103872 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_301
timestamp 1679585382
transform 1 0 104544 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_308
timestamp 1679585382
transform 1 0 105216 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_315
timestamp 1679585382
transform 1 0 105888 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_322
timestamp 1679585382
transform 1 0 106560 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_329
timestamp 1679585382
transform 1 0 107232 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_336
timestamp 1679585382
transform 1 0 107904 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_343
timestamp 1679585382
transform 1 0 108576 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_350
timestamp 1679585382
transform 1 0 109248 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_357
timestamp 1679585382
transform 1 0 109920 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_364
timestamp 1679585382
transform 1 0 110592 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_371
timestamp 1679585382
transform 1 0 111264 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_378
timestamp 1679585382
transform 1 0 111936 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_385
timestamp 1679585382
transform 1 0 112608 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_392
timestamp 1679585382
transform 1 0 113280 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_399
timestamp 1679585382
transform 1 0 113952 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_406
timestamp 1679585382
transform 1 0 114624 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_413
timestamp 1679585382
transform 1 0 115296 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_420
timestamp 1679585382
transform 1 0 115968 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_427
timestamp 1679585382
transform 1 0 116640 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_434
timestamp 1679585382
transform 1 0 117312 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_441
timestamp 1679585382
transform 1 0 117984 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_448
timestamp 1679585382
transform 1 0 118656 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_455
timestamp 1679585382
transform 1 0 119328 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_462
timestamp 1679585382
transform 1 0 120000 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_469
timestamp 1679585382
transform 1 0 120672 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_476
timestamp 1679585382
transform 1 0 121344 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_483
timestamp 1679585382
transform 1 0 122016 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_490
timestamp 1679585382
transform 1 0 122688 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_497
timestamp 1679585382
transform 1 0 123360 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_504
timestamp 1679585382
transform 1 0 124032 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_511
timestamp 1679585382
transform 1 0 124704 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_518
timestamp 1679585382
transform 1 0 125376 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_525
timestamp 1679585382
transform 1 0 126048 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_532
timestamp 1679585382
transform 1 0 126720 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_539
timestamp 1679585382
transform 1 0 127392 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_546
timestamp 1679585382
transform 1 0 128064 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_553
timestamp 1679585382
transform 1 0 128736 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_560
timestamp 1679585382
transform 1 0 129408 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_567
timestamp 1679585382
transform 1 0 130080 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_574
timestamp 1679585382
transform 1 0 130752 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_581
timestamp 1679585382
transform 1 0 131424 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_588
timestamp 1679585382
transform 1 0 132096 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_595
timestamp 1679585382
transform 1 0 132768 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_602
timestamp 1679585382
transform 1 0 133440 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_609
timestamp 1679585382
transform 1 0 134112 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_616
timestamp 1679585382
transform 1 0 134784 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_623
timestamp 1679585382
transform 1 0 135456 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_630
timestamp 1679585382
transform 1 0 136128 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_637
timestamp 1679585382
transform 1 0 136800 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_644
timestamp 1679585382
transform 1 0 137472 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_651
timestamp 1679585382
transform 1 0 138144 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_658
timestamp 1679585382
transform 1 0 138816 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_665
timestamp 1679585382
transform 1 0 139488 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_672
timestamp 1679585382
transform 1 0 140160 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_679
timestamp 1679585382
transform 1 0 140832 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_686
timestamp 1679585382
transform 1 0 141504 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_693
timestamp 1679585382
transform 1 0 142176 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_700
timestamp 1679585382
transform 1 0 142848 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_707
timestamp 1679585382
transform 1 0 143520 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_714
timestamp 1679585382
transform 1 0 144192 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_721
timestamp 1679585382
transform 1 0 144864 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_728
timestamp 1679585382
transform 1 0 145536 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_735
timestamp 1679585382
transform 1 0 146208 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_742
timestamp 1679585382
transform 1 0 146880 0 1 78624
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_749
timestamp 1679585382
transform 1 0 147552 0 1 78624
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_756
timestamp 1677583258
transform 1 0 148224 0 1 78624
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_0
timestamp 1679585382
transform 1 0 75648 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_7
timestamp 1679585382
transform 1 0 76320 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_14
timestamp 1679585382
transform 1 0 76992 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_21
timestamp 1679585382
transform 1 0 77664 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_28
timestamp 1679585382
transform 1 0 78336 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_35
timestamp 1679585382
transform 1 0 79008 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_42
timestamp 1679585382
transform 1 0 79680 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_49
timestamp 1679585382
transform 1 0 80352 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_56
timestamp 1679585382
transform 1 0 81024 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_63
timestamp 1679585382
transform 1 0 81696 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_70
timestamp 1679585382
transform 1 0 82368 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_77
timestamp 1679585382
transform 1 0 83040 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_84
timestamp 1679585382
transform 1 0 83712 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_91
timestamp 1679585382
transform 1 0 84384 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_98
timestamp 1679585382
transform 1 0 85056 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_105
timestamp 1679585382
transform 1 0 85728 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_112
timestamp 1679585382
transform 1 0 86400 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_119
timestamp 1679585382
transform 1 0 87072 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_126
timestamp 1679585382
transform 1 0 87744 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_133
timestamp 1679585382
transform 1 0 88416 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_140
timestamp 1679585382
transform 1 0 89088 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_147
timestamp 1679585382
transform 1 0 89760 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_154
timestamp 1679585382
transform 1 0 90432 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_161
timestamp 1679585382
transform 1 0 91104 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_168
timestamp 1679585382
transform 1 0 91776 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_175
timestamp 1679585382
transform 1 0 92448 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_182
timestamp 1679585382
transform 1 0 93120 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_189
timestamp 1679585382
transform 1 0 93792 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_196
timestamp 1679585382
transform 1 0 94464 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_203
timestamp 1679585382
transform 1 0 95136 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_210
timestamp 1679585382
transform 1 0 95808 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_217
timestamp 1679585382
transform 1 0 96480 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_224
timestamp 1679585382
transform 1 0 97152 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_231
timestamp 1679585382
transform 1 0 97824 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_238
timestamp 1679585382
transform 1 0 98496 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_245
timestamp 1679585382
transform 1 0 99168 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_252
timestamp 1679585382
transform 1 0 99840 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_259
timestamp 1679585382
transform 1 0 100512 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_266
timestamp 1679585382
transform 1 0 101184 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_273
timestamp 1679585382
transform 1 0 101856 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_280
timestamp 1679585382
transform 1 0 102528 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_287
timestamp 1679585382
transform 1 0 103200 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_294
timestamp 1679585382
transform 1 0 103872 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_301
timestamp 1679585382
transform 1 0 104544 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_308
timestamp 1679585382
transform 1 0 105216 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_315
timestamp 1679585382
transform 1 0 105888 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_322
timestamp 1679585382
transform 1 0 106560 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_329
timestamp 1679585382
transform 1 0 107232 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_336
timestamp 1679585382
transform 1 0 107904 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_343
timestamp 1679585382
transform 1 0 108576 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_350
timestamp 1679585382
transform 1 0 109248 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_357
timestamp 1679585382
transform 1 0 109920 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_364
timestamp 1679585382
transform 1 0 110592 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_371
timestamp 1679585382
transform 1 0 111264 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_378
timestamp 1679585382
transform 1 0 111936 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_385
timestamp 1679585382
transform 1 0 112608 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_392
timestamp 1679585382
transform 1 0 113280 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_399
timestamp 1679585382
transform 1 0 113952 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_406
timestamp 1679585382
transform 1 0 114624 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_413
timestamp 1679585382
transform 1 0 115296 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_420
timestamp 1679585382
transform 1 0 115968 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_427
timestamp 1679585382
transform 1 0 116640 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_434
timestamp 1679585382
transform 1 0 117312 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_441
timestamp 1679585382
transform 1 0 117984 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_448
timestamp 1679585382
transform 1 0 118656 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_455
timestamp 1679585382
transform 1 0 119328 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_462
timestamp 1679585382
transform 1 0 120000 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_469
timestamp 1679585382
transform 1 0 120672 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_476
timestamp 1679585382
transform 1 0 121344 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_483
timestamp 1679585382
transform 1 0 122016 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_490
timestamp 1679585382
transform 1 0 122688 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_497
timestamp 1679585382
transform 1 0 123360 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_504
timestamp 1679585382
transform 1 0 124032 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_511
timestamp 1679585382
transform 1 0 124704 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_518
timestamp 1679585382
transform 1 0 125376 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_525
timestamp 1679585382
transform 1 0 126048 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_532
timestamp 1679585382
transform 1 0 126720 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_539
timestamp 1679585382
transform 1 0 127392 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_546
timestamp 1679585382
transform 1 0 128064 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_553
timestamp 1679585382
transform 1 0 128736 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_560
timestamp 1679585382
transform 1 0 129408 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_567
timestamp 1679585382
transform 1 0 130080 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_574
timestamp 1679585382
transform 1 0 130752 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_581
timestamp 1679585382
transform 1 0 131424 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_588
timestamp 1679585382
transform 1 0 132096 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_595
timestamp 1679585382
transform 1 0 132768 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_602
timestamp 1679585382
transform 1 0 133440 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_609
timestamp 1679585382
transform 1 0 134112 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_616
timestamp 1679585382
transform 1 0 134784 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_623
timestamp 1679585382
transform 1 0 135456 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_630
timestamp 1679585382
transform 1 0 136128 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_637
timestamp 1679585382
transform 1 0 136800 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_644
timestamp 1679585382
transform 1 0 137472 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_651
timestamp 1679585382
transform 1 0 138144 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_658
timestamp 1679585382
transform 1 0 138816 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_665
timestamp 1679585382
transform 1 0 139488 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_672
timestamp 1679585382
transform 1 0 140160 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_679
timestamp 1679585382
transform 1 0 140832 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_686
timestamp 1679585382
transform 1 0 141504 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_693
timestamp 1679585382
transform 1 0 142176 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_700
timestamp 1679585382
transform 1 0 142848 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_707
timestamp 1679585382
transform 1 0 143520 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_714
timestamp 1679585382
transform 1 0 144192 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_721
timestamp 1679585382
transform 1 0 144864 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_728
timestamp 1679585382
transform 1 0 145536 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_735
timestamp 1679585382
transform 1 0 146208 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_742
timestamp 1679585382
transform 1 0 146880 0 -1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_749
timestamp 1679585382
transform 1 0 147552 0 -1 80136
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_756
timestamp 1677583258
transform 1 0 148224 0 -1 80136
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_0
timestamp 1679585382
transform 1 0 75648 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_7
timestamp 1679585382
transform 1 0 76320 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_14
timestamp 1679585382
transform 1 0 76992 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_21
timestamp 1679585382
transform 1 0 77664 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_28
timestamp 1679585382
transform 1 0 78336 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_35
timestamp 1679585382
transform 1 0 79008 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_42
timestamp 1679585382
transform 1 0 79680 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_49
timestamp 1679585382
transform 1 0 80352 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_56
timestamp 1679585382
transform 1 0 81024 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_63
timestamp 1679585382
transform 1 0 81696 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_70
timestamp 1679585382
transform 1 0 82368 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_77
timestamp 1679585382
transform 1 0 83040 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_84
timestamp 1679585382
transform 1 0 83712 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_91
timestamp 1679585382
transform 1 0 84384 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_98
timestamp 1679585382
transform 1 0 85056 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_105
timestamp 1679585382
transform 1 0 85728 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_112
timestamp 1679585382
transform 1 0 86400 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_119
timestamp 1679585382
transform 1 0 87072 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_126
timestamp 1679585382
transform 1 0 87744 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_133
timestamp 1679585382
transform 1 0 88416 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_140
timestamp 1679585382
transform 1 0 89088 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_147
timestamp 1679585382
transform 1 0 89760 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_154
timestamp 1679585382
transform 1 0 90432 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_161
timestamp 1679585382
transform 1 0 91104 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_168
timestamp 1679585382
transform 1 0 91776 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_175
timestamp 1679585382
transform 1 0 92448 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_182
timestamp 1679585382
transform 1 0 93120 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_189
timestamp 1679585382
transform 1 0 93792 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_196
timestamp 1679585382
transform 1 0 94464 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_203
timestamp 1679585382
transform 1 0 95136 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_210
timestamp 1679585382
transform 1 0 95808 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_217
timestamp 1679585382
transform 1 0 96480 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_224
timestamp 1679585382
transform 1 0 97152 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_231
timestamp 1679585382
transform 1 0 97824 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_238
timestamp 1679585382
transform 1 0 98496 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_245
timestamp 1679585382
transform 1 0 99168 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_252
timestamp 1679585382
transform 1 0 99840 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_259
timestamp 1679585382
transform 1 0 100512 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_266
timestamp 1679585382
transform 1 0 101184 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_273
timestamp 1679585382
transform 1 0 101856 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_280
timestamp 1679585382
transform 1 0 102528 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_287
timestamp 1679585382
transform 1 0 103200 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_294
timestamp 1679585382
transform 1 0 103872 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_301
timestamp 1679585382
transform 1 0 104544 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_308
timestamp 1679585382
transform 1 0 105216 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_315
timestamp 1679585382
transform 1 0 105888 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_322
timestamp 1679585382
transform 1 0 106560 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_329
timestamp 1679585382
transform 1 0 107232 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_336
timestamp 1679585382
transform 1 0 107904 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_343
timestamp 1679585382
transform 1 0 108576 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_350
timestamp 1679585382
transform 1 0 109248 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_357
timestamp 1679585382
transform 1 0 109920 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_364
timestamp 1679585382
transform 1 0 110592 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_371
timestamp 1679585382
transform 1 0 111264 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_378
timestamp 1679585382
transform 1 0 111936 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_385
timestamp 1679585382
transform 1 0 112608 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_392
timestamp 1679585382
transform 1 0 113280 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_399
timestamp 1679585382
transform 1 0 113952 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_406
timestamp 1679585382
transform 1 0 114624 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_413
timestamp 1679585382
transform 1 0 115296 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_420
timestamp 1679585382
transform 1 0 115968 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_427
timestamp 1679585382
transform 1 0 116640 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_434
timestamp 1679585382
transform 1 0 117312 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_441
timestamp 1679585382
transform 1 0 117984 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_448
timestamp 1679585382
transform 1 0 118656 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_455
timestamp 1679585382
transform 1 0 119328 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_462
timestamp 1679585382
transform 1 0 120000 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_469
timestamp 1679585382
transform 1 0 120672 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_476
timestamp 1679585382
transform 1 0 121344 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_483
timestamp 1679585382
transform 1 0 122016 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_490
timestamp 1679585382
transform 1 0 122688 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_497
timestamp 1679585382
transform 1 0 123360 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_504
timestamp 1679585382
transform 1 0 124032 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_511
timestamp 1679585382
transform 1 0 124704 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_518
timestamp 1679585382
transform 1 0 125376 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_525
timestamp 1679585382
transform 1 0 126048 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_532
timestamp 1679585382
transform 1 0 126720 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_539
timestamp 1679585382
transform 1 0 127392 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_546
timestamp 1679585382
transform 1 0 128064 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_553
timestamp 1679585382
transform 1 0 128736 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_560
timestamp 1679585382
transform 1 0 129408 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_567
timestamp 1679585382
transform 1 0 130080 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_574
timestamp 1679585382
transform 1 0 130752 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_581
timestamp 1679585382
transform 1 0 131424 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_588
timestamp 1679585382
transform 1 0 132096 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_595
timestamp 1679585382
transform 1 0 132768 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_602
timestamp 1679585382
transform 1 0 133440 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_609
timestamp 1679585382
transform 1 0 134112 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_616
timestamp 1679585382
transform 1 0 134784 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_623
timestamp 1679585382
transform 1 0 135456 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_630
timestamp 1679585382
transform 1 0 136128 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_637
timestamp 1679585382
transform 1 0 136800 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_644
timestamp 1679585382
transform 1 0 137472 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_651
timestamp 1679585382
transform 1 0 138144 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_658
timestamp 1679585382
transform 1 0 138816 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_665
timestamp 1679585382
transform 1 0 139488 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_672
timestamp 1679585382
transform 1 0 140160 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_679
timestamp 1679585382
transform 1 0 140832 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_686
timestamp 1679585382
transform 1 0 141504 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_693
timestamp 1679585382
transform 1 0 142176 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_700
timestamp 1679585382
transform 1 0 142848 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_707
timestamp 1679585382
transform 1 0 143520 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_714
timestamp 1679585382
transform 1 0 144192 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_721
timestamp 1679585382
transform 1 0 144864 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_728
timestamp 1679585382
transform 1 0 145536 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_735
timestamp 1679585382
transform 1 0 146208 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_742
timestamp 1679585382
transform 1 0 146880 0 1 80136
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_749
timestamp 1679585382
transform 1 0 147552 0 1 80136
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_756
timestamp 1677583258
transform 1 0 148224 0 1 80136
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_0
timestamp 1679585382
transform 1 0 75648 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_7
timestamp 1679585382
transform 1 0 76320 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_14
timestamp 1679585382
transform 1 0 76992 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_21
timestamp 1679585382
transform 1 0 77664 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_28
timestamp 1679585382
transform 1 0 78336 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_35
timestamp 1679585382
transform 1 0 79008 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_42
timestamp 1679585382
transform 1 0 79680 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_49
timestamp 1679585382
transform 1 0 80352 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_56
timestamp 1679585382
transform 1 0 81024 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_63
timestamp 1679585382
transform 1 0 81696 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_70
timestamp 1679585382
transform 1 0 82368 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_77
timestamp 1679585382
transform 1 0 83040 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_84
timestamp 1679585382
transform 1 0 83712 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_91
timestamp 1679585382
transform 1 0 84384 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_98
timestamp 1679585382
transform 1 0 85056 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679585382
transform 1 0 85728 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_112
timestamp 1679585382
transform 1 0 86400 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_119
timestamp 1679585382
transform 1 0 87072 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_126
timestamp 1679585382
transform 1 0 87744 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679585382
transform 1 0 88416 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_140
timestamp 1679585382
transform 1 0 89088 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_147
timestamp 1679585382
transform 1 0 89760 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_154
timestamp 1679585382
transform 1 0 90432 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_161
timestamp 1679585382
transform 1 0 91104 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_168
timestamp 1679585382
transform 1 0 91776 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_175
timestamp 1679585382
transform 1 0 92448 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_182
timestamp 1679585382
transform 1 0 93120 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_189
timestamp 1679585382
transform 1 0 93792 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_196
timestamp 1679585382
transform 1 0 94464 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_203
timestamp 1679585382
transform 1 0 95136 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_210
timestamp 1679585382
transform 1 0 95808 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_217
timestamp 1679585382
transform 1 0 96480 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_224
timestamp 1679585382
transform 1 0 97152 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_231
timestamp 1679585382
transform 1 0 97824 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_238
timestamp 1679585382
transform 1 0 98496 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_245
timestamp 1679585382
transform 1 0 99168 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_252
timestamp 1679585382
transform 1 0 99840 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_259
timestamp 1679585382
transform 1 0 100512 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_266
timestamp 1679585382
transform 1 0 101184 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_273
timestamp 1679585382
transform 1 0 101856 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_280
timestamp 1679585382
transform 1 0 102528 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_287
timestamp 1679585382
transform 1 0 103200 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_294
timestamp 1679585382
transform 1 0 103872 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_301
timestamp 1679585382
transform 1 0 104544 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_308
timestamp 1679585382
transform 1 0 105216 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_315
timestamp 1679585382
transform 1 0 105888 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_322
timestamp 1679585382
transform 1 0 106560 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_329
timestamp 1679585382
transform 1 0 107232 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_336
timestamp 1679585382
transform 1 0 107904 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_343
timestamp 1679585382
transform 1 0 108576 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_350
timestamp 1679585382
transform 1 0 109248 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_357
timestamp 1679585382
transform 1 0 109920 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_364
timestamp 1679585382
transform 1 0 110592 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_371
timestamp 1679585382
transform 1 0 111264 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_378
timestamp 1679585382
transform 1 0 111936 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_385
timestamp 1679585382
transform 1 0 112608 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_392
timestamp 1679585382
transform 1 0 113280 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_399
timestamp 1679585382
transform 1 0 113952 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_406
timestamp 1679585382
transform 1 0 114624 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_413
timestamp 1679585382
transform 1 0 115296 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_420
timestamp 1679585382
transform 1 0 115968 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_427
timestamp 1679585382
transform 1 0 116640 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_434
timestamp 1679585382
transform 1 0 117312 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_441
timestamp 1679585382
transform 1 0 117984 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_448
timestamp 1679585382
transform 1 0 118656 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_455
timestamp 1679585382
transform 1 0 119328 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_462
timestamp 1679585382
transform 1 0 120000 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_469
timestamp 1679585382
transform 1 0 120672 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_476
timestamp 1679585382
transform 1 0 121344 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_483
timestamp 1679585382
transform 1 0 122016 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_490
timestamp 1679585382
transform 1 0 122688 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_497
timestamp 1679585382
transform 1 0 123360 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_504
timestamp 1679585382
transform 1 0 124032 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_511
timestamp 1679585382
transform 1 0 124704 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_518
timestamp 1679585382
transform 1 0 125376 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_525
timestamp 1679585382
transform 1 0 126048 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_532
timestamp 1679585382
transform 1 0 126720 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_539
timestamp 1679585382
transform 1 0 127392 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_546
timestamp 1679585382
transform 1 0 128064 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_553
timestamp 1679585382
transform 1 0 128736 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_560
timestamp 1679585382
transform 1 0 129408 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_567
timestamp 1679585382
transform 1 0 130080 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_574
timestamp 1679585382
transform 1 0 130752 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_581
timestamp 1679585382
transform 1 0 131424 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_588
timestamp 1679585382
transform 1 0 132096 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_595
timestamp 1679585382
transform 1 0 132768 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_602
timestamp 1679585382
transform 1 0 133440 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_609
timestamp 1679585382
transform 1 0 134112 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_616
timestamp 1679585382
transform 1 0 134784 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_623
timestamp 1679585382
transform 1 0 135456 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_630
timestamp 1679585382
transform 1 0 136128 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_637
timestamp 1679585382
transform 1 0 136800 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_644
timestamp 1679585382
transform 1 0 137472 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_651
timestamp 1679585382
transform 1 0 138144 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_658
timestamp 1679585382
transform 1 0 138816 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_665
timestamp 1679585382
transform 1 0 139488 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_672
timestamp 1679585382
transform 1 0 140160 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_679
timestamp 1679585382
transform 1 0 140832 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_686
timestamp 1679585382
transform 1 0 141504 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_693
timestamp 1679585382
transform 1 0 142176 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_700
timestamp 1679585382
transform 1 0 142848 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_707
timestamp 1679585382
transform 1 0 143520 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_714
timestamp 1679585382
transform 1 0 144192 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_721
timestamp 1679585382
transform 1 0 144864 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_728
timestamp 1679585382
transform 1 0 145536 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_735
timestamp 1679585382
transform 1 0 146208 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_742
timestamp 1679585382
transform 1 0 146880 0 -1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_749
timestamp 1679585382
transform 1 0 147552 0 -1 81648
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_756
timestamp 1677583258
transform 1 0 148224 0 -1 81648
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_0
timestamp 1679585382
transform 1 0 75648 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_7
timestamp 1679585382
transform 1 0 76320 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_14
timestamp 1679585382
transform 1 0 76992 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_21
timestamp 1679585382
transform 1 0 77664 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_28
timestamp 1679585382
transform 1 0 78336 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_35
timestamp 1679585382
transform 1 0 79008 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_42
timestamp 1679585382
transform 1 0 79680 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_49
timestamp 1679585382
transform 1 0 80352 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_56
timestamp 1679585382
transform 1 0 81024 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_63
timestamp 1679585382
transform 1 0 81696 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_70
timestamp 1679585382
transform 1 0 82368 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_77
timestamp 1679585382
transform 1 0 83040 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_84
timestamp 1679585382
transform 1 0 83712 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_91
timestamp 1679585382
transform 1 0 84384 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_98
timestamp 1679585382
transform 1 0 85056 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_105
timestamp 1679585382
transform 1 0 85728 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_112
timestamp 1679585382
transform 1 0 86400 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_119
timestamp 1679585382
transform 1 0 87072 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_126
timestamp 1679585382
transform 1 0 87744 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_133
timestamp 1679585382
transform 1 0 88416 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_140
timestamp 1679585382
transform 1 0 89088 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_147
timestamp 1679585382
transform 1 0 89760 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_154
timestamp 1679585382
transform 1 0 90432 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_161
timestamp 1679585382
transform 1 0 91104 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_168
timestamp 1679585382
transform 1 0 91776 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_175
timestamp 1679585382
transform 1 0 92448 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_182
timestamp 1679585382
transform 1 0 93120 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_189
timestamp 1679585382
transform 1 0 93792 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_196
timestamp 1679585382
transform 1 0 94464 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_203
timestamp 1679585382
transform 1 0 95136 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_210
timestamp 1679585382
transform 1 0 95808 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_217
timestamp 1679585382
transform 1 0 96480 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_224
timestamp 1679585382
transform 1 0 97152 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_231
timestamp 1679585382
transform 1 0 97824 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_238
timestamp 1679585382
transform 1 0 98496 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_245
timestamp 1679585382
transform 1 0 99168 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_252
timestamp 1679585382
transform 1 0 99840 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_259
timestamp 1679585382
transform 1 0 100512 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_266
timestamp 1679585382
transform 1 0 101184 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_273
timestamp 1679585382
transform 1 0 101856 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_280
timestamp 1679585382
transform 1 0 102528 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_287
timestamp 1679585382
transform 1 0 103200 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_294
timestamp 1679585382
transform 1 0 103872 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_301
timestamp 1679585382
transform 1 0 104544 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_308
timestamp 1679585382
transform 1 0 105216 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_315
timestamp 1679585382
transform 1 0 105888 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_322
timestamp 1679585382
transform 1 0 106560 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_329
timestamp 1679585382
transform 1 0 107232 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_336
timestamp 1679585382
transform 1 0 107904 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_343
timestamp 1679585382
transform 1 0 108576 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_350
timestamp 1679585382
transform 1 0 109248 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_357
timestamp 1679585382
transform 1 0 109920 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_364
timestamp 1679585382
transform 1 0 110592 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_371
timestamp 1679585382
transform 1 0 111264 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_378
timestamp 1679585382
transform 1 0 111936 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_385
timestamp 1679585382
transform 1 0 112608 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_392
timestamp 1679585382
transform 1 0 113280 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_399
timestamp 1679585382
transform 1 0 113952 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_406
timestamp 1679585382
transform 1 0 114624 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_413
timestamp 1679585382
transform 1 0 115296 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_420
timestamp 1679585382
transform 1 0 115968 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_427
timestamp 1679585382
transform 1 0 116640 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_434
timestamp 1679585382
transform 1 0 117312 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_441
timestamp 1679585382
transform 1 0 117984 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_448
timestamp 1679585382
transform 1 0 118656 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_455
timestamp 1679585382
transform 1 0 119328 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_462
timestamp 1679585382
transform 1 0 120000 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_469
timestamp 1679585382
transform 1 0 120672 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_476
timestamp 1679585382
transform 1 0 121344 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_483
timestamp 1679585382
transform 1 0 122016 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_490
timestamp 1679585382
transform 1 0 122688 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_497
timestamp 1679585382
transform 1 0 123360 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_504
timestamp 1679585382
transform 1 0 124032 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_511
timestamp 1679585382
transform 1 0 124704 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_518
timestamp 1679585382
transform 1 0 125376 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_525
timestamp 1679585382
transform 1 0 126048 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_532
timestamp 1679585382
transform 1 0 126720 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_539
timestamp 1679585382
transform 1 0 127392 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_546
timestamp 1679585382
transform 1 0 128064 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_553
timestamp 1679585382
transform 1 0 128736 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_560
timestamp 1679585382
transform 1 0 129408 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_567
timestamp 1679585382
transform 1 0 130080 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_574
timestamp 1679585382
transform 1 0 130752 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_581
timestamp 1679585382
transform 1 0 131424 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_588
timestamp 1679585382
transform 1 0 132096 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_595
timestamp 1679585382
transform 1 0 132768 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_602
timestamp 1679585382
transform 1 0 133440 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_609
timestamp 1679585382
transform 1 0 134112 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_616
timestamp 1679585382
transform 1 0 134784 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_623
timestamp 1679585382
transform 1 0 135456 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_630
timestamp 1679585382
transform 1 0 136128 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_637
timestamp 1679585382
transform 1 0 136800 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_644
timestamp 1679585382
transform 1 0 137472 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_651
timestamp 1679585382
transform 1 0 138144 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_658
timestamp 1679585382
transform 1 0 138816 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_665
timestamp 1679585382
transform 1 0 139488 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_672
timestamp 1679585382
transform 1 0 140160 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_679
timestamp 1679585382
transform 1 0 140832 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_686
timestamp 1679585382
transform 1 0 141504 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_693
timestamp 1679585382
transform 1 0 142176 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_700
timestamp 1679585382
transform 1 0 142848 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_707
timestamp 1679585382
transform 1 0 143520 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_714
timestamp 1679585382
transform 1 0 144192 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_721
timestamp 1679585382
transform 1 0 144864 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_728
timestamp 1679585382
transform 1 0 145536 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_735
timestamp 1679585382
transform 1 0 146208 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_742
timestamp 1679585382
transform 1 0 146880 0 1 81648
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_749
timestamp 1679585382
transform 1 0 147552 0 1 81648
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_756
timestamp 1677583258
transform 1 0 148224 0 1 81648
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679585382
transform 1 0 75648 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_7
timestamp 1679585382
transform 1 0 76320 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_14
timestamp 1679585382
transform 1 0 76992 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_21
timestamp 1679585382
transform 1 0 77664 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_28
timestamp 1679585382
transform 1 0 78336 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_35
timestamp 1679585382
transform 1 0 79008 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_42
timestamp 1679585382
transform 1 0 79680 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_49
timestamp 1679585382
transform 1 0 80352 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_56
timestamp 1679585382
transform 1 0 81024 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_63
timestamp 1679585382
transform 1 0 81696 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_70
timestamp 1679585382
transform 1 0 82368 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_77
timestamp 1679585382
transform 1 0 83040 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_84
timestamp 1679585382
transform 1 0 83712 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_91
timestamp 1679585382
transform 1 0 84384 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_98
timestamp 1679585382
transform 1 0 85056 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_105
timestamp 1679585382
transform 1 0 85728 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_112
timestamp 1679585382
transform 1 0 86400 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_119
timestamp 1679585382
transform 1 0 87072 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_126
timestamp 1679585382
transform 1 0 87744 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_133
timestamp 1679585382
transform 1 0 88416 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_140
timestamp 1679585382
transform 1 0 89088 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_147
timestamp 1679585382
transform 1 0 89760 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_154
timestamp 1679585382
transform 1 0 90432 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_161
timestamp 1679585382
transform 1 0 91104 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_168
timestamp 1679585382
transform 1 0 91776 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_175
timestamp 1679585382
transform 1 0 92448 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_182
timestamp 1679585382
transform 1 0 93120 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_189
timestamp 1679585382
transform 1 0 93792 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_196
timestamp 1679585382
transform 1 0 94464 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_203
timestamp 1679585382
transform 1 0 95136 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_210
timestamp 1679585382
transform 1 0 95808 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_217
timestamp 1679585382
transform 1 0 96480 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_224
timestamp 1679585382
transform 1 0 97152 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_231
timestamp 1679585382
transform 1 0 97824 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_238
timestamp 1679585382
transform 1 0 98496 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_245
timestamp 1679585382
transform 1 0 99168 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_252
timestamp 1679585382
transform 1 0 99840 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_259
timestamp 1679585382
transform 1 0 100512 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_266
timestamp 1679585382
transform 1 0 101184 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_273
timestamp 1679585382
transform 1 0 101856 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_280
timestamp 1679585382
transform 1 0 102528 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_287
timestamp 1679585382
transform 1 0 103200 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_294
timestamp 1679585382
transform 1 0 103872 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_301
timestamp 1679585382
transform 1 0 104544 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_308
timestamp 1679585382
transform 1 0 105216 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_315
timestamp 1679585382
transform 1 0 105888 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_322
timestamp 1679585382
transform 1 0 106560 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_329
timestamp 1679585382
transform 1 0 107232 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_336
timestamp 1679585382
transform 1 0 107904 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_343
timestamp 1679585382
transform 1 0 108576 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_350
timestamp 1679585382
transform 1 0 109248 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_357
timestamp 1679585382
transform 1 0 109920 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_364
timestamp 1679585382
transform 1 0 110592 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_371
timestamp 1679585382
transform 1 0 111264 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_378
timestamp 1679585382
transform 1 0 111936 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_385
timestamp 1679585382
transform 1 0 112608 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_392
timestamp 1679585382
transform 1 0 113280 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_399
timestamp 1679585382
transform 1 0 113952 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_406
timestamp 1679585382
transform 1 0 114624 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_413
timestamp 1679585382
transform 1 0 115296 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_420
timestamp 1679585382
transform 1 0 115968 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_427
timestamp 1679585382
transform 1 0 116640 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_434
timestamp 1679585382
transform 1 0 117312 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_441
timestamp 1679585382
transform 1 0 117984 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_448
timestamp 1679585382
transform 1 0 118656 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_455
timestamp 1679585382
transform 1 0 119328 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_462
timestamp 1679585382
transform 1 0 120000 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_469
timestamp 1679585382
transform 1 0 120672 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_476
timestamp 1679585382
transform 1 0 121344 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_483
timestamp 1679585382
transform 1 0 122016 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_490
timestamp 1679585382
transform 1 0 122688 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_497
timestamp 1679585382
transform 1 0 123360 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_504
timestamp 1679585382
transform 1 0 124032 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_511
timestamp 1679585382
transform 1 0 124704 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_518
timestamp 1679585382
transform 1 0 125376 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_525
timestamp 1679585382
transform 1 0 126048 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_532
timestamp 1679585382
transform 1 0 126720 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_539
timestamp 1679585382
transform 1 0 127392 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_546
timestamp 1679585382
transform 1 0 128064 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_553
timestamp 1679585382
transform 1 0 128736 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_560
timestamp 1679585382
transform 1 0 129408 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_567
timestamp 1679585382
transform 1 0 130080 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_574
timestamp 1679585382
transform 1 0 130752 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_581
timestamp 1679585382
transform 1 0 131424 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_588
timestamp 1679585382
transform 1 0 132096 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_595
timestamp 1679585382
transform 1 0 132768 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_602
timestamp 1679585382
transform 1 0 133440 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_609
timestamp 1679585382
transform 1 0 134112 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_616
timestamp 1679585382
transform 1 0 134784 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_623
timestamp 1679585382
transform 1 0 135456 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_630
timestamp 1679585382
transform 1 0 136128 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_637
timestamp 1679585382
transform 1 0 136800 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_644
timestamp 1679585382
transform 1 0 137472 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_651
timestamp 1679585382
transform 1 0 138144 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_658
timestamp 1679585382
transform 1 0 138816 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_665
timestamp 1679585382
transform 1 0 139488 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_672
timestamp 1679585382
transform 1 0 140160 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_679
timestamp 1679585382
transform 1 0 140832 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_686
timestamp 1679585382
transform 1 0 141504 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_693
timestamp 1679585382
transform 1 0 142176 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_700
timestamp 1679585382
transform 1 0 142848 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_707
timestamp 1679585382
transform 1 0 143520 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_714
timestamp 1679585382
transform 1 0 144192 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_721
timestamp 1679585382
transform 1 0 144864 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_728
timestamp 1679585382
transform 1 0 145536 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_735
timestamp 1679585382
transform 1 0 146208 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_742
timestamp 1679585382
transform 1 0 146880 0 -1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_9_749
timestamp 1679585382
transform 1 0 147552 0 -1 83160
box -48 -56 720 834
use sg13g2_fill_1  FILLER_9_756
timestamp 1677583258
transform 1 0 148224 0 -1 83160
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_0
timestamp 1679585382
transform 1 0 75648 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_7
timestamp 1679585382
transform 1 0 76320 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_14
timestamp 1679585382
transform 1 0 76992 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_21
timestamp 1679585382
transform 1 0 77664 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_28
timestamp 1679585382
transform 1 0 78336 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_35
timestamp 1679585382
transform 1 0 79008 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_42
timestamp 1679585382
transform 1 0 79680 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_49
timestamp 1679585382
transform 1 0 80352 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_56
timestamp 1679585382
transform 1 0 81024 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_63
timestamp 1679585382
transform 1 0 81696 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_70
timestamp 1679585382
transform 1 0 82368 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_77
timestamp 1679585382
transform 1 0 83040 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_84
timestamp 1679585382
transform 1 0 83712 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_91
timestamp 1679585382
transform 1 0 84384 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_98
timestamp 1679585382
transform 1 0 85056 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_105
timestamp 1679585382
transform 1 0 85728 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_112
timestamp 1679585382
transform 1 0 86400 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_119
timestamp 1679585382
transform 1 0 87072 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_126
timestamp 1679585382
transform 1 0 87744 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_133
timestamp 1679585382
transform 1 0 88416 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_140
timestamp 1679585382
transform 1 0 89088 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_147
timestamp 1679585382
transform 1 0 89760 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_154
timestamp 1679585382
transform 1 0 90432 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_161
timestamp 1679585382
transform 1 0 91104 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_168
timestamp 1679585382
transform 1 0 91776 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_175
timestamp 1679585382
transform 1 0 92448 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_182
timestamp 1679585382
transform 1 0 93120 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_189
timestamp 1679585382
transform 1 0 93792 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_196
timestamp 1679585382
transform 1 0 94464 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_203
timestamp 1679585382
transform 1 0 95136 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_210
timestamp 1679585382
transform 1 0 95808 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_217
timestamp 1679585382
transform 1 0 96480 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_224
timestamp 1679585382
transform 1 0 97152 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_231
timestamp 1679585382
transform 1 0 97824 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_238
timestamp 1679585382
transform 1 0 98496 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_245
timestamp 1679585382
transform 1 0 99168 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_252
timestamp 1679585382
transform 1 0 99840 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_259
timestamp 1679585382
transform 1 0 100512 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_266
timestamp 1679585382
transform 1 0 101184 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_273
timestamp 1679585382
transform 1 0 101856 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_280
timestamp 1679585382
transform 1 0 102528 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_287
timestamp 1679585382
transform 1 0 103200 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_294
timestamp 1679585382
transform 1 0 103872 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_301
timestamp 1679585382
transform 1 0 104544 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_308
timestamp 1679585382
transform 1 0 105216 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_315
timestamp 1679585382
transform 1 0 105888 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_322
timestamp 1679585382
transform 1 0 106560 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_329
timestamp 1679585382
transform 1 0 107232 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_336
timestamp 1679585382
transform 1 0 107904 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_343
timestamp 1679585382
transform 1 0 108576 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_350
timestamp 1679585382
transform 1 0 109248 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_357
timestamp 1679585382
transform 1 0 109920 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_364
timestamp 1679585382
transform 1 0 110592 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_371
timestamp 1679585382
transform 1 0 111264 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_378
timestamp 1679585382
transform 1 0 111936 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_385
timestamp 1679585382
transform 1 0 112608 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_392
timestamp 1679585382
transform 1 0 113280 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_399
timestamp 1679585382
transform 1 0 113952 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_406
timestamp 1679585382
transform 1 0 114624 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_413
timestamp 1679585382
transform 1 0 115296 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_420
timestamp 1679585382
transform 1 0 115968 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_427
timestamp 1679585382
transform 1 0 116640 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_434
timestamp 1679585382
transform 1 0 117312 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_441
timestamp 1679585382
transform 1 0 117984 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_448
timestamp 1679585382
transform 1 0 118656 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_455
timestamp 1679585382
transform 1 0 119328 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_462
timestamp 1679585382
transform 1 0 120000 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_469
timestamp 1679585382
transform 1 0 120672 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_476
timestamp 1679585382
transform 1 0 121344 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_483
timestamp 1679585382
transform 1 0 122016 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_490
timestamp 1679585382
transform 1 0 122688 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_497
timestamp 1679585382
transform 1 0 123360 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_504
timestamp 1679585382
transform 1 0 124032 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_511
timestamp 1679585382
transform 1 0 124704 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_518
timestamp 1679585382
transform 1 0 125376 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_525
timestamp 1679585382
transform 1 0 126048 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_532
timestamp 1679585382
transform 1 0 126720 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_539
timestamp 1679585382
transform 1 0 127392 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_546
timestamp 1679585382
transform 1 0 128064 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_553
timestamp 1679585382
transform 1 0 128736 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_560
timestamp 1679585382
transform 1 0 129408 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_567
timestamp 1679585382
transform 1 0 130080 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_574
timestamp 1679585382
transform 1 0 130752 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_581
timestamp 1679585382
transform 1 0 131424 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_588
timestamp 1679585382
transform 1 0 132096 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_595
timestamp 1679585382
transform 1 0 132768 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_602
timestamp 1679585382
transform 1 0 133440 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_609
timestamp 1679585382
transform 1 0 134112 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_616
timestamp 1679585382
transform 1 0 134784 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_623
timestamp 1679585382
transform 1 0 135456 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_630
timestamp 1679585382
transform 1 0 136128 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_637
timestamp 1679585382
transform 1 0 136800 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_644
timestamp 1679585382
transform 1 0 137472 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_651
timestamp 1679585382
transform 1 0 138144 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_658
timestamp 1679585382
transform 1 0 138816 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_665
timestamp 1679585382
transform 1 0 139488 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_672
timestamp 1679585382
transform 1 0 140160 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_679
timestamp 1679585382
transform 1 0 140832 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_686
timestamp 1679585382
transform 1 0 141504 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_693
timestamp 1679585382
transform 1 0 142176 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_700
timestamp 1679585382
transform 1 0 142848 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_707
timestamp 1679585382
transform 1 0 143520 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_714
timestamp 1679585382
transform 1 0 144192 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_721
timestamp 1679585382
transform 1 0 144864 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_728
timestamp 1679585382
transform 1 0 145536 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_735
timestamp 1679585382
transform 1 0 146208 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_742
timestamp 1679585382
transform 1 0 146880 0 1 83160
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_749
timestamp 1679585382
transform 1 0 147552 0 1 83160
box -48 -56 720 834
use sg13g2_fill_1  FILLER_10_756
timestamp 1677583258
transform 1 0 148224 0 1 83160
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_0
timestamp 1679585382
transform 1 0 75648 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_7
timestamp 1679585382
transform 1 0 76320 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_14
timestamp 1679585382
transform 1 0 76992 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_21
timestamp 1679585382
transform 1 0 77664 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_28
timestamp 1679585382
transform 1 0 78336 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_35
timestamp 1679585382
transform 1 0 79008 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_42
timestamp 1679585382
transform 1 0 79680 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_49
timestamp 1679585382
transform 1 0 80352 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_56
timestamp 1679585382
transform 1 0 81024 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_63
timestamp 1679585382
transform 1 0 81696 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_70
timestamp 1679585382
transform 1 0 82368 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_77
timestamp 1679585382
transform 1 0 83040 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_84
timestamp 1679585382
transform 1 0 83712 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_91
timestamp 1679585382
transform 1 0 84384 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_98
timestamp 1679585382
transform 1 0 85056 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_105
timestamp 1679585382
transform 1 0 85728 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_112
timestamp 1679585382
transform 1 0 86400 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_119
timestamp 1679585382
transform 1 0 87072 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_126
timestamp 1679585382
transform 1 0 87744 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_133
timestamp 1679585382
transform 1 0 88416 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_140
timestamp 1679585382
transform 1 0 89088 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_147
timestamp 1679585382
transform 1 0 89760 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_154
timestamp 1679585382
transform 1 0 90432 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_161
timestamp 1679585382
transform 1 0 91104 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_168
timestamp 1679585382
transform 1 0 91776 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_175
timestamp 1679585382
transform 1 0 92448 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_182
timestamp 1679585382
transform 1 0 93120 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_189
timestamp 1679585382
transform 1 0 93792 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_196
timestamp 1679585382
transform 1 0 94464 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_203
timestamp 1679585382
transform 1 0 95136 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_210
timestamp 1679585382
transform 1 0 95808 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_217
timestamp 1679585382
transform 1 0 96480 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_224
timestamp 1679585382
transform 1 0 97152 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_231
timestamp 1679585382
transform 1 0 97824 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_238
timestamp 1679585382
transform 1 0 98496 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_245
timestamp 1679585382
transform 1 0 99168 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_252
timestamp 1679585382
transform 1 0 99840 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_259
timestamp 1679585382
transform 1 0 100512 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_266
timestamp 1679585382
transform 1 0 101184 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_273
timestamp 1679585382
transform 1 0 101856 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_280
timestamp 1679585382
transform 1 0 102528 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_287
timestamp 1679585382
transform 1 0 103200 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_294
timestamp 1679585382
transform 1 0 103872 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_301
timestamp 1679585382
transform 1 0 104544 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_308
timestamp 1679585382
transform 1 0 105216 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_315
timestamp 1679585382
transform 1 0 105888 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_322
timestamp 1679585382
transform 1 0 106560 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_329
timestamp 1679585382
transform 1 0 107232 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_336
timestamp 1679585382
transform 1 0 107904 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_343
timestamp 1679585382
transform 1 0 108576 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_350
timestamp 1679585382
transform 1 0 109248 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_357
timestamp 1679585382
transform 1 0 109920 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_364
timestamp 1679585382
transform 1 0 110592 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_371
timestamp 1679585382
transform 1 0 111264 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_378
timestamp 1679585382
transform 1 0 111936 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_385
timestamp 1679585382
transform 1 0 112608 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_392
timestamp 1679585382
transform 1 0 113280 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_399
timestamp 1679585382
transform 1 0 113952 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_406
timestamp 1679585382
transform 1 0 114624 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_413
timestamp 1679585382
transform 1 0 115296 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_420
timestamp 1679585382
transform 1 0 115968 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_427
timestamp 1679585382
transform 1 0 116640 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_434
timestamp 1679585382
transform 1 0 117312 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_441
timestamp 1679585382
transform 1 0 117984 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_448
timestamp 1679585382
transform 1 0 118656 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_455
timestamp 1679585382
transform 1 0 119328 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_462
timestamp 1679585382
transform 1 0 120000 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_469
timestamp 1679585382
transform 1 0 120672 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_476
timestamp 1679585382
transform 1 0 121344 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_483
timestamp 1679585382
transform 1 0 122016 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_490
timestamp 1679585382
transform 1 0 122688 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_497
timestamp 1679585382
transform 1 0 123360 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_504
timestamp 1679585382
transform 1 0 124032 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_511
timestamp 1679585382
transform 1 0 124704 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_518
timestamp 1679585382
transform 1 0 125376 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_525
timestamp 1679585382
transform 1 0 126048 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_532
timestamp 1679585382
transform 1 0 126720 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_539
timestamp 1679585382
transform 1 0 127392 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_546
timestamp 1679585382
transform 1 0 128064 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_553
timestamp 1679585382
transform 1 0 128736 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_560
timestamp 1679585382
transform 1 0 129408 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_567
timestamp 1679585382
transform 1 0 130080 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_574
timestamp 1679585382
transform 1 0 130752 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_581
timestamp 1679585382
transform 1 0 131424 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_588
timestamp 1679585382
transform 1 0 132096 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_595
timestamp 1679585382
transform 1 0 132768 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_602
timestamp 1679585382
transform 1 0 133440 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_609
timestamp 1679585382
transform 1 0 134112 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_616
timestamp 1679585382
transform 1 0 134784 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_623
timestamp 1679585382
transform 1 0 135456 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_630
timestamp 1679585382
transform 1 0 136128 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_637
timestamp 1679585382
transform 1 0 136800 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_644
timestamp 1679585382
transform 1 0 137472 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_651
timestamp 1679585382
transform 1 0 138144 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_658
timestamp 1679585382
transform 1 0 138816 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_665
timestamp 1679585382
transform 1 0 139488 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_672
timestamp 1679585382
transform 1 0 140160 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_679
timestamp 1679585382
transform 1 0 140832 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_686
timestamp 1679585382
transform 1 0 141504 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_693
timestamp 1679585382
transform 1 0 142176 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_700
timestamp 1679585382
transform 1 0 142848 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_707
timestamp 1679585382
transform 1 0 143520 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_714
timestamp 1679585382
transform 1 0 144192 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_721
timestamp 1679585382
transform 1 0 144864 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_728
timestamp 1679585382
transform 1 0 145536 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_735
timestamp 1679585382
transform 1 0 146208 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_742
timestamp 1679585382
transform 1 0 146880 0 -1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_749
timestamp 1679585382
transform 1 0 147552 0 -1 84672
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_756
timestamp 1677583258
transform 1 0 148224 0 -1 84672
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_0
timestamp 1679585382
transform 1 0 75648 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_7
timestamp 1679585382
transform 1 0 76320 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_14
timestamp 1679585382
transform 1 0 76992 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_21
timestamp 1679585382
transform 1 0 77664 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_28
timestamp 1679585382
transform 1 0 78336 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_35
timestamp 1679585382
transform 1 0 79008 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_42
timestamp 1679585382
transform 1 0 79680 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_49
timestamp 1679585382
transform 1 0 80352 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_56
timestamp 1679585382
transform 1 0 81024 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_63
timestamp 1679585382
transform 1 0 81696 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_70
timestamp 1679585382
transform 1 0 82368 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_77
timestamp 1679585382
transform 1 0 83040 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_84
timestamp 1679585382
transform 1 0 83712 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_91
timestamp 1679585382
transform 1 0 84384 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_98
timestamp 1679585382
transform 1 0 85056 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_105
timestamp 1679585382
transform 1 0 85728 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_112
timestamp 1679585382
transform 1 0 86400 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_119
timestamp 1679585382
transform 1 0 87072 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_126
timestamp 1679585382
transform 1 0 87744 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_133
timestamp 1679585382
transform 1 0 88416 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_140
timestamp 1679585382
transform 1 0 89088 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_147
timestamp 1679585382
transform 1 0 89760 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_154
timestamp 1679585382
transform 1 0 90432 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_161
timestamp 1679585382
transform 1 0 91104 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_168
timestamp 1679585382
transform 1 0 91776 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_175
timestamp 1679585382
transform 1 0 92448 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_182
timestamp 1679585382
transform 1 0 93120 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_189
timestamp 1679585382
transform 1 0 93792 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_196
timestamp 1679585382
transform 1 0 94464 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_203
timestamp 1679585382
transform 1 0 95136 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_210
timestamp 1679585382
transform 1 0 95808 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_217
timestamp 1679585382
transform 1 0 96480 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_224
timestamp 1679585382
transform 1 0 97152 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_231
timestamp 1679585382
transform 1 0 97824 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_238
timestamp 1679585382
transform 1 0 98496 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_245
timestamp 1679585382
transform 1 0 99168 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_252
timestamp 1679585382
transform 1 0 99840 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_259
timestamp 1679585382
transform 1 0 100512 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_266
timestamp 1679585382
transform 1 0 101184 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_273
timestamp 1679585382
transform 1 0 101856 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_280
timestamp 1679585382
transform 1 0 102528 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_287
timestamp 1679585382
transform 1 0 103200 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_294
timestamp 1679585382
transform 1 0 103872 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_301
timestamp 1679585382
transform 1 0 104544 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_308
timestamp 1679585382
transform 1 0 105216 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_315
timestamp 1679585382
transform 1 0 105888 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_322
timestamp 1679585382
transform 1 0 106560 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_329
timestamp 1679585382
transform 1 0 107232 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_336
timestamp 1679585382
transform 1 0 107904 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_343
timestamp 1679585382
transform 1 0 108576 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_350
timestamp 1679585382
transform 1 0 109248 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_357
timestamp 1679585382
transform 1 0 109920 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_364
timestamp 1679585382
transform 1 0 110592 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_371
timestamp 1679585382
transform 1 0 111264 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_378
timestamp 1679585382
transform 1 0 111936 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_385
timestamp 1679585382
transform 1 0 112608 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_392
timestamp 1679585382
transform 1 0 113280 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_399
timestamp 1679585382
transform 1 0 113952 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_406
timestamp 1679585382
transform 1 0 114624 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_413
timestamp 1679585382
transform 1 0 115296 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_420
timestamp 1679585382
transform 1 0 115968 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_427
timestamp 1679585382
transform 1 0 116640 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_434
timestamp 1679585382
transform 1 0 117312 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_441
timestamp 1679585382
transform 1 0 117984 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_448
timestamp 1679585382
transform 1 0 118656 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_455
timestamp 1679585382
transform 1 0 119328 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_462
timestamp 1679585382
transform 1 0 120000 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_469
timestamp 1679585382
transform 1 0 120672 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_476
timestamp 1679585382
transform 1 0 121344 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_483
timestamp 1679585382
transform 1 0 122016 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_490
timestamp 1679585382
transform 1 0 122688 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_497
timestamp 1679585382
transform 1 0 123360 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_504
timestamp 1679585382
transform 1 0 124032 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_511
timestamp 1679585382
transform 1 0 124704 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_518
timestamp 1679585382
transform 1 0 125376 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_525
timestamp 1679585382
transform 1 0 126048 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_532
timestamp 1679585382
transform 1 0 126720 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_539
timestamp 1679585382
transform 1 0 127392 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_546
timestamp 1679585382
transform 1 0 128064 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_553
timestamp 1679585382
transform 1 0 128736 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_560
timestamp 1679585382
transform 1 0 129408 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_567
timestamp 1679585382
transform 1 0 130080 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_574
timestamp 1679585382
transform 1 0 130752 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_581
timestamp 1679585382
transform 1 0 131424 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_588
timestamp 1679585382
transform 1 0 132096 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_595
timestamp 1679585382
transform 1 0 132768 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_602
timestamp 1679585382
transform 1 0 133440 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_609
timestamp 1679585382
transform 1 0 134112 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_616
timestamp 1679585382
transform 1 0 134784 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_623
timestamp 1679585382
transform 1 0 135456 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_630
timestamp 1679585382
transform 1 0 136128 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_637
timestamp 1679585382
transform 1 0 136800 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_644
timestamp 1679585382
transform 1 0 137472 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_651
timestamp 1679585382
transform 1 0 138144 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_658
timestamp 1679585382
transform 1 0 138816 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_665
timestamp 1679585382
transform 1 0 139488 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_672
timestamp 1679585382
transform 1 0 140160 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_679
timestamp 1679585382
transform 1 0 140832 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_686
timestamp 1679585382
transform 1 0 141504 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_693
timestamp 1679585382
transform 1 0 142176 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_700
timestamp 1679585382
transform 1 0 142848 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_707
timestamp 1679585382
transform 1 0 143520 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_714
timestamp 1679585382
transform 1 0 144192 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_721
timestamp 1679585382
transform 1 0 144864 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_728
timestamp 1679585382
transform 1 0 145536 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_735
timestamp 1679585382
transform 1 0 146208 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_742
timestamp 1679585382
transform 1 0 146880 0 1 84672
box -48 -56 720 834
use sg13g2_decap_8  FILLER_12_749
timestamp 1679585382
transform 1 0 147552 0 1 84672
box -48 -56 720 834
use sg13g2_fill_1  FILLER_12_756
timestamp 1677583258
transform 1 0 148224 0 1 84672
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_0
timestamp 1679585382
transform 1 0 75648 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_7
timestamp 1679585382
transform 1 0 76320 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_14
timestamp 1679585382
transform 1 0 76992 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_21
timestamp 1679585382
transform 1 0 77664 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_28
timestamp 1679585382
transform 1 0 78336 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_35
timestamp 1679585382
transform 1 0 79008 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_42
timestamp 1679585382
transform 1 0 79680 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_49
timestamp 1679585382
transform 1 0 80352 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_56
timestamp 1679585382
transform 1 0 81024 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_63
timestamp 1679585382
transform 1 0 81696 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_70
timestamp 1679585382
transform 1 0 82368 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_77
timestamp 1679585382
transform 1 0 83040 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_84
timestamp 1679585382
transform 1 0 83712 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_91
timestamp 1679585382
transform 1 0 84384 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_98
timestamp 1679585382
transform 1 0 85056 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_105
timestamp 1679585382
transform 1 0 85728 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_112
timestamp 1679585382
transform 1 0 86400 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_119
timestamp 1679585382
transform 1 0 87072 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_126
timestamp 1679585382
transform 1 0 87744 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_133
timestamp 1679585382
transform 1 0 88416 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_140
timestamp 1679585382
transform 1 0 89088 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_147
timestamp 1679585382
transform 1 0 89760 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_154
timestamp 1679585382
transform 1 0 90432 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_161
timestamp 1679585382
transform 1 0 91104 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_168
timestamp 1679585382
transform 1 0 91776 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_175
timestamp 1679585382
transform 1 0 92448 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_182
timestamp 1679585382
transform 1 0 93120 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_189
timestamp 1679585382
transform 1 0 93792 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_196
timestamp 1679585382
transform 1 0 94464 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_203
timestamp 1679585382
transform 1 0 95136 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_210
timestamp 1679585382
transform 1 0 95808 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_217
timestamp 1679585382
transform 1 0 96480 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_224
timestamp 1679585382
transform 1 0 97152 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_231
timestamp 1679585382
transform 1 0 97824 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_238
timestamp 1679585382
transform 1 0 98496 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_245
timestamp 1679585382
transform 1 0 99168 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_252
timestamp 1679585382
transform 1 0 99840 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_259
timestamp 1679585382
transform 1 0 100512 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_266
timestamp 1679585382
transform 1 0 101184 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_273
timestamp 1679585382
transform 1 0 101856 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_280
timestamp 1679585382
transform 1 0 102528 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_287
timestamp 1679585382
transform 1 0 103200 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_294
timestamp 1679585382
transform 1 0 103872 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_301
timestamp 1679585382
transform 1 0 104544 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_308
timestamp 1679585382
transform 1 0 105216 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_315
timestamp 1679585382
transform 1 0 105888 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_322
timestamp 1679585382
transform 1 0 106560 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_329
timestamp 1679585382
transform 1 0 107232 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_336
timestamp 1679585382
transform 1 0 107904 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_343
timestamp 1679585382
transform 1 0 108576 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_350
timestamp 1679585382
transform 1 0 109248 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_357
timestamp 1679585382
transform 1 0 109920 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_364
timestamp 1679585382
transform 1 0 110592 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_371
timestamp 1679585382
transform 1 0 111264 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_378
timestamp 1679585382
transform 1 0 111936 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_385
timestamp 1679585382
transform 1 0 112608 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_392
timestamp 1679585382
transform 1 0 113280 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_399
timestamp 1679585382
transform 1 0 113952 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_406
timestamp 1679585382
transform 1 0 114624 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_413
timestamp 1679585382
transform 1 0 115296 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_420
timestamp 1679585382
transform 1 0 115968 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_427
timestamp 1679585382
transform 1 0 116640 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_434
timestamp 1679585382
transform 1 0 117312 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_441
timestamp 1679585382
transform 1 0 117984 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_448
timestamp 1679585382
transform 1 0 118656 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_455
timestamp 1679585382
transform 1 0 119328 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_462
timestamp 1679585382
transform 1 0 120000 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_469
timestamp 1679585382
transform 1 0 120672 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_476
timestamp 1679585382
transform 1 0 121344 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_483
timestamp 1679585382
transform 1 0 122016 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_490
timestamp 1679585382
transform 1 0 122688 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_497
timestamp 1679585382
transform 1 0 123360 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_504
timestamp 1679585382
transform 1 0 124032 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_511
timestamp 1679585382
transform 1 0 124704 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_518
timestamp 1679585382
transform 1 0 125376 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_525
timestamp 1679585382
transform 1 0 126048 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_532
timestamp 1679585382
transform 1 0 126720 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_539
timestamp 1679585382
transform 1 0 127392 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_546
timestamp 1679585382
transform 1 0 128064 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_553
timestamp 1679585382
transform 1 0 128736 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_560
timestamp 1679585382
transform 1 0 129408 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_567
timestamp 1679585382
transform 1 0 130080 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_574
timestamp 1679585382
transform 1 0 130752 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_581
timestamp 1679585382
transform 1 0 131424 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_588
timestamp 1679585382
transform 1 0 132096 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_595
timestamp 1679585382
transform 1 0 132768 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_602
timestamp 1679585382
transform 1 0 133440 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_609
timestamp 1679585382
transform 1 0 134112 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_616
timestamp 1679585382
transform 1 0 134784 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_623
timestamp 1679585382
transform 1 0 135456 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_630
timestamp 1679585382
transform 1 0 136128 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_637
timestamp 1679585382
transform 1 0 136800 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_644
timestamp 1679585382
transform 1 0 137472 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_651
timestamp 1679585382
transform 1 0 138144 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_658
timestamp 1679585382
transform 1 0 138816 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_665
timestamp 1679585382
transform 1 0 139488 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_672
timestamp 1679585382
transform 1 0 140160 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_679
timestamp 1679585382
transform 1 0 140832 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_686
timestamp 1679585382
transform 1 0 141504 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_693
timestamp 1679585382
transform 1 0 142176 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_700
timestamp 1679585382
transform 1 0 142848 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_707
timestamp 1679585382
transform 1 0 143520 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_714
timestamp 1679585382
transform 1 0 144192 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_721
timestamp 1679585382
transform 1 0 144864 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_728
timestamp 1679585382
transform 1 0 145536 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_735
timestamp 1679585382
transform 1 0 146208 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_742
timestamp 1679585382
transform 1 0 146880 0 -1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_13_749
timestamp 1679585382
transform 1 0 147552 0 -1 86184
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_756
timestamp 1677583258
transform 1 0 148224 0 -1 86184
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_0
timestamp 1679585382
transform 1 0 75648 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_7
timestamp 1679585382
transform 1 0 76320 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_14
timestamp 1679585382
transform 1 0 76992 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_21
timestamp 1679585382
transform 1 0 77664 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_28
timestamp 1679585382
transform 1 0 78336 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_35
timestamp 1679585382
transform 1 0 79008 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_42
timestamp 1679585382
transform 1 0 79680 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_49
timestamp 1679585382
transform 1 0 80352 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_56
timestamp 1679585382
transform 1 0 81024 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_63
timestamp 1679585382
transform 1 0 81696 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_70
timestamp 1679585382
transform 1 0 82368 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_77
timestamp 1679585382
transform 1 0 83040 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_84
timestamp 1679585382
transform 1 0 83712 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_91
timestamp 1679585382
transform 1 0 84384 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_98
timestamp 1679585382
transform 1 0 85056 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_105
timestamp 1679585382
transform 1 0 85728 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_112
timestamp 1679585382
transform 1 0 86400 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_119
timestamp 1679585382
transform 1 0 87072 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_126
timestamp 1679585382
transform 1 0 87744 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_133
timestamp 1679585382
transform 1 0 88416 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_140
timestamp 1679585382
transform 1 0 89088 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_147
timestamp 1679585382
transform 1 0 89760 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_154
timestamp 1679585382
transform 1 0 90432 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_161
timestamp 1679585382
transform 1 0 91104 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_168
timestamp 1679585382
transform 1 0 91776 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_175
timestamp 1679585382
transform 1 0 92448 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_182
timestamp 1679585382
transform 1 0 93120 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_189
timestamp 1679585382
transform 1 0 93792 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_196
timestamp 1679585382
transform 1 0 94464 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_203
timestamp 1679585382
transform 1 0 95136 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_210
timestamp 1679585382
transform 1 0 95808 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_217
timestamp 1679585382
transform 1 0 96480 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_224
timestamp 1679585382
transform 1 0 97152 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_231
timestamp 1679585382
transform 1 0 97824 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_238
timestamp 1679585382
transform 1 0 98496 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_245
timestamp 1679585382
transform 1 0 99168 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_252
timestamp 1679585382
transform 1 0 99840 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_259
timestamp 1679585382
transform 1 0 100512 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_266
timestamp 1679585382
transform 1 0 101184 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_273
timestamp 1679585382
transform 1 0 101856 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_280
timestamp 1679585382
transform 1 0 102528 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_287
timestamp 1679585382
transform 1 0 103200 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_294
timestamp 1679585382
transform 1 0 103872 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_301
timestamp 1679585382
transform 1 0 104544 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_308
timestamp 1679585382
transform 1 0 105216 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_315
timestamp 1679585382
transform 1 0 105888 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_322
timestamp 1679585382
transform 1 0 106560 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_329
timestamp 1679585382
transform 1 0 107232 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_336
timestamp 1679585382
transform 1 0 107904 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_343
timestamp 1679585382
transform 1 0 108576 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_350
timestamp 1679585382
transform 1 0 109248 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_357
timestamp 1679585382
transform 1 0 109920 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_364
timestamp 1679585382
transform 1 0 110592 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_371
timestamp 1679585382
transform 1 0 111264 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_378
timestamp 1679585382
transform 1 0 111936 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_385
timestamp 1679585382
transform 1 0 112608 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_392
timestamp 1679585382
transform 1 0 113280 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_399
timestamp 1679585382
transform 1 0 113952 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_406
timestamp 1679585382
transform 1 0 114624 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_413
timestamp 1679585382
transform 1 0 115296 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_420
timestamp 1679585382
transform 1 0 115968 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_427
timestamp 1679585382
transform 1 0 116640 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_434
timestamp 1679585382
transform 1 0 117312 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_441
timestamp 1679585382
transform 1 0 117984 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_448
timestamp 1679585382
transform 1 0 118656 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_455
timestamp 1679585382
transform 1 0 119328 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_462
timestamp 1679585382
transform 1 0 120000 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_469
timestamp 1679585382
transform 1 0 120672 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_476
timestamp 1679585382
transform 1 0 121344 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_483
timestamp 1679585382
transform 1 0 122016 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_490
timestamp 1679585382
transform 1 0 122688 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_497
timestamp 1679585382
transform 1 0 123360 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_504
timestamp 1679585382
transform 1 0 124032 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_511
timestamp 1679585382
transform 1 0 124704 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_518
timestamp 1679585382
transform 1 0 125376 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_525
timestamp 1679585382
transform 1 0 126048 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_532
timestamp 1679585382
transform 1 0 126720 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_539
timestamp 1679585382
transform 1 0 127392 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_546
timestamp 1679585382
transform 1 0 128064 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_553
timestamp 1679585382
transform 1 0 128736 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_560
timestamp 1679585382
transform 1 0 129408 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_567
timestamp 1679585382
transform 1 0 130080 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_574
timestamp 1679585382
transform 1 0 130752 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_581
timestamp 1679585382
transform 1 0 131424 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_588
timestamp 1679585382
transform 1 0 132096 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_595
timestamp 1679585382
transform 1 0 132768 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_602
timestamp 1679585382
transform 1 0 133440 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_609
timestamp 1679585382
transform 1 0 134112 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_616
timestamp 1679585382
transform 1 0 134784 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_623
timestamp 1679585382
transform 1 0 135456 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_630
timestamp 1679585382
transform 1 0 136128 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_637
timestamp 1679585382
transform 1 0 136800 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_644
timestamp 1679585382
transform 1 0 137472 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_651
timestamp 1679585382
transform 1 0 138144 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_658
timestamp 1679585382
transform 1 0 138816 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_665
timestamp 1679585382
transform 1 0 139488 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_672
timestamp 1679585382
transform 1 0 140160 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_679
timestamp 1679585382
transform 1 0 140832 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_686
timestamp 1679585382
transform 1 0 141504 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_693
timestamp 1679585382
transform 1 0 142176 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_700
timestamp 1679585382
transform 1 0 142848 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_707
timestamp 1679585382
transform 1 0 143520 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_714
timestamp 1679585382
transform 1 0 144192 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_721
timestamp 1679585382
transform 1 0 144864 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_728
timestamp 1679585382
transform 1 0 145536 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_735
timestamp 1679585382
transform 1 0 146208 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_742
timestamp 1679585382
transform 1 0 146880 0 1 86184
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_749
timestamp 1679585382
transform 1 0 147552 0 1 86184
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_756
timestamp 1677583258
transform 1 0 148224 0 1 86184
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_0
timestamp 1679585382
transform 1 0 75648 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_7
timestamp 1679585382
transform 1 0 76320 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_14
timestamp 1679585382
transform 1 0 76992 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_21
timestamp 1679585382
transform 1 0 77664 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_28
timestamp 1679585382
transform 1 0 78336 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_35
timestamp 1679585382
transform 1 0 79008 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_42
timestamp 1679585382
transform 1 0 79680 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_49
timestamp 1679585382
transform 1 0 80352 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_56
timestamp 1679585382
transform 1 0 81024 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_63
timestamp 1679585382
transform 1 0 81696 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_70
timestamp 1679585382
transform 1 0 82368 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_77
timestamp 1679585382
transform 1 0 83040 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_84
timestamp 1679585382
transform 1 0 83712 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_91
timestamp 1679585382
transform 1 0 84384 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_98
timestamp 1679585382
transform 1 0 85056 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_105
timestamp 1679585382
transform 1 0 85728 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_112
timestamp 1679585382
transform 1 0 86400 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_119
timestamp 1679585382
transform 1 0 87072 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_126
timestamp 1679585382
transform 1 0 87744 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_133
timestamp 1679585382
transform 1 0 88416 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_140
timestamp 1679585382
transform 1 0 89088 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_147
timestamp 1679585382
transform 1 0 89760 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_154
timestamp 1679585382
transform 1 0 90432 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_161
timestamp 1679585382
transform 1 0 91104 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_168
timestamp 1679585382
transform 1 0 91776 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_175
timestamp 1679585382
transform 1 0 92448 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_182
timestamp 1679585382
transform 1 0 93120 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_189
timestamp 1679585382
transform 1 0 93792 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_196
timestamp 1679585382
transform 1 0 94464 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_203
timestamp 1679585382
transform 1 0 95136 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_210
timestamp 1679585382
transform 1 0 95808 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_217
timestamp 1679585382
transform 1 0 96480 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_224
timestamp 1679585382
transform 1 0 97152 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_231
timestamp 1679585382
transform 1 0 97824 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_238
timestamp 1679585382
transform 1 0 98496 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_245
timestamp 1679585382
transform 1 0 99168 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_252
timestamp 1679585382
transform 1 0 99840 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_259
timestamp 1679585382
transform 1 0 100512 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_266
timestamp 1679585382
transform 1 0 101184 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_273
timestamp 1679585382
transform 1 0 101856 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_280
timestamp 1679585382
transform 1 0 102528 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_287
timestamp 1679585382
transform 1 0 103200 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_294
timestamp 1679585382
transform 1 0 103872 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_301
timestamp 1679585382
transform 1 0 104544 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_308
timestamp 1679585382
transform 1 0 105216 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_315
timestamp 1679585382
transform 1 0 105888 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_322
timestamp 1679585382
transform 1 0 106560 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_329
timestamp 1679585382
transform 1 0 107232 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_336
timestamp 1679585382
transform 1 0 107904 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_343
timestamp 1679585382
transform 1 0 108576 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_350
timestamp 1679585382
transform 1 0 109248 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_357
timestamp 1679585382
transform 1 0 109920 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_364
timestamp 1679585382
transform 1 0 110592 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_371
timestamp 1679585382
transform 1 0 111264 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_378
timestamp 1679585382
transform 1 0 111936 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_385
timestamp 1679585382
transform 1 0 112608 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_392
timestamp 1679585382
transform 1 0 113280 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_399
timestamp 1679585382
transform 1 0 113952 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_406
timestamp 1679585382
transform 1 0 114624 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_413
timestamp 1679585382
transform 1 0 115296 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_420
timestamp 1679585382
transform 1 0 115968 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_427
timestamp 1679585382
transform 1 0 116640 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_434
timestamp 1679585382
transform 1 0 117312 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_441
timestamp 1679585382
transform 1 0 117984 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_448
timestamp 1679585382
transform 1 0 118656 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_455
timestamp 1679585382
transform 1 0 119328 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_462
timestamp 1679585382
transform 1 0 120000 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_469
timestamp 1679585382
transform 1 0 120672 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_476
timestamp 1679585382
transform 1 0 121344 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_483
timestamp 1679585382
transform 1 0 122016 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_490
timestamp 1679585382
transform 1 0 122688 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_497
timestamp 1679585382
transform 1 0 123360 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_504
timestamp 1679585382
transform 1 0 124032 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_511
timestamp 1679585382
transform 1 0 124704 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_518
timestamp 1679585382
transform 1 0 125376 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_525
timestamp 1679585382
transform 1 0 126048 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_532
timestamp 1679585382
transform 1 0 126720 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_539
timestamp 1679585382
transform 1 0 127392 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_546
timestamp 1679585382
transform 1 0 128064 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_553
timestamp 1679585382
transform 1 0 128736 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_560
timestamp 1679585382
transform 1 0 129408 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_567
timestamp 1679585382
transform 1 0 130080 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_574
timestamp 1679585382
transform 1 0 130752 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_581
timestamp 1679585382
transform 1 0 131424 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_588
timestamp 1679585382
transform 1 0 132096 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_595
timestamp 1679585382
transform 1 0 132768 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_602
timestamp 1679585382
transform 1 0 133440 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_609
timestamp 1679585382
transform 1 0 134112 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_616
timestamp 1679585382
transform 1 0 134784 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_623
timestamp 1679585382
transform 1 0 135456 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_630
timestamp 1679585382
transform 1 0 136128 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_637
timestamp 1679585382
transform 1 0 136800 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_644
timestamp 1679585382
transform 1 0 137472 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_651
timestamp 1679585382
transform 1 0 138144 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_658
timestamp 1679585382
transform 1 0 138816 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_665
timestamp 1679585382
transform 1 0 139488 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_672
timestamp 1679585382
transform 1 0 140160 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_679
timestamp 1679585382
transform 1 0 140832 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_686
timestamp 1679585382
transform 1 0 141504 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_693
timestamp 1679585382
transform 1 0 142176 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_700
timestamp 1679585382
transform 1 0 142848 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_707
timestamp 1679585382
transform 1 0 143520 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_714
timestamp 1679585382
transform 1 0 144192 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_721
timestamp 1679585382
transform 1 0 144864 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_728
timestamp 1679585382
transform 1 0 145536 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_735
timestamp 1679585382
transform 1 0 146208 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_742
timestamp 1679585382
transform 1 0 146880 0 -1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_15_749
timestamp 1679585382
transform 1 0 147552 0 -1 87696
box -48 -56 720 834
use sg13g2_fill_1  FILLER_15_756
timestamp 1677583258
transform 1 0 148224 0 -1 87696
box -48 -56 144 834
use sg13g2_decap_8  FILLER_16_0
timestamp 1679585382
transform 1 0 75648 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_7
timestamp 1679585382
transform 1 0 76320 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_14
timestamp 1679585382
transform 1 0 76992 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_21
timestamp 1679585382
transform 1 0 77664 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_28
timestamp 1679585382
transform 1 0 78336 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_35
timestamp 1679585382
transform 1 0 79008 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_42
timestamp 1679585382
transform 1 0 79680 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_49
timestamp 1679585382
transform 1 0 80352 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_56
timestamp 1679585382
transform 1 0 81024 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_63
timestamp 1679585382
transform 1 0 81696 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_70
timestamp 1679585382
transform 1 0 82368 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_77
timestamp 1679585382
transform 1 0 83040 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_84
timestamp 1679585382
transform 1 0 83712 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_91
timestamp 1679585382
transform 1 0 84384 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_98
timestamp 1679585382
transform 1 0 85056 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_105
timestamp 1679585382
transform 1 0 85728 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_112
timestamp 1679585382
transform 1 0 86400 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_119
timestamp 1679585382
transform 1 0 87072 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_126
timestamp 1679585382
transform 1 0 87744 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_133
timestamp 1679585382
transform 1 0 88416 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_140
timestamp 1679585382
transform 1 0 89088 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_147
timestamp 1679585382
transform 1 0 89760 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_154
timestamp 1679585382
transform 1 0 90432 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_161
timestamp 1679585382
transform 1 0 91104 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_168
timestamp 1679585382
transform 1 0 91776 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_175
timestamp 1679585382
transform 1 0 92448 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_182
timestamp 1679585382
transform 1 0 93120 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_189
timestamp 1679585382
transform 1 0 93792 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_196
timestamp 1679585382
transform 1 0 94464 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_203
timestamp 1679585382
transform 1 0 95136 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_210
timestamp 1679585382
transform 1 0 95808 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_217
timestamp 1679585382
transform 1 0 96480 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_224
timestamp 1679585382
transform 1 0 97152 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_231
timestamp 1679585382
transform 1 0 97824 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_238
timestamp 1679585382
transform 1 0 98496 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_245
timestamp 1679585382
transform 1 0 99168 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_252
timestamp 1679585382
transform 1 0 99840 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_259
timestamp 1679585382
transform 1 0 100512 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_266
timestamp 1679585382
transform 1 0 101184 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_273
timestamp 1679585382
transform 1 0 101856 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_280
timestamp 1679585382
transform 1 0 102528 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_287
timestamp 1679585382
transform 1 0 103200 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_294
timestamp 1679585382
transform 1 0 103872 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_301
timestamp 1679585382
transform 1 0 104544 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_308
timestamp 1679585382
transform 1 0 105216 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_315
timestamp 1679585382
transform 1 0 105888 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_322
timestamp 1679585382
transform 1 0 106560 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_329
timestamp 1679585382
transform 1 0 107232 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_336
timestamp 1679585382
transform 1 0 107904 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_343
timestamp 1679585382
transform 1 0 108576 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_350
timestamp 1679585382
transform 1 0 109248 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_357
timestamp 1679585382
transform 1 0 109920 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_364
timestamp 1679585382
transform 1 0 110592 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_371
timestamp 1679585382
transform 1 0 111264 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_378
timestamp 1679585382
transform 1 0 111936 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_385
timestamp 1679585382
transform 1 0 112608 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_392
timestamp 1679585382
transform 1 0 113280 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_399
timestamp 1679585382
transform 1 0 113952 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_406
timestamp 1679585382
transform 1 0 114624 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_413
timestamp 1679585382
transform 1 0 115296 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_420
timestamp 1679585382
transform 1 0 115968 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_427
timestamp 1679585382
transform 1 0 116640 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_434
timestamp 1679585382
transform 1 0 117312 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_441
timestamp 1679585382
transform 1 0 117984 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_448
timestamp 1679585382
transform 1 0 118656 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_455
timestamp 1679585382
transform 1 0 119328 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_462
timestamp 1679585382
transform 1 0 120000 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_469
timestamp 1679585382
transform 1 0 120672 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_476
timestamp 1679585382
transform 1 0 121344 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_483
timestamp 1679585382
transform 1 0 122016 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_490
timestamp 1679585382
transform 1 0 122688 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_497
timestamp 1679585382
transform 1 0 123360 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_504
timestamp 1679585382
transform 1 0 124032 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_511
timestamp 1679585382
transform 1 0 124704 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_518
timestamp 1679585382
transform 1 0 125376 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_525
timestamp 1679585382
transform 1 0 126048 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_532
timestamp 1679585382
transform 1 0 126720 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_539
timestamp 1679585382
transform 1 0 127392 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_546
timestamp 1679585382
transform 1 0 128064 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_553
timestamp 1679585382
transform 1 0 128736 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_560
timestamp 1679585382
transform 1 0 129408 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_567
timestamp 1679585382
transform 1 0 130080 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_574
timestamp 1679585382
transform 1 0 130752 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_581
timestamp 1679585382
transform 1 0 131424 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_588
timestamp 1679585382
transform 1 0 132096 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_595
timestamp 1679585382
transform 1 0 132768 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_602
timestamp 1679585382
transform 1 0 133440 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_609
timestamp 1679585382
transform 1 0 134112 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_616
timestamp 1679585382
transform 1 0 134784 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_623
timestamp 1679585382
transform 1 0 135456 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_630
timestamp 1679585382
transform 1 0 136128 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_637
timestamp 1679585382
transform 1 0 136800 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_644
timestamp 1679585382
transform 1 0 137472 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_651
timestamp 1679585382
transform 1 0 138144 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_658
timestamp 1679585382
transform 1 0 138816 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_665
timestamp 1679585382
transform 1 0 139488 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_672
timestamp 1679585382
transform 1 0 140160 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_679
timestamp 1679585382
transform 1 0 140832 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_686
timestamp 1679585382
transform 1 0 141504 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_693
timestamp 1679585382
transform 1 0 142176 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_700
timestamp 1679585382
transform 1 0 142848 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_707
timestamp 1679585382
transform 1 0 143520 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_714
timestamp 1679585382
transform 1 0 144192 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_721
timestamp 1679585382
transform 1 0 144864 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_728
timestamp 1679585382
transform 1 0 145536 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_735
timestamp 1679585382
transform 1 0 146208 0 1 87696
box -48 -56 720 834
use sg13g2_decap_8  FILLER_16_742
timestamp 1679585382
transform 1 0 146880 0 1 87696
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_749
timestamp 1679581501
transform 1 0 147552 0 1 87696
box -48 -56 432 834
use sg13g2_decap_8  FILLER_17_0
timestamp 1679585382
transform 1 0 75648 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_7
timestamp 1679585382
transform 1 0 76320 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_14
timestamp 1679585382
transform 1 0 76992 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_21
timestamp 1679585382
transform 1 0 77664 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_28
timestamp 1679585382
transform 1 0 78336 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_35
timestamp 1679585382
transform 1 0 79008 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_42
timestamp 1679585382
transform 1 0 79680 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_49
timestamp 1679585382
transform 1 0 80352 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_56
timestamp 1679585382
transform 1 0 81024 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_63
timestamp 1679585382
transform 1 0 81696 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_70
timestamp 1679585382
transform 1 0 82368 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_77
timestamp 1679585382
transform 1 0 83040 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_84
timestamp 1679585382
transform 1 0 83712 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_91
timestamp 1679585382
transform 1 0 84384 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_98
timestamp 1679585382
transform 1 0 85056 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_105
timestamp 1679585382
transform 1 0 85728 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_112
timestamp 1679585382
transform 1 0 86400 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_119
timestamp 1679585382
transform 1 0 87072 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_126
timestamp 1679585382
transform 1 0 87744 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_133
timestamp 1679585382
transform 1 0 88416 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_140
timestamp 1679585382
transform 1 0 89088 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_147
timestamp 1679585382
transform 1 0 89760 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_154
timestamp 1679585382
transform 1 0 90432 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_161
timestamp 1679585382
transform 1 0 91104 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_168
timestamp 1679585382
transform 1 0 91776 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_175
timestamp 1679585382
transform 1 0 92448 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_182
timestamp 1679585382
transform 1 0 93120 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_189
timestamp 1679585382
transform 1 0 93792 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_196
timestamp 1679585382
transform 1 0 94464 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_203
timestamp 1679585382
transform 1 0 95136 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_210
timestamp 1679585382
transform 1 0 95808 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_217
timestamp 1679585382
transform 1 0 96480 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_224
timestamp 1679585382
transform 1 0 97152 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_231
timestamp 1679585382
transform 1 0 97824 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_238
timestamp 1679585382
transform 1 0 98496 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_245
timestamp 1679585382
transform 1 0 99168 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_252
timestamp 1679585382
transform 1 0 99840 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_259
timestamp 1679585382
transform 1 0 100512 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_266
timestamp 1679585382
transform 1 0 101184 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_273
timestamp 1679585382
transform 1 0 101856 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_280
timestamp 1679585382
transform 1 0 102528 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_287
timestamp 1679585382
transform 1 0 103200 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_294
timestamp 1679585382
transform 1 0 103872 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_301
timestamp 1679585382
transform 1 0 104544 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_308
timestamp 1679585382
transform 1 0 105216 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_315
timestamp 1679585382
transform 1 0 105888 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_322
timestamp 1679585382
transform 1 0 106560 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_329
timestamp 1679585382
transform 1 0 107232 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_336
timestamp 1679585382
transform 1 0 107904 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_343
timestamp 1679585382
transform 1 0 108576 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_350
timestamp 1679585382
transform 1 0 109248 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_357
timestamp 1679585382
transform 1 0 109920 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_364
timestamp 1679585382
transform 1 0 110592 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_371
timestamp 1679585382
transform 1 0 111264 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_378
timestamp 1679585382
transform 1 0 111936 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_385
timestamp 1679585382
transform 1 0 112608 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_392
timestamp 1679585382
transform 1 0 113280 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_399
timestamp 1679585382
transform 1 0 113952 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_406
timestamp 1679585382
transform 1 0 114624 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_413
timestamp 1679585382
transform 1 0 115296 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_420
timestamp 1679585382
transform 1 0 115968 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_427
timestamp 1679585382
transform 1 0 116640 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_434
timestamp 1679585382
transform 1 0 117312 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_441
timestamp 1679585382
transform 1 0 117984 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_448
timestamp 1679585382
transform 1 0 118656 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_455
timestamp 1679585382
transform 1 0 119328 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_462
timestamp 1679585382
transform 1 0 120000 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_469
timestamp 1679585382
transform 1 0 120672 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_476
timestamp 1679585382
transform 1 0 121344 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_483
timestamp 1679585382
transform 1 0 122016 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_490
timestamp 1679585382
transform 1 0 122688 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_497
timestamp 1679585382
transform 1 0 123360 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_504
timestamp 1679585382
transform 1 0 124032 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_511
timestamp 1679585382
transform 1 0 124704 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_518
timestamp 1679585382
transform 1 0 125376 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_525
timestamp 1679585382
transform 1 0 126048 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_532
timestamp 1679585382
transform 1 0 126720 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_539
timestamp 1679585382
transform 1 0 127392 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_546
timestamp 1679585382
transform 1 0 128064 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_553
timestamp 1679585382
transform 1 0 128736 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_560
timestamp 1679585382
transform 1 0 129408 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_567
timestamp 1679585382
transform 1 0 130080 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_574
timestamp 1679585382
transform 1 0 130752 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_581
timestamp 1679585382
transform 1 0 131424 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_588
timestamp 1679585382
transform 1 0 132096 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_595
timestamp 1679585382
transform 1 0 132768 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_602
timestamp 1679585382
transform 1 0 133440 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_609
timestamp 1679585382
transform 1 0 134112 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_616
timestamp 1679585382
transform 1 0 134784 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_623
timestamp 1679585382
transform 1 0 135456 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_630
timestamp 1679585382
transform 1 0 136128 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_637
timestamp 1679585382
transform 1 0 136800 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_644
timestamp 1679585382
transform 1 0 137472 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_651
timestamp 1679585382
transform 1 0 138144 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_658
timestamp 1679585382
transform 1 0 138816 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_665
timestamp 1679585382
transform 1 0 139488 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_672
timestamp 1679585382
transform 1 0 140160 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_679
timestamp 1679585382
transform 1 0 140832 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_686
timestamp 1679585382
transform 1 0 141504 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_693
timestamp 1679585382
transform 1 0 142176 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_700
timestamp 1679585382
transform 1 0 142848 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_707
timestamp 1679585382
transform 1 0 143520 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_714
timestamp 1679585382
transform 1 0 144192 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_721
timestamp 1679585382
transform 1 0 144864 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_728
timestamp 1679585382
transform 1 0 145536 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_735
timestamp 1679585382
transform 1 0 146208 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_742
timestamp 1679585382
transform 1 0 146880 0 -1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_749
timestamp 1679585382
transform 1 0 147552 0 -1 89208
box -48 -56 720 834
use sg13g2_fill_1  FILLER_17_756
timestamp 1677583258
transform 1 0 148224 0 -1 89208
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_0
timestamp 1679585382
transform 1 0 75648 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_7
timestamp 1679585382
transform 1 0 76320 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_14
timestamp 1679585382
transform 1 0 76992 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_21
timestamp 1679585382
transform 1 0 77664 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_28
timestamp 1679585382
transform 1 0 78336 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_35
timestamp 1679585382
transform 1 0 79008 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_42
timestamp 1679585382
transform 1 0 79680 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_49
timestamp 1679585382
transform 1 0 80352 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_56
timestamp 1679585382
transform 1 0 81024 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_63
timestamp 1679585382
transform 1 0 81696 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_70
timestamp 1679585382
transform 1 0 82368 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_77
timestamp 1679585382
transform 1 0 83040 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_84
timestamp 1679585382
transform 1 0 83712 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_91
timestamp 1679585382
transform 1 0 84384 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_98
timestamp 1679585382
transform 1 0 85056 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_105
timestamp 1679585382
transform 1 0 85728 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_112
timestamp 1679585382
transform 1 0 86400 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_119
timestamp 1679585382
transform 1 0 87072 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_126
timestamp 1679585382
transform 1 0 87744 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_133
timestamp 1679585382
transform 1 0 88416 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_140
timestamp 1679585382
transform 1 0 89088 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_147
timestamp 1679585382
transform 1 0 89760 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_154
timestamp 1679585382
transform 1 0 90432 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_161
timestamp 1679585382
transform 1 0 91104 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_168
timestamp 1679585382
transform 1 0 91776 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_175
timestamp 1679585382
transform 1 0 92448 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_182
timestamp 1679585382
transform 1 0 93120 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_189
timestamp 1679585382
transform 1 0 93792 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_196
timestamp 1679585382
transform 1 0 94464 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_203
timestamp 1679585382
transform 1 0 95136 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_210
timestamp 1679585382
transform 1 0 95808 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_217
timestamp 1679585382
transform 1 0 96480 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_224
timestamp 1679585382
transform 1 0 97152 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_231
timestamp 1679585382
transform 1 0 97824 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_238
timestamp 1679585382
transform 1 0 98496 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_245
timestamp 1679585382
transform 1 0 99168 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_252
timestamp 1679585382
transform 1 0 99840 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_259
timestamp 1679585382
transform 1 0 100512 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_266
timestamp 1679585382
transform 1 0 101184 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_273
timestamp 1679585382
transform 1 0 101856 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_280
timestamp 1679585382
transform 1 0 102528 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_287
timestamp 1679585382
transform 1 0 103200 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_294
timestamp 1679585382
transform 1 0 103872 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_301
timestamp 1679585382
transform 1 0 104544 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_308
timestamp 1679585382
transform 1 0 105216 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_315
timestamp 1679585382
transform 1 0 105888 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_322
timestamp 1679585382
transform 1 0 106560 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_329
timestamp 1679585382
transform 1 0 107232 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_336
timestamp 1679585382
transform 1 0 107904 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_343
timestamp 1679585382
transform 1 0 108576 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_350
timestamp 1679585382
transform 1 0 109248 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_357
timestamp 1679585382
transform 1 0 109920 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_364
timestamp 1679585382
transform 1 0 110592 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_371
timestamp 1679585382
transform 1 0 111264 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_378
timestamp 1679585382
transform 1 0 111936 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_385
timestamp 1679585382
transform 1 0 112608 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_392
timestamp 1679585382
transform 1 0 113280 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_399
timestamp 1679585382
transform 1 0 113952 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_406
timestamp 1679585382
transform 1 0 114624 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_413
timestamp 1679585382
transform 1 0 115296 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_420
timestamp 1679585382
transform 1 0 115968 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_427
timestamp 1679585382
transform 1 0 116640 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_434
timestamp 1679585382
transform 1 0 117312 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_441
timestamp 1679585382
transform 1 0 117984 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_448
timestamp 1679585382
transform 1 0 118656 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_455
timestamp 1679585382
transform 1 0 119328 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_462
timestamp 1679585382
transform 1 0 120000 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_469
timestamp 1679585382
transform 1 0 120672 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_476
timestamp 1679585382
transform 1 0 121344 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_483
timestamp 1679585382
transform 1 0 122016 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_490
timestamp 1679585382
transform 1 0 122688 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_497
timestamp 1679585382
transform 1 0 123360 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_504
timestamp 1679585382
transform 1 0 124032 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_511
timestamp 1679585382
transform 1 0 124704 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_518
timestamp 1679585382
transform 1 0 125376 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_525
timestamp 1679585382
transform 1 0 126048 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_532
timestamp 1679585382
transform 1 0 126720 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_539
timestamp 1679585382
transform 1 0 127392 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_546
timestamp 1679585382
transform 1 0 128064 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_553
timestamp 1679585382
transform 1 0 128736 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_560
timestamp 1679585382
transform 1 0 129408 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_567
timestamp 1679585382
transform 1 0 130080 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_574
timestamp 1679585382
transform 1 0 130752 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_581
timestamp 1679585382
transform 1 0 131424 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_588
timestamp 1679585382
transform 1 0 132096 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_595
timestamp 1679585382
transform 1 0 132768 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_602
timestamp 1679585382
transform 1 0 133440 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_609
timestamp 1679585382
transform 1 0 134112 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_616
timestamp 1679585382
transform 1 0 134784 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_623
timestamp 1679585382
transform 1 0 135456 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_630
timestamp 1679585382
transform 1 0 136128 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_637
timestamp 1679585382
transform 1 0 136800 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_644
timestamp 1679585382
transform 1 0 137472 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_651
timestamp 1679585382
transform 1 0 138144 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_658
timestamp 1679585382
transform 1 0 138816 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_665
timestamp 1679585382
transform 1 0 139488 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_672
timestamp 1679585382
transform 1 0 140160 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_679
timestamp 1679585382
transform 1 0 140832 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_686
timestamp 1679585382
transform 1 0 141504 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_693
timestamp 1679585382
transform 1 0 142176 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_700
timestamp 1679585382
transform 1 0 142848 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_707
timestamp 1679585382
transform 1 0 143520 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_714
timestamp 1679585382
transform 1 0 144192 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_721
timestamp 1679585382
transform 1 0 144864 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_728
timestamp 1679585382
transform 1 0 145536 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_735
timestamp 1679585382
transform 1 0 146208 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_742
timestamp 1679585382
transform 1 0 146880 0 1 89208
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_749
timestamp 1679585382
transform 1 0 147552 0 1 89208
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_756
timestamp 1677583258
transform 1 0 148224 0 1 89208
box -48 -56 144 834
use sg13g2_decap_8  FILLER_19_0
timestamp 1679585382
transform 1 0 75648 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_7
timestamp 1679585382
transform 1 0 76320 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_14
timestamp 1679585382
transform 1 0 76992 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_21
timestamp 1679585382
transform 1 0 77664 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_28
timestamp 1679585382
transform 1 0 78336 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_35
timestamp 1679585382
transform 1 0 79008 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_42
timestamp 1679585382
transform 1 0 79680 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_49
timestamp 1679585382
transform 1 0 80352 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_56
timestamp 1679585382
transform 1 0 81024 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_63
timestamp 1679585382
transform 1 0 81696 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_70
timestamp 1679585382
transform 1 0 82368 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_77
timestamp 1679585382
transform 1 0 83040 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_84
timestamp 1679585382
transform 1 0 83712 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_91
timestamp 1679585382
transform 1 0 84384 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_98
timestamp 1679585382
transform 1 0 85056 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_105
timestamp 1679585382
transform 1 0 85728 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_112
timestamp 1679585382
transform 1 0 86400 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_119
timestamp 1679585382
transform 1 0 87072 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_126
timestamp 1679585382
transform 1 0 87744 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_133
timestamp 1679585382
transform 1 0 88416 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_140
timestamp 1679585382
transform 1 0 89088 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_147
timestamp 1679585382
transform 1 0 89760 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_154
timestamp 1679585382
transform 1 0 90432 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_161
timestamp 1679585382
transform 1 0 91104 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_168
timestamp 1679585382
transform 1 0 91776 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_175
timestamp 1679585382
transform 1 0 92448 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_182
timestamp 1679585382
transform 1 0 93120 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_189
timestamp 1679585382
transform 1 0 93792 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_196
timestamp 1679585382
transform 1 0 94464 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_203
timestamp 1679585382
transform 1 0 95136 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_210
timestamp 1679585382
transform 1 0 95808 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_217
timestamp 1679585382
transform 1 0 96480 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_224
timestamp 1679585382
transform 1 0 97152 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_231
timestamp 1679585382
transform 1 0 97824 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_238
timestamp 1679585382
transform 1 0 98496 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_245
timestamp 1679585382
transform 1 0 99168 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_252
timestamp 1679585382
transform 1 0 99840 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_259
timestamp 1679585382
transform 1 0 100512 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_266
timestamp 1679585382
transform 1 0 101184 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_273
timestamp 1679585382
transform 1 0 101856 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_280
timestamp 1679585382
transform 1 0 102528 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_287
timestamp 1679585382
transform 1 0 103200 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_294
timestamp 1679585382
transform 1 0 103872 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_301
timestamp 1679585382
transform 1 0 104544 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_308
timestamp 1679585382
transform 1 0 105216 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_315
timestamp 1679585382
transform 1 0 105888 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_322
timestamp 1679585382
transform 1 0 106560 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_329
timestamp 1679585382
transform 1 0 107232 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_336
timestamp 1679585382
transform 1 0 107904 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_343
timestamp 1679585382
transform 1 0 108576 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_350
timestamp 1679585382
transform 1 0 109248 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_357
timestamp 1679585382
transform 1 0 109920 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_364
timestamp 1679585382
transform 1 0 110592 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_371
timestamp 1679585382
transform 1 0 111264 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_378
timestamp 1679585382
transform 1 0 111936 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_385
timestamp 1679585382
transform 1 0 112608 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_392
timestamp 1679585382
transform 1 0 113280 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_399
timestamp 1679585382
transform 1 0 113952 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_406
timestamp 1679585382
transform 1 0 114624 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_413
timestamp 1679585382
transform 1 0 115296 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_420
timestamp 1679585382
transform 1 0 115968 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_427
timestamp 1679585382
transform 1 0 116640 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_434
timestamp 1679585382
transform 1 0 117312 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_441
timestamp 1679585382
transform 1 0 117984 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_448
timestamp 1679585382
transform 1 0 118656 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_455
timestamp 1679585382
transform 1 0 119328 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_462
timestamp 1679585382
transform 1 0 120000 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_469
timestamp 1679585382
transform 1 0 120672 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_476
timestamp 1679585382
transform 1 0 121344 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_483
timestamp 1679585382
transform 1 0 122016 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_490
timestamp 1679585382
transform 1 0 122688 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_497
timestamp 1679585382
transform 1 0 123360 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_504
timestamp 1679585382
transform 1 0 124032 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_511
timestamp 1679585382
transform 1 0 124704 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_518
timestamp 1679585382
transform 1 0 125376 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_525
timestamp 1679585382
transform 1 0 126048 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_532
timestamp 1679585382
transform 1 0 126720 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_539
timestamp 1679585382
transform 1 0 127392 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_546
timestamp 1679585382
transform 1 0 128064 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_553
timestamp 1679585382
transform 1 0 128736 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_560
timestamp 1679585382
transform 1 0 129408 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_567
timestamp 1679585382
transform 1 0 130080 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_574
timestamp 1679585382
transform 1 0 130752 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_581
timestamp 1679585382
transform 1 0 131424 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_588
timestamp 1679585382
transform 1 0 132096 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_595
timestamp 1679585382
transform 1 0 132768 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_602
timestamp 1679585382
transform 1 0 133440 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_609
timestamp 1679585382
transform 1 0 134112 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_616
timestamp 1679585382
transform 1 0 134784 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_623
timestamp 1679585382
transform 1 0 135456 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_630
timestamp 1679585382
transform 1 0 136128 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_637
timestamp 1679585382
transform 1 0 136800 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_644
timestamp 1679585382
transform 1 0 137472 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_651
timestamp 1679585382
transform 1 0 138144 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_658
timestamp 1679585382
transform 1 0 138816 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_665
timestamp 1679585382
transform 1 0 139488 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_672
timestamp 1679585382
transform 1 0 140160 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_679
timestamp 1679585382
transform 1 0 140832 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_686
timestamp 1679585382
transform 1 0 141504 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_693
timestamp 1679585382
transform 1 0 142176 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_700
timestamp 1679585382
transform 1 0 142848 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_707
timestamp 1679585382
transform 1 0 143520 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_714
timestamp 1679585382
transform 1 0 144192 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_721
timestamp 1679585382
transform 1 0 144864 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_728
timestamp 1679585382
transform 1 0 145536 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_735
timestamp 1679585382
transform 1 0 146208 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_742
timestamp 1679585382
transform 1 0 146880 0 -1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_19_749
timestamp 1679585382
transform 1 0 147552 0 -1 90720
box -48 -56 720 834
use sg13g2_fill_1  FILLER_19_756
timestamp 1677583258
transform 1 0 148224 0 -1 90720
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_0
timestamp 1679585382
transform 1 0 75648 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_7
timestamp 1679585382
transform 1 0 76320 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_14
timestamp 1679585382
transform 1 0 76992 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_21
timestamp 1679585382
transform 1 0 77664 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_28
timestamp 1679585382
transform 1 0 78336 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_35
timestamp 1679585382
transform 1 0 79008 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_42
timestamp 1679585382
transform 1 0 79680 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_49
timestamp 1679585382
transform 1 0 80352 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_56
timestamp 1679585382
transform 1 0 81024 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_63
timestamp 1679585382
transform 1 0 81696 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_70
timestamp 1679585382
transform 1 0 82368 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_77
timestamp 1679585382
transform 1 0 83040 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_84
timestamp 1679585382
transform 1 0 83712 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_91
timestamp 1679585382
transform 1 0 84384 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_98
timestamp 1679585382
transform 1 0 85056 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_105
timestamp 1679585382
transform 1 0 85728 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_112
timestamp 1679585382
transform 1 0 86400 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_119
timestamp 1679585382
transform 1 0 87072 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_126
timestamp 1679585382
transform 1 0 87744 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_133
timestamp 1679585382
transform 1 0 88416 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_140
timestamp 1679585382
transform 1 0 89088 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_147
timestamp 1679585382
transform 1 0 89760 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_154
timestamp 1679585382
transform 1 0 90432 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_161
timestamp 1679585382
transform 1 0 91104 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_168
timestamp 1679585382
transform 1 0 91776 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_175
timestamp 1679585382
transform 1 0 92448 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_182
timestamp 1679585382
transform 1 0 93120 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_189
timestamp 1679585382
transform 1 0 93792 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_196
timestamp 1679585382
transform 1 0 94464 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_203
timestamp 1679585382
transform 1 0 95136 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_210
timestamp 1679585382
transform 1 0 95808 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_217
timestamp 1679585382
transform 1 0 96480 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_224
timestamp 1679585382
transform 1 0 97152 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_231
timestamp 1679585382
transform 1 0 97824 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_238
timestamp 1679585382
transform 1 0 98496 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_245
timestamp 1679585382
transform 1 0 99168 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_252
timestamp 1679585382
transform 1 0 99840 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_259
timestamp 1679585382
transform 1 0 100512 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_266
timestamp 1679585382
transform 1 0 101184 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_273
timestamp 1679585382
transform 1 0 101856 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_280
timestamp 1679585382
transform 1 0 102528 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_287
timestamp 1679585382
transform 1 0 103200 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_294
timestamp 1679585382
transform 1 0 103872 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_301
timestamp 1679585382
transform 1 0 104544 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_308
timestamp 1679585382
transform 1 0 105216 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_315
timestamp 1679585382
transform 1 0 105888 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_322
timestamp 1679585382
transform 1 0 106560 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_329
timestamp 1679585382
transform 1 0 107232 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_336
timestamp 1679585382
transform 1 0 107904 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_343
timestamp 1679585382
transform 1 0 108576 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_350
timestamp 1679585382
transform 1 0 109248 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_357
timestamp 1679585382
transform 1 0 109920 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_364
timestamp 1679585382
transform 1 0 110592 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_371
timestamp 1679585382
transform 1 0 111264 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_378
timestamp 1679585382
transform 1 0 111936 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_385
timestamp 1679585382
transform 1 0 112608 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_392
timestamp 1679585382
transform 1 0 113280 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_399
timestamp 1679585382
transform 1 0 113952 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_406
timestamp 1679585382
transform 1 0 114624 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_413
timestamp 1679585382
transform 1 0 115296 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_420
timestamp 1679585382
transform 1 0 115968 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_427
timestamp 1679585382
transform 1 0 116640 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_434
timestamp 1679585382
transform 1 0 117312 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_441
timestamp 1679585382
transform 1 0 117984 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_448
timestamp 1679585382
transform 1 0 118656 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_455
timestamp 1679585382
transform 1 0 119328 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_462
timestamp 1679585382
transform 1 0 120000 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_469
timestamp 1679585382
transform 1 0 120672 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_476
timestamp 1679585382
transform 1 0 121344 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_483
timestamp 1679585382
transform 1 0 122016 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_490
timestamp 1679585382
transform 1 0 122688 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_497
timestamp 1679585382
transform 1 0 123360 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_504
timestamp 1679585382
transform 1 0 124032 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_511
timestamp 1679585382
transform 1 0 124704 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_518
timestamp 1679585382
transform 1 0 125376 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_525
timestamp 1679585382
transform 1 0 126048 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_532
timestamp 1679585382
transform 1 0 126720 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_539
timestamp 1679585382
transform 1 0 127392 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_546
timestamp 1679585382
transform 1 0 128064 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_553
timestamp 1679585382
transform 1 0 128736 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_560
timestamp 1679585382
transform 1 0 129408 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_567
timestamp 1679585382
transform 1 0 130080 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_574
timestamp 1679585382
transform 1 0 130752 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_581
timestamp 1679585382
transform 1 0 131424 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_588
timestamp 1679585382
transform 1 0 132096 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_595
timestamp 1679585382
transform 1 0 132768 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_602
timestamp 1679585382
transform 1 0 133440 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_609
timestamp 1679585382
transform 1 0 134112 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_616
timestamp 1679585382
transform 1 0 134784 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_623
timestamp 1679585382
transform 1 0 135456 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_630
timestamp 1679585382
transform 1 0 136128 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_637
timestamp 1679585382
transform 1 0 136800 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_644
timestamp 1679585382
transform 1 0 137472 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_651
timestamp 1679585382
transform 1 0 138144 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_658
timestamp 1679585382
transform 1 0 138816 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_665
timestamp 1679585382
transform 1 0 139488 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_672
timestamp 1679585382
transform 1 0 140160 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_679
timestamp 1679585382
transform 1 0 140832 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_686
timestamp 1679585382
transform 1 0 141504 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_693
timestamp 1679585382
transform 1 0 142176 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_700
timestamp 1679585382
transform 1 0 142848 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_707
timestamp 1679585382
transform 1 0 143520 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_714
timestamp 1679585382
transform 1 0 144192 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_721
timestamp 1679585382
transform 1 0 144864 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_728
timestamp 1679585382
transform 1 0 145536 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_735
timestamp 1679585382
transform 1 0 146208 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_742
timestamp 1679585382
transform 1 0 146880 0 1 90720
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_749
timestamp 1679585382
transform 1 0 147552 0 1 90720
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_756
timestamp 1677583258
transform 1 0 148224 0 1 90720
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_0
timestamp 1679585382
transform 1 0 75648 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_7
timestamp 1679585382
transform 1 0 76320 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_14
timestamp 1679585382
transform 1 0 76992 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_21
timestamp 1679585382
transform 1 0 77664 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_28
timestamp 1679585382
transform 1 0 78336 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_35
timestamp 1679585382
transform 1 0 79008 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_42
timestamp 1679585382
transform 1 0 79680 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_49
timestamp 1679585382
transform 1 0 80352 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_56
timestamp 1679585382
transform 1 0 81024 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_63
timestamp 1679585382
transform 1 0 81696 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_70
timestamp 1679585382
transform 1 0 82368 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_77
timestamp 1679585382
transform 1 0 83040 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_84
timestamp 1679585382
transform 1 0 83712 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_91
timestamp 1679585382
transform 1 0 84384 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_98
timestamp 1679585382
transform 1 0 85056 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_105
timestamp 1679585382
transform 1 0 85728 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_112
timestamp 1679585382
transform 1 0 86400 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_119
timestamp 1679585382
transform 1 0 87072 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_126
timestamp 1679585382
transform 1 0 87744 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_133
timestamp 1679585382
transform 1 0 88416 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_140
timestamp 1679585382
transform 1 0 89088 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_147
timestamp 1679585382
transform 1 0 89760 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_154
timestamp 1679585382
transform 1 0 90432 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_161
timestamp 1679585382
transform 1 0 91104 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_168
timestamp 1679585382
transform 1 0 91776 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_175
timestamp 1679585382
transform 1 0 92448 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_182
timestamp 1679585382
transform 1 0 93120 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_189
timestamp 1679585382
transform 1 0 93792 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_196
timestamp 1679585382
transform 1 0 94464 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_203
timestamp 1679585382
transform 1 0 95136 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_210
timestamp 1679585382
transform 1 0 95808 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_217
timestamp 1679585382
transform 1 0 96480 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_224
timestamp 1679585382
transform 1 0 97152 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_231
timestamp 1679585382
transform 1 0 97824 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_238
timestamp 1679585382
transform 1 0 98496 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_245
timestamp 1679585382
transform 1 0 99168 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_252
timestamp 1679585382
transform 1 0 99840 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_259
timestamp 1679585382
transform 1 0 100512 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_266
timestamp 1679585382
transform 1 0 101184 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_273
timestamp 1679585382
transform 1 0 101856 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_280
timestamp 1679585382
transform 1 0 102528 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_287
timestamp 1679585382
transform 1 0 103200 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_294
timestamp 1679585382
transform 1 0 103872 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_301
timestamp 1679585382
transform 1 0 104544 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_308
timestamp 1679585382
transform 1 0 105216 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_315
timestamp 1679585382
transform 1 0 105888 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_322
timestamp 1679585382
transform 1 0 106560 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_329
timestamp 1679585382
transform 1 0 107232 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_336
timestamp 1679585382
transform 1 0 107904 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_343
timestamp 1679585382
transform 1 0 108576 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_350
timestamp 1679585382
transform 1 0 109248 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_357
timestamp 1679585382
transform 1 0 109920 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_364
timestamp 1679585382
transform 1 0 110592 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_371
timestamp 1679585382
transform 1 0 111264 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_378
timestamp 1679585382
transform 1 0 111936 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_385
timestamp 1679585382
transform 1 0 112608 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_392
timestamp 1679585382
transform 1 0 113280 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_399
timestamp 1679585382
transform 1 0 113952 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_406
timestamp 1679585382
transform 1 0 114624 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_413
timestamp 1679585382
transform 1 0 115296 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_420
timestamp 1679585382
transform 1 0 115968 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_427
timestamp 1679585382
transform 1 0 116640 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_434
timestamp 1679585382
transform 1 0 117312 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_441
timestamp 1679585382
transform 1 0 117984 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_448
timestamp 1679585382
transform 1 0 118656 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_455
timestamp 1679585382
transform 1 0 119328 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_462
timestamp 1679585382
transform 1 0 120000 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_469
timestamp 1679585382
transform 1 0 120672 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_476
timestamp 1679585382
transform 1 0 121344 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_483
timestamp 1679585382
transform 1 0 122016 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_490
timestamp 1679585382
transform 1 0 122688 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_497
timestamp 1679585382
transform 1 0 123360 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_504
timestamp 1679585382
transform 1 0 124032 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_511
timestamp 1679585382
transform 1 0 124704 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_518
timestamp 1679585382
transform 1 0 125376 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_525
timestamp 1679585382
transform 1 0 126048 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_532
timestamp 1679585382
transform 1 0 126720 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_539
timestamp 1679585382
transform 1 0 127392 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_546
timestamp 1679585382
transform 1 0 128064 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_553
timestamp 1679585382
transform 1 0 128736 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_560
timestamp 1679585382
transform 1 0 129408 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_567
timestamp 1679585382
transform 1 0 130080 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_574
timestamp 1679585382
transform 1 0 130752 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_581
timestamp 1679585382
transform 1 0 131424 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_588
timestamp 1679585382
transform 1 0 132096 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_595
timestamp 1679585382
transform 1 0 132768 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_602
timestamp 1679585382
transform 1 0 133440 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_609
timestamp 1679585382
transform 1 0 134112 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_616
timestamp 1679585382
transform 1 0 134784 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_623
timestamp 1679585382
transform 1 0 135456 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_630
timestamp 1679585382
transform 1 0 136128 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_637
timestamp 1679585382
transform 1 0 136800 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_644
timestamp 1679585382
transform 1 0 137472 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_651
timestamp 1679585382
transform 1 0 138144 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_658
timestamp 1679585382
transform 1 0 138816 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_665
timestamp 1679585382
transform 1 0 139488 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_672
timestamp 1679585382
transform 1 0 140160 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_679
timestamp 1679585382
transform 1 0 140832 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_686
timestamp 1679585382
transform 1 0 141504 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_693
timestamp 1679585382
transform 1 0 142176 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_700
timestamp 1679585382
transform 1 0 142848 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_707
timestamp 1679585382
transform 1 0 143520 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_714
timestamp 1679585382
transform 1 0 144192 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_721
timestamp 1679585382
transform 1 0 144864 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_728
timestamp 1679585382
transform 1 0 145536 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_735
timestamp 1679585382
transform 1 0 146208 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_742
timestamp 1679585382
transform 1 0 146880 0 -1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_749
timestamp 1679585382
transform 1 0 147552 0 -1 92232
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_756
timestamp 1677583258
transform 1 0 148224 0 -1 92232
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_0
timestamp 1679585382
transform 1 0 75648 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_7
timestamp 1679585382
transform 1 0 76320 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_14
timestamp 1679585382
transform 1 0 76992 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_21
timestamp 1679585382
transform 1 0 77664 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_28
timestamp 1679585382
transform 1 0 78336 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_35
timestamp 1679585382
transform 1 0 79008 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_42
timestamp 1679585382
transform 1 0 79680 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_49
timestamp 1679585382
transform 1 0 80352 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_56
timestamp 1679585382
transform 1 0 81024 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_63
timestamp 1679585382
transform 1 0 81696 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_70
timestamp 1679585382
transform 1 0 82368 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_77
timestamp 1679585382
transform 1 0 83040 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_84
timestamp 1679585382
transform 1 0 83712 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_91
timestamp 1679585382
transform 1 0 84384 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_98
timestamp 1679585382
transform 1 0 85056 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_105
timestamp 1679585382
transform 1 0 85728 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_112
timestamp 1679585382
transform 1 0 86400 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_119
timestamp 1679585382
transform 1 0 87072 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_126
timestamp 1679585382
transform 1 0 87744 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_133
timestamp 1679585382
transform 1 0 88416 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_140
timestamp 1679585382
transform 1 0 89088 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_147
timestamp 1679585382
transform 1 0 89760 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_154
timestamp 1679585382
transform 1 0 90432 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_161
timestamp 1679585382
transform 1 0 91104 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_168
timestamp 1679585382
transform 1 0 91776 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_175
timestamp 1679585382
transform 1 0 92448 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_182
timestamp 1679585382
transform 1 0 93120 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_189
timestamp 1679585382
transform 1 0 93792 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_196
timestamp 1679585382
transform 1 0 94464 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_203
timestamp 1679585382
transform 1 0 95136 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_210
timestamp 1679585382
transform 1 0 95808 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_217
timestamp 1679585382
transform 1 0 96480 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_224
timestamp 1679585382
transform 1 0 97152 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_231
timestamp 1679585382
transform 1 0 97824 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_238
timestamp 1679585382
transform 1 0 98496 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_245
timestamp 1679585382
transform 1 0 99168 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_252
timestamp 1679585382
transform 1 0 99840 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_259
timestamp 1679585382
transform 1 0 100512 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_266
timestamp 1679585382
transform 1 0 101184 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_273
timestamp 1679585382
transform 1 0 101856 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_280
timestamp 1679585382
transform 1 0 102528 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_287
timestamp 1679585382
transform 1 0 103200 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_294
timestamp 1679585382
transform 1 0 103872 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_301
timestamp 1679585382
transform 1 0 104544 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_308
timestamp 1679585382
transform 1 0 105216 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_315
timestamp 1679585382
transform 1 0 105888 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_322
timestamp 1679585382
transform 1 0 106560 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_329
timestamp 1679585382
transform 1 0 107232 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_336
timestamp 1679585382
transform 1 0 107904 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_343
timestamp 1679585382
transform 1 0 108576 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_350
timestamp 1679585382
transform 1 0 109248 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_357
timestamp 1679585382
transform 1 0 109920 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_364
timestamp 1679585382
transform 1 0 110592 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_371
timestamp 1679585382
transform 1 0 111264 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_378
timestamp 1679585382
transform 1 0 111936 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_385
timestamp 1679585382
transform 1 0 112608 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_392
timestamp 1679585382
transform 1 0 113280 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_399
timestamp 1679585382
transform 1 0 113952 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_406
timestamp 1679585382
transform 1 0 114624 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_413
timestamp 1679585382
transform 1 0 115296 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_420
timestamp 1679585382
transform 1 0 115968 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_427
timestamp 1679585382
transform 1 0 116640 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_434
timestamp 1679585382
transform 1 0 117312 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_441
timestamp 1679585382
transform 1 0 117984 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_448
timestamp 1679585382
transform 1 0 118656 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_455
timestamp 1679585382
transform 1 0 119328 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_462
timestamp 1679585382
transform 1 0 120000 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_469
timestamp 1679585382
transform 1 0 120672 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_476
timestamp 1679585382
transform 1 0 121344 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_483
timestamp 1679585382
transform 1 0 122016 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_490
timestamp 1679585382
transform 1 0 122688 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_497
timestamp 1679585382
transform 1 0 123360 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_504
timestamp 1679585382
transform 1 0 124032 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_511
timestamp 1679585382
transform 1 0 124704 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_518
timestamp 1679585382
transform 1 0 125376 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_525
timestamp 1679585382
transform 1 0 126048 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_532
timestamp 1679585382
transform 1 0 126720 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_539
timestamp 1679585382
transform 1 0 127392 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_546
timestamp 1679585382
transform 1 0 128064 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_553
timestamp 1679585382
transform 1 0 128736 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_560
timestamp 1679585382
transform 1 0 129408 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_567
timestamp 1679585382
transform 1 0 130080 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_574
timestamp 1679585382
transform 1 0 130752 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_581
timestamp 1679585382
transform 1 0 131424 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_588
timestamp 1679585382
transform 1 0 132096 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_595
timestamp 1679585382
transform 1 0 132768 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_602
timestamp 1679585382
transform 1 0 133440 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_609
timestamp 1679585382
transform 1 0 134112 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_616
timestamp 1679585382
transform 1 0 134784 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_623
timestamp 1679585382
transform 1 0 135456 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_630
timestamp 1679585382
transform 1 0 136128 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_637
timestamp 1679585382
transform 1 0 136800 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_644
timestamp 1679585382
transform 1 0 137472 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_651
timestamp 1679585382
transform 1 0 138144 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_658
timestamp 1679585382
transform 1 0 138816 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_665
timestamp 1679585382
transform 1 0 139488 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_672
timestamp 1679585382
transform 1 0 140160 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_679
timestamp 1679585382
transform 1 0 140832 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_686
timestamp 1679585382
transform 1 0 141504 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_693
timestamp 1679585382
transform 1 0 142176 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_700
timestamp 1679585382
transform 1 0 142848 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_707
timestamp 1679585382
transform 1 0 143520 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_714
timestamp 1679585382
transform 1 0 144192 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_721
timestamp 1679585382
transform 1 0 144864 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_728
timestamp 1679585382
transform 1 0 145536 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_735
timestamp 1679585382
transform 1 0 146208 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_742
timestamp 1679585382
transform 1 0 146880 0 1 92232
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_749
timestamp 1679585382
transform 1 0 147552 0 1 92232
box -48 -56 720 834
use sg13g2_fill_1  FILLER_22_756
timestamp 1677583258
transform 1 0 148224 0 1 92232
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_0
timestamp 1679585382
transform 1 0 75648 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_7
timestamp 1679585382
transform 1 0 76320 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_14
timestamp 1679585382
transform 1 0 76992 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_21
timestamp 1679585382
transform 1 0 77664 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_28
timestamp 1679585382
transform 1 0 78336 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_35
timestamp 1679585382
transform 1 0 79008 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_42
timestamp 1679585382
transform 1 0 79680 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_49
timestamp 1679585382
transform 1 0 80352 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_56
timestamp 1679585382
transform 1 0 81024 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_63
timestamp 1679585382
transform 1 0 81696 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_70
timestamp 1679585382
transform 1 0 82368 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_77
timestamp 1679585382
transform 1 0 83040 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_84
timestamp 1679585382
transform 1 0 83712 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_91
timestamp 1679585382
transform 1 0 84384 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_98
timestamp 1679585382
transform 1 0 85056 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_105
timestamp 1679585382
transform 1 0 85728 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_112
timestamp 1679585382
transform 1 0 86400 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_119
timestamp 1679585382
transform 1 0 87072 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_126
timestamp 1679585382
transform 1 0 87744 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_133
timestamp 1679585382
transform 1 0 88416 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_140
timestamp 1679585382
transform 1 0 89088 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_147
timestamp 1679585382
transform 1 0 89760 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_154
timestamp 1679585382
transform 1 0 90432 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_161
timestamp 1679585382
transform 1 0 91104 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_168
timestamp 1679585382
transform 1 0 91776 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_175
timestamp 1679585382
transform 1 0 92448 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_182
timestamp 1679585382
transform 1 0 93120 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_189
timestamp 1679585382
transform 1 0 93792 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_196
timestamp 1679585382
transform 1 0 94464 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_203
timestamp 1679585382
transform 1 0 95136 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_210
timestamp 1679585382
transform 1 0 95808 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_217
timestamp 1679585382
transform 1 0 96480 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_224
timestamp 1679585382
transform 1 0 97152 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_231
timestamp 1679585382
transform 1 0 97824 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_238
timestamp 1679585382
transform 1 0 98496 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_245
timestamp 1679585382
transform 1 0 99168 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_252
timestamp 1679585382
transform 1 0 99840 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_259
timestamp 1679585382
transform 1 0 100512 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_266
timestamp 1679585382
transform 1 0 101184 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_273
timestamp 1679585382
transform 1 0 101856 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_280
timestamp 1679585382
transform 1 0 102528 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_287
timestamp 1679585382
transform 1 0 103200 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_294
timestamp 1679585382
transform 1 0 103872 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_301
timestamp 1679585382
transform 1 0 104544 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_308
timestamp 1679585382
transform 1 0 105216 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_315
timestamp 1679585382
transform 1 0 105888 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_322
timestamp 1679585382
transform 1 0 106560 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_329
timestamp 1679585382
transform 1 0 107232 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_336
timestamp 1679585382
transform 1 0 107904 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_343
timestamp 1679585382
transform 1 0 108576 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_350
timestamp 1679585382
transform 1 0 109248 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_357
timestamp 1679585382
transform 1 0 109920 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_364
timestamp 1679585382
transform 1 0 110592 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_371
timestamp 1679585382
transform 1 0 111264 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_378
timestamp 1679585382
transform 1 0 111936 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_385
timestamp 1679585382
transform 1 0 112608 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_392
timestamp 1679585382
transform 1 0 113280 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_399
timestamp 1679585382
transform 1 0 113952 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_406
timestamp 1679585382
transform 1 0 114624 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_413
timestamp 1679585382
transform 1 0 115296 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_420
timestamp 1679585382
transform 1 0 115968 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_427
timestamp 1679585382
transform 1 0 116640 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_434
timestamp 1679585382
transform 1 0 117312 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_441
timestamp 1679585382
transform 1 0 117984 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_448
timestamp 1679585382
transform 1 0 118656 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_455
timestamp 1679585382
transform 1 0 119328 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_462
timestamp 1679585382
transform 1 0 120000 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_469
timestamp 1679585382
transform 1 0 120672 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_476
timestamp 1679585382
transform 1 0 121344 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_483
timestamp 1679585382
transform 1 0 122016 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_490
timestamp 1679585382
transform 1 0 122688 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_497
timestamp 1679585382
transform 1 0 123360 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_504
timestamp 1679585382
transform 1 0 124032 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_511
timestamp 1679585382
transform 1 0 124704 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_518
timestamp 1679585382
transform 1 0 125376 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_525
timestamp 1679585382
transform 1 0 126048 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_532
timestamp 1679585382
transform 1 0 126720 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_539
timestamp 1679585382
transform 1 0 127392 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_546
timestamp 1679585382
transform 1 0 128064 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_553
timestamp 1679585382
transform 1 0 128736 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_560
timestamp 1679585382
transform 1 0 129408 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_567
timestamp 1679585382
transform 1 0 130080 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_574
timestamp 1679585382
transform 1 0 130752 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_581
timestamp 1679585382
transform 1 0 131424 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_588
timestamp 1679585382
transform 1 0 132096 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_595
timestamp 1679585382
transform 1 0 132768 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_602
timestamp 1679585382
transform 1 0 133440 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_609
timestamp 1679585382
transform 1 0 134112 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_616
timestamp 1679585382
transform 1 0 134784 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_623
timestamp 1679585382
transform 1 0 135456 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_630
timestamp 1679585382
transform 1 0 136128 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_637
timestamp 1679585382
transform 1 0 136800 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_644
timestamp 1679585382
transform 1 0 137472 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_651
timestamp 1679585382
transform 1 0 138144 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_658
timestamp 1679585382
transform 1 0 138816 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_665
timestamp 1679585382
transform 1 0 139488 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_672
timestamp 1679585382
transform 1 0 140160 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_679
timestamp 1679585382
transform 1 0 140832 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_686
timestamp 1679585382
transform 1 0 141504 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_693
timestamp 1679585382
transform 1 0 142176 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_700
timestamp 1679585382
transform 1 0 142848 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_707
timestamp 1679585382
transform 1 0 143520 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_714
timestamp 1679585382
transform 1 0 144192 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_721
timestamp 1679585382
transform 1 0 144864 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_728
timestamp 1679585382
transform 1 0 145536 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_735
timestamp 1679585382
transform 1 0 146208 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_742
timestamp 1679585382
transform 1 0 146880 0 -1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_749
timestamp 1679585382
transform 1 0 147552 0 -1 93744
box -48 -56 720 834
use sg13g2_fill_1  FILLER_23_756
timestamp 1677583258
transform 1 0 148224 0 -1 93744
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_0
timestamp 1679585382
transform 1 0 75648 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_7
timestamp 1679585382
transform 1 0 76320 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_14
timestamp 1679585382
transform 1 0 76992 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_21
timestamp 1679585382
transform 1 0 77664 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_28
timestamp 1679585382
transform 1 0 78336 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_35
timestamp 1679585382
transform 1 0 79008 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_42
timestamp 1679585382
transform 1 0 79680 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_49
timestamp 1679585382
transform 1 0 80352 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_56
timestamp 1679585382
transform 1 0 81024 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_63
timestamp 1679585382
transform 1 0 81696 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_70
timestamp 1679585382
transform 1 0 82368 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_77
timestamp 1679585382
transform 1 0 83040 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_84
timestamp 1679585382
transform 1 0 83712 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_91
timestamp 1679585382
transform 1 0 84384 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_98
timestamp 1679585382
transform 1 0 85056 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_105
timestamp 1679585382
transform 1 0 85728 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_112
timestamp 1679585382
transform 1 0 86400 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_119
timestamp 1679585382
transform 1 0 87072 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_126
timestamp 1679585382
transform 1 0 87744 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_133
timestamp 1679585382
transform 1 0 88416 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_140
timestamp 1679585382
transform 1 0 89088 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_147
timestamp 1679585382
transform 1 0 89760 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_154
timestamp 1679585382
transform 1 0 90432 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_161
timestamp 1679585382
transform 1 0 91104 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_168
timestamp 1679585382
transform 1 0 91776 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_175
timestamp 1679585382
transform 1 0 92448 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_182
timestamp 1679585382
transform 1 0 93120 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_189
timestamp 1679585382
transform 1 0 93792 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_196
timestamp 1679585382
transform 1 0 94464 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_203
timestamp 1679585382
transform 1 0 95136 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_210
timestamp 1679585382
transform 1 0 95808 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_217
timestamp 1679585382
transform 1 0 96480 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_224
timestamp 1679585382
transform 1 0 97152 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_231
timestamp 1679585382
transform 1 0 97824 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_238
timestamp 1679585382
transform 1 0 98496 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_245
timestamp 1679585382
transform 1 0 99168 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_252
timestamp 1679585382
transform 1 0 99840 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_259
timestamp 1679585382
transform 1 0 100512 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_266
timestamp 1679585382
transform 1 0 101184 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_273
timestamp 1679585382
transform 1 0 101856 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_280
timestamp 1679585382
transform 1 0 102528 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_287
timestamp 1679585382
transform 1 0 103200 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_294
timestamp 1679585382
transform 1 0 103872 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_301
timestamp 1679585382
transform 1 0 104544 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_308
timestamp 1679585382
transform 1 0 105216 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_315
timestamp 1679585382
transform 1 0 105888 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_322
timestamp 1679585382
transform 1 0 106560 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_329
timestamp 1679585382
transform 1 0 107232 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_336
timestamp 1679585382
transform 1 0 107904 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_343
timestamp 1679585382
transform 1 0 108576 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_350
timestamp 1679585382
transform 1 0 109248 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_357
timestamp 1679585382
transform 1 0 109920 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_364
timestamp 1679585382
transform 1 0 110592 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_371
timestamp 1679585382
transform 1 0 111264 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_378
timestamp 1679585382
transform 1 0 111936 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_385
timestamp 1679585382
transform 1 0 112608 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_392
timestamp 1679585382
transform 1 0 113280 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_399
timestamp 1679585382
transform 1 0 113952 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_406
timestamp 1679585382
transform 1 0 114624 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_413
timestamp 1679585382
transform 1 0 115296 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_420
timestamp 1679585382
transform 1 0 115968 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_427
timestamp 1679585382
transform 1 0 116640 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_434
timestamp 1679585382
transform 1 0 117312 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_441
timestamp 1679585382
transform 1 0 117984 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_448
timestamp 1679585382
transform 1 0 118656 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_455
timestamp 1679585382
transform 1 0 119328 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_462
timestamp 1679585382
transform 1 0 120000 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_469
timestamp 1679585382
transform 1 0 120672 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_476
timestamp 1679585382
transform 1 0 121344 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_483
timestamp 1679585382
transform 1 0 122016 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_490
timestamp 1679585382
transform 1 0 122688 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_497
timestamp 1679585382
transform 1 0 123360 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_504
timestamp 1679585382
transform 1 0 124032 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_511
timestamp 1679585382
transform 1 0 124704 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_518
timestamp 1679585382
transform 1 0 125376 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_525
timestamp 1679585382
transform 1 0 126048 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_532
timestamp 1679585382
transform 1 0 126720 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_539
timestamp 1679585382
transform 1 0 127392 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_546
timestamp 1679585382
transform 1 0 128064 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_553
timestamp 1679585382
transform 1 0 128736 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_560
timestamp 1679585382
transform 1 0 129408 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_567
timestamp 1679585382
transform 1 0 130080 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_574
timestamp 1679585382
transform 1 0 130752 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_581
timestamp 1679585382
transform 1 0 131424 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_588
timestamp 1679585382
transform 1 0 132096 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_595
timestamp 1679585382
transform 1 0 132768 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_602
timestamp 1679585382
transform 1 0 133440 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_609
timestamp 1679585382
transform 1 0 134112 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_616
timestamp 1679585382
transform 1 0 134784 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_623
timestamp 1679585382
transform 1 0 135456 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_630
timestamp 1679585382
transform 1 0 136128 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_637
timestamp 1679585382
transform 1 0 136800 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_644
timestamp 1679585382
transform 1 0 137472 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_651
timestamp 1679585382
transform 1 0 138144 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_658
timestamp 1679585382
transform 1 0 138816 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_665
timestamp 1679585382
transform 1 0 139488 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_672
timestamp 1679585382
transform 1 0 140160 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_679
timestamp 1679585382
transform 1 0 140832 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_686
timestamp 1679585382
transform 1 0 141504 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_693
timestamp 1679585382
transform 1 0 142176 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_700
timestamp 1679585382
transform 1 0 142848 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_707
timestamp 1679585382
transform 1 0 143520 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_714
timestamp 1679585382
transform 1 0 144192 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_721
timestamp 1679585382
transform 1 0 144864 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_728
timestamp 1679585382
transform 1 0 145536 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_735
timestamp 1679585382
transform 1 0 146208 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_742
timestamp 1679585382
transform 1 0 146880 0 1 93744
box -48 -56 720 834
use sg13g2_decap_8  FILLER_24_749
timestamp 1679585382
transform 1 0 147552 0 1 93744
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_756
timestamp 1677583258
transform 1 0 148224 0 1 93744
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_0
timestamp 1679585382
transform 1 0 75648 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_7
timestamp 1679585382
transform 1 0 76320 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_14
timestamp 1679585382
transform 1 0 76992 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_21
timestamp 1679585382
transform 1 0 77664 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_28
timestamp 1679585382
transform 1 0 78336 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_35
timestamp 1679585382
transform 1 0 79008 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_42
timestamp 1679585382
transform 1 0 79680 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_49
timestamp 1679585382
transform 1 0 80352 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_56
timestamp 1679585382
transform 1 0 81024 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_63
timestamp 1679585382
transform 1 0 81696 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_70
timestamp 1679585382
transform 1 0 82368 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_77
timestamp 1679585382
transform 1 0 83040 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_84
timestamp 1679585382
transform 1 0 83712 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_91
timestamp 1679585382
transform 1 0 84384 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_98
timestamp 1679585382
transform 1 0 85056 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_105
timestamp 1679585382
transform 1 0 85728 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_112
timestamp 1679585382
transform 1 0 86400 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_119
timestamp 1679585382
transform 1 0 87072 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_126
timestamp 1679585382
transform 1 0 87744 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_133
timestamp 1679585382
transform 1 0 88416 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_140
timestamp 1679585382
transform 1 0 89088 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_147
timestamp 1679585382
transform 1 0 89760 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_154
timestamp 1679585382
transform 1 0 90432 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_161
timestamp 1679585382
transform 1 0 91104 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_168
timestamp 1679585382
transform 1 0 91776 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_175
timestamp 1679585382
transform 1 0 92448 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_182
timestamp 1679585382
transform 1 0 93120 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_189
timestamp 1679585382
transform 1 0 93792 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_196
timestamp 1679585382
transform 1 0 94464 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_203
timestamp 1679585382
transform 1 0 95136 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_210
timestamp 1679585382
transform 1 0 95808 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_217
timestamp 1679585382
transform 1 0 96480 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_224
timestamp 1679585382
transform 1 0 97152 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_231
timestamp 1679585382
transform 1 0 97824 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_238
timestamp 1679585382
transform 1 0 98496 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_245
timestamp 1679585382
transform 1 0 99168 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_252
timestamp 1679585382
transform 1 0 99840 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_259
timestamp 1679585382
transform 1 0 100512 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_266
timestamp 1679585382
transform 1 0 101184 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_273
timestamp 1679585382
transform 1 0 101856 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_280
timestamp 1679585382
transform 1 0 102528 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_287
timestamp 1679585382
transform 1 0 103200 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_294
timestamp 1679585382
transform 1 0 103872 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_301
timestamp 1679585382
transform 1 0 104544 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_308
timestamp 1679585382
transform 1 0 105216 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_315
timestamp 1679585382
transform 1 0 105888 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_322
timestamp 1679585382
transform 1 0 106560 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_329
timestamp 1679585382
transform 1 0 107232 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_336
timestamp 1679585382
transform 1 0 107904 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_343
timestamp 1679585382
transform 1 0 108576 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_350
timestamp 1679585382
transform 1 0 109248 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_357
timestamp 1679585382
transform 1 0 109920 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_364
timestamp 1679585382
transform 1 0 110592 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_371
timestamp 1679585382
transform 1 0 111264 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_378
timestamp 1679585382
transform 1 0 111936 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_385
timestamp 1679585382
transform 1 0 112608 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_392
timestamp 1679585382
transform 1 0 113280 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_399
timestamp 1679585382
transform 1 0 113952 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_406
timestamp 1679585382
transform 1 0 114624 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_413
timestamp 1679585382
transform 1 0 115296 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_420
timestamp 1679585382
transform 1 0 115968 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_427
timestamp 1679585382
transform 1 0 116640 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_434
timestamp 1679585382
transform 1 0 117312 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_441
timestamp 1679585382
transform 1 0 117984 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_448
timestamp 1679585382
transform 1 0 118656 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_455
timestamp 1679585382
transform 1 0 119328 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_462
timestamp 1679585382
transform 1 0 120000 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_469
timestamp 1679585382
transform 1 0 120672 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_476
timestamp 1679585382
transform 1 0 121344 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_483
timestamp 1679585382
transform 1 0 122016 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_490
timestamp 1679585382
transform 1 0 122688 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_497
timestamp 1679585382
transform 1 0 123360 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_504
timestamp 1679585382
transform 1 0 124032 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_511
timestamp 1679585382
transform 1 0 124704 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_518
timestamp 1679585382
transform 1 0 125376 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_525
timestamp 1679585382
transform 1 0 126048 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_532
timestamp 1679585382
transform 1 0 126720 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_539
timestamp 1679585382
transform 1 0 127392 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_546
timestamp 1679585382
transform 1 0 128064 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_553
timestamp 1679585382
transform 1 0 128736 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_560
timestamp 1679585382
transform 1 0 129408 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_567
timestamp 1679585382
transform 1 0 130080 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_574
timestamp 1679585382
transform 1 0 130752 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_581
timestamp 1679585382
transform 1 0 131424 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_588
timestamp 1679585382
transform 1 0 132096 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_595
timestamp 1679585382
transform 1 0 132768 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_602
timestamp 1679585382
transform 1 0 133440 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_609
timestamp 1679585382
transform 1 0 134112 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_616
timestamp 1679585382
transform 1 0 134784 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_623
timestamp 1679585382
transform 1 0 135456 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_630
timestamp 1679585382
transform 1 0 136128 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_637
timestamp 1679585382
transform 1 0 136800 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_644
timestamp 1679585382
transform 1 0 137472 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_651
timestamp 1679585382
transform 1 0 138144 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_658
timestamp 1679585382
transform 1 0 138816 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_665
timestamp 1679585382
transform 1 0 139488 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_672
timestamp 1679585382
transform 1 0 140160 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_679
timestamp 1679585382
transform 1 0 140832 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_686
timestamp 1679585382
transform 1 0 141504 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_693
timestamp 1679585382
transform 1 0 142176 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_700
timestamp 1679585382
transform 1 0 142848 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_707
timestamp 1679585382
transform 1 0 143520 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_714
timestamp 1679585382
transform 1 0 144192 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_721
timestamp 1679585382
transform 1 0 144864 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_728
timestamp 1679585382
transform 1 0 145536 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_735
timestamp 1679585382
transform 1 0 146208 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_742
timestamp 1679585382
transform 1 0 146880 0 -1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_25_749
timestamp 1679585382
transform 1 0 147552 0 -1 95256
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_756
timestamp 1677583258
transform 1 0 148224 0 -1 95256
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_0
timestamp 1679585382
transform 1 0 75648 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_7
timestamp 1679585382
transform 1 0 76320 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_14
timestamp 1679585382
transform 1 0 76992 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_21
timestamp 1679585382
transform 1 0 77664 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_28
timestamp 1679585382
transform 1 0 78336 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_35
timestamp 1679585382
transform 1 0 79008 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_42
timestamp 1679585382
transform 1 0 79680 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_49
timestamp 1679585382
transform 1 0 80352 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_56
timestamp 1679585382
transform 1 0 81024 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_63
timestamp 1679585382
transform 1 0 81696 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_70
timestamp 1679585382
transform 1 0 82368 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_77
timestamp 1679585382
transform 1 0 83040 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_84
timestamp 1679585382
transform 1 0 83712 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_91
timestamp 1679585382
transform 1 0 84384 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_98
timestamp 1679585382
transform 1 0 85056 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_105
timestamp 1679585382
transform 1 0 85728 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_112
timestamp 1679585382
transform 1 0 86400 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_119
timestamp 1679585382
transform 1 0 87072 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_126
timestamp 1679585382
transform 1 0 87744 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_133
timestamp 1679585382
transform 1 0 88416 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_140
timestamp 1679585382
transform 1 0 89088 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_147
timestamp 1679585382
transform 1 0 89760 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_154
timestamp 1679585382
transform 1 0 90432 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_161
timestamp 1679585382
transform 1 0 91104 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_168
timestamp 1679585382
transform 1 0 91776 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_175
timestamp 1679585382
transform 1 0 92448 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_182
timestamp 1679585382
transform 1 0 93120 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_189
timestamp 1679585382
transform 1 0 93792 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_196
timestamp 1679585382
transform 1 0 94464 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_203
timestamp 1679585382
transform 1 0 95136 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_210
timestamp 1679585382
transform 1 0 95808 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_217
timestamp 1679585382
transform 1 0 96480 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_224
timestamp 1679585382
transform 1 0 97152 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_231
timestamp 1679585382
transform 1 0 97824 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_238
timestamp 1679585382
transform 1 0 98496 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_245
timestamp 1679585382
transform 1 0 99168 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_252
timestamp 1679585382
transform 1 0 99840 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_259
timestamp 1679585382
transform 1 0 100512 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_266
timestamp 1679585382
transform 1 0 101184 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_273
timestamp 1679585382
transform 1 0 101856 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_280
timestamp 1679585382
transform 1 0 102528 0 1 95256
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_287
timestamp 1679581501
transform 1 0 103200 0 1 95256
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_300
timestamp 1679585382
transform 1 0 104448 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_307
timestamp 1679585382
transform 1 0 105120 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_314
timestamp 1679585382
transform 1 0 105792 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_321
timestamp 1679585382
transform 1 0 106464 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_328
timestamp 1679585382
transform 1 0 107136 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_335
timestamp 1679585382
transform 1 0 107808 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_342
timestamp 1679585382
transform 1 0 108480 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_349
timestamp 1679585382
transform 1 0 109152 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_356
timestamp 1679585382
transform 1 0 109824 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_363
timestamp 1679585382
transform 1 0 110496 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_370
timestamp 1679585382
transform 1 0 111168 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_377
timestamp 1679585382
transform 1 0 111840 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_384
timestamp 1679585382
transform 1 0 112512 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_391
timestamp 1679585382
transform 1 0 113184 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_398
timestamp 1679585382
transform 1 0 113856 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_405
timestamp 1679585382
transform 1 0 114528 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_412
timestamp 1679585382
transform 1 0 115200 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_419
timestamp 1679585382
transform 1 0 115872 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_426
timestamp 1679585382
transform 1 0 116544 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_433
timestamp 1679585382
transform 1 0 117216 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_440
timestamp 1679585382
transform 1 0 117888 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_447
timestamp 1679585382
transform 1 0 118560 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_454
timestamp 1679585382
transform 1 0 119232 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_461
timestamp 1679585382
transform 1 0 119904 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_468
timestamp 1679585382
transform 1 0 120576 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_475
timestamp 1679585382
transform 1 0 121248 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_482
timestamp 1679585382
transform 1 0 121920 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_489
timestamp 1679585382
transform 1 0 122592 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_496
timestamp 1679585382
transform 1 0 123264 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_503
timestamp 1679585382
transform 1 0 123936 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_510
timestamp 1679585382
transform 1 0 124608 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_517
timestamp 1679585382
transform 1 0 125280 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_524
timestamp 1679585382
transform 1 0 125952 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_531
timestamp 1679585382
transform 1 0 126624 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_538
timestamp 1679585382
transform 1 0 127296 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_545
timestamp 1679585382
transform 1 0 127968 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_552
timestamp 1679585382
transform 1 0 128640 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_559
timestamp 1679585382
transform 1 0 129312 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_566
timestamp 1679585382
transform 1 0 129984 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_573
timestamp 1679585382
transform 1 0 130656 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_580
timestamp 1679585382
transform 1 0 131328 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_587
timestamp 1679585382
transform 1 0 132000 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_594
timestamp 1679585382
transform 1 0 132672 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_601
timestamp 1679585382
transform 1 0 133344 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_608
timestamp 1679585382
transform 1 0 134016 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_615
timestamp 1679585382
transform 1 0 134688 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_622
timestamp 1679585382
transform 1 0 135360 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_629
timestamp 1679585382
transform 1 0 136032 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_636
timestamp 1679585382
transform 1 0 136704 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_643
timestamp 1679585382
transform 1 0 137376 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_650
timestamp 1679585382
transform 1 0 138048 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_657
timestamp 1679585382
transform 1 0 138720 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_664
timestamp 1679585382
transform 1 0 139392 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_671
timestamp 1679585382
transform 1 0 140064 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_678
timestamp 1679585382
transform 1 0 140736 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_685
timestamp 1679585382
transform 1 0 141408 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_692
timestamp 1679585382
transform 1 0 142080 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_699
timestamp 1679585382
transform 1 0 142752 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_706
timestamp 1679585382
transform 1 0 143424 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_713
timestamp 1679585382
transform 1 0 144096 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_720
timestamp 1679585382
transform 1 0 144768 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_727
timestamp 1679585382
transform 1 0 145440 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_734
timestamp 1679585382
transform 1 0 146112 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_741
timestamp 1679585382
transform 1 0 146784 0 1 95256
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_748
timestamp 1679585382
transform 1 0 147456 0 1 95256
box -48 -56 720 834
use sg13g2_fill_2  FILLER_26_755
timestamp 1677583704
transform 1 0 148128 0 1 95256
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679585382
transform 1 0 75648 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_7
timestamp 1679585382
transform 1 0 76320 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_14
timestamp 1679585382
transform 1 0 76992 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_21
timestamp 1679585382
transform 1 0 77664 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_28
timestamp 1679585382
transform 1 0 78336 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_35
timestamp 1679585382
transform 1 0 79008 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_42
timestamp 1679585382
transform 1 0 79680 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_49
timestamp 1679585382
transform 1 0 80352 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_56
timestamp 1679585382
transform 1 0 81024 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_63
timestamp 1679585382
transform 1 0 81696 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_70
timestamp 1679585382
transform 1 0 82368 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_77
timestamp 1679585382
transform 1 0 83040 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_84
timestamp 1679585382
transform 1 0 83712 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_91
timestamp 1679585382
transform 1 0 84384 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_98
timestamp 1679585382
transform 1 0 85056 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_105
timestamp 1679585382
transform 1 0 85728 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_112
timestamp 1679585382
transform 1 0 86400 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_119
timestamp 1679585382
transform 1 0 87072 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_126
timestamp 1679585382
transform 1 0 87744 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_133
timestamp 1679585382
transform 1 0 88416 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_140
timestamp 1679585382
transform 1 0 89088 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_147
timestamp 1679585382
transform 1 0 89760 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_154
timestamp 1679585382
transform 1 0 90432 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_161
timestamp 1679585382
transform 1 0 91104 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_168
timestamp 1679585382
transform 1 0 91776 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_175
timestamp 1679585382
transform 1 0 92448 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_182
timestamp 1679585382
transform 1 0 93120 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_189
timestamp 1679585382
transform 1 0 93792 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_196
timestamp 1679585382
transform 1 0 94464 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_203
timestamp 1679585382
transform 1 0 95136 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_210
timestamp 1679585382
transform 1 0 95808 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_217
timestamp 1679585382
transform 1 0 96480 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_224
timestamp 1679585382
transform 1 0 97152 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_231
timestamp 1679585382
transform 1 0 97824 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_238
timestamp 1679585382
transform 1 0 98496 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_245
timestamp 1679585382
transform 1 0 99168 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_252
timestamp 1679585382
transform 1 0 99840 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_259
timestamp 1679585382
transform 1 0 100512 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_266
timestamp 1679585382
transform 1 0 101184 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_273
timestamp 1679585382
transform 1 0 101856 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_280
timestamp 1679585382
transform 1 0 102528 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_287
timestamp 1679585382
transform 1 0 103200 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_294
timestamp 1679585382
transform 1 0 103872 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_301
timestamp 1679585382
transform 1 0 104544 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_308
timestamp 1679585382
transform 1 0 105216 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_315
timestamp 1679585382
transform 1 0 105888 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_322
timestamp 1679585382
transform 1 0 106560 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_329
timestamp 1679585382
transform 1 0 107232 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_336
timestamp 1679585382
transform 1 0 107904 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_343
timestamp 1679585382
transform 1 0 108576 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_350
timestamp 1679585382
transform 1 0 109248 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_357
timestamp 1679585382
transform 1 0 109920 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_364
timestamp 1679585382
transform 1 0 110592 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_371
timestamp 1679585382
transform 1 0 111264 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_378
timestamp 1679585382
transform 1 0 111936 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_385
timestamp 1679585382
transform 1 0 112608 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_392
timestamp 1679585382
transform 1 0 113280 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_399
timestamp 1679585382
transform 1 0 113952 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_406
timestamp 1679585382
transform 1 0 114624 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_413
timestamp 1679585382
transform 1 0 115296 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_420
timestamp 1679585382
transform 1 0 115968 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_427
timestamp 1679585382
transform 1 0 116640 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_434
timestamp 1679585382
transform 1 0 117312 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_441
timestamp 1679585382
transform 1 0 117984 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_448
timestamp 1679585382
transform 1 0 118656 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_455
timestamp 1679585382
transform 1 0 119328 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_462
timestamp 1679585382
transform 1 0 120000 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_469
timestamp 1679585382
transform 1 0 120672 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_476
timestamp 1679585382
transform 1 0 121344 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_483
timestamp 1679585382
transform 1 0 122016 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_490
timestamp 1679585382
transform 1 0 122688 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_497
timestamp 1679585382
transform 1 0 123360 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_504
timestamp 1679585382
transform 1 0 124032 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_511
timestamp 1679585382
transform 1 0 124704 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_518
timestamp 1679585382
transform 1 0 125376 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_525
timestamp 1679585382
transform 1 0 126048 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_532
timestamp 1679585382
transform 1 0 126720 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_539
timestamp 1679585382
transform 1 0 127392 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_546
timestamp 1679585382
transform 1 0 128064 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_553
timestamp 1679585382
transform 1 0 128736 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_560
timestamp 1679585382
transform 1 0 129408 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_567
timestamp 1679585382
transform 1 0 130080 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_574
timestamp 1679585382
transform 1 0 130752 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_581
timestamp 1679585382
transform 1 0 131424 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_588
timestamp 1679585382
transform 1 0 132096 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_595
timestamp 1679585382
transform 1 0 132768 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_602
timestamp 1679585382
transform 1 0 133440 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_609
timestamp 1679585382
transform 1 0 134112 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_616
timestamp 1679585382
transform 1 0 134784 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_623
timestamp 1679585382
transform 1 0 135456 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_630
timestamp 1679585382
transform 1 0 136128 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_637
timestamp 1679585382
transform 1 0 136800 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_644
timestamp 1679585382
transform 1 0 137472 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_651
timestamp 1679585382
transform 1 0 138144 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_658
timestamp 1679585382
transform 1 0 138816 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_665
timestamp 1679585382
transform 1 0 139488 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_672
timestamp 1679585382
transform 1 0 140160 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_679
timestamp 1679585382
transform 1 0 140832 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_686
timestamp 1679585382
transform 1 0 141504 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_693
timestamp 1679585382
transform 1 0 142176 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_700
timestamp 1679585382
transform 1 0 142848 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_707
timestamp 1679585382
transform 1 0 143520 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_714
timestamp 1679585382
transform 1 0 144192 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_721
timestamp 1679585382
transform 1 0 144864 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_728
timestamp 1679585382
transform 1 0 145536 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_735
timestamp 1679585382
transform 1 0 146208 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_742
timestamp 1679585382
transform 1 0 146880 0 -1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_749
timestamp 1679585382
transform 1 0 147552 0 -1 96768
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_756
timestamp 1677583258
transform 1 0 148224 0 -1 96768
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_0
timestamp 1679585382
transform 1 0 75648 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_7
timestamp 1679585382
transform 1 0 76320 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_14
timestamp 1679585382
transform 1 0 76992 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_21
timestamp 1679585382
transform 1 0 77664 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_28
timestamp 1679585382
transform 1 0 78336 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_35
timestamp 1679585382
transform 1 0 79008 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_42
timestamp 1679585382
transform 1 0 79680 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_49
timestamp 1679585382
transform 1 0 80352 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_56
timestamp 1679585382
transform 1 0 81024 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_63
timestamp 1679585382
transform 1 0 81696 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_70
timestamp 1679585382
transform 1 0 82368 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_77
timestamp 1679585382
transform 1 0 83040 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_84
timestamp 1679585382
transform 1 0 83712 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_91
timestamp 1679585382
transform 1 0 84384 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_98
timestamp 1679585382
transform 1 0 85056 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_105
timestamp 1679585382
transform 1 0 85728 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_112
timestamp 1679585382
transform 1 0 86400 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_119
timestamp 1679585382
transform 1 0 87072 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_126
timestamp 1679585382
transform 1 0 87744 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_133
timestamp 1679585382
transform 1 0 88416 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_140
timestamp 1679585382
transform 1 0 89088 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_147
timestamp 1679585382
transform 1 0 89760 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_154
timestamp 1679585382
transform 1 0 90432 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_161
timestamp 1679585382
transform 1 0 91104 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_168
timestamp 1679585382
transform 1 0 91776 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_175
timestamp 1679585382
transform 1 0 92448 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_182
timestamp 1679585382
transform 1 0 93120 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_189
timestamp 1679585382
transform 1 0 93792 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_196
timestamp 1679585382
transform 1 0 94464 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_203
timestamp 1679585382
transform 1 0 95136 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_210
timestamp 1679585382
transform 1 0 95808 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_217
timestamp 1679585382
transform 1 0 96480 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_224
timestamp 1679585382
transform 1 0 97152 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_231
timestamp 1679585382
transform 1 0 97824 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_238
timestamp 1679585382
transform 1 0 98496 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_245
timestamp 1679585382
transform 1 0 99168 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_252
timestamp 1679585382
transform 1 0 99840 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_259
timestamp 1679585382
transform 1 0 100512 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_266
timestamp 1679585382
transform 1 0 101184 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_273
timestamp 1679585382
transform 1 0 101856 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_280
timestamp 1679585382
transform 1 0 102528 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_287
timestamp 1679585382
transform 1 0 103200 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_294
timestamp 1679585382
transform 1 0 103872 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_301
timestamp 1679585382
transform 1 0 104544 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_308
timestamp 1679585382
transform 1 0 105216 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_315
timestamp 1679585382
transform 1 0 105888 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_322
timestamp 1679585382
transform 1 0 106560 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_329
timestamp 1679585382
transform 1 0 107232 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_336
timestamp 1679585382
transform 1 0 107904 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_343
timestamp 1679585382
transform 1 0 108576 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_350
timestamp 1679585382
transform 1 0 109248 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_357
timestamp 1679585382
transform 1 0 109920 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_364
timestamp 1679585382
transform 1 0 110592 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_371
timestamp 1679585382
transform 1 0 111264 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_378
timestamp 1679585382
transform 1 0 111936 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_385
timestamp 1679585382
transform 1 0 112608 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_392
timestamp 1679585382
transform 1 0 113280 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_399
timestamp 1679585382
transform 1 0 113952 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_406
timestamp 1679585382
transform 1 0 114624 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_413
timestamp 1679585382
transform 1 0 115296 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_420
timestamp 1679585382
transform 1 0 115968 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_427
timestamp 1679585382
transform 1 0 116640 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_434
timestamp 1679585382
transform 1 0 117312 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_441
timestamp 1679585382
transform 1 0 117984 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_448
timestamp 1679585382
transform 1 0 118656 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_455
timestamp 1679585382
transform 1 0 119328 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_462
timestamp 1679585382
transform 1 0 120000 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_469
timestamp 1679585382
transform 1 0 120672 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_476
timestamp 1679585382
transform 1 0 121344 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_483
timestamp 1679585382
transform 1 0 122016 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_490
timestamp 1679585382
transform 1 0 122688 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_497
timestamp 1679585382
transform 1 0 123360 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_504
timestamp 1679585382
transform 1 0 124032 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_511
timestamp 1679585382
transform 1 0 124704 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_518
timestamp 1679585382
transform 1 0 125376 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_525
timestamp 1679585382
transform 1 0 126048 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_532
timestamp 1679585382
transform 1 0 126720 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_539
timestamp 1679585382
transform 1 0 127392 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_546
timestamp 1679585382
transform 1 0 128064 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_553
timestamp 1679585382
transform 1 0 128736 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_560
timestamp 1679585382
transform 1 0 129408 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_567
timestamp 1679585382
transform 1 0 130080 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_574
timestamp 1679585382
transform 1 0 130752 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_581
timestamp 1679585382
transform 1 0 131424 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_588
timestamp 1679585382
transform 1 0 132096 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_595
timestamp 1679585382
transform 1 0 132768 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_602
timestamp 1679585382
transform 1 0 133440 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_609
timestamp 1679585382
transform 1 0 134112 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_616
timestamp 1679585382
transform 1 0 134784 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_623
timestamp 1679585382
transform 1 0 135456 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_630
timestamp 1679585382
transform 1 0 136128 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_637
timestamp 1679585382
transform 1 0 136800 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_644
timestamp 1679585382
transform 1 0 137472 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_651
timestamp 1679585382
transform 1 0 138144 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_658
timestamp 1679585382
transform 1 0 138816 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_665
timestamp 1679585382
transform 1 0 139488 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_672
timestamp 1679585382
transform 1 0 140160 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_679
timestamp 1679585382
transform 1 0 140832 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_686
timestamp 1679585382
transform 1 0 141504 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_693
timestamp 1679585382
transform 1 0 142176 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_700
timestamp 1679585382
transform 1 0 142848 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_707
timestamp 1679585382
transform 1 0 143520 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_714
timestamp 1679585382
transform 1 0 144192 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_721
timestamp 1679585382
transform 1 0 144864 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_728
timestamp 1679585382
transform 1 0 145536 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_735
timestamp 1679585382
transform 1 0 146208 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_742
timestamp 1679585382
transform 1 0 146880 0 1 96768
box -48 -56 720 834
use sg13g2_decap_8  FILLER_28_749
timestamp 1679585382
transform 1 0 147552 0 1 96768
box -48 -56 720 834
use sg13g2_fill_1  FILLER_28_756
timestamp 1677583258
transform 1 0 148224 0 1 96768
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_0
timestamp 1679585382
transform 1 0 75648 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_7
timestamp 1679585382
transform 1 0 76320 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_14
timestamp 1679585382
transform 1 0 76992 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_21
timestamp 1679585382
transform 1 0 77664 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_28
timestamp 1679585382
transform 1 0 78336 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_35
timestamp 1679585382
transform 1 0 79008 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_42
timestamp 1679585382
transform 1 0 79680 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_49
timestamp 1679585382
transform 1 0 80352 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_56
timestamp 1679585382
transform 1 0 81024 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_63
timestamp 1679585382
transform 1 0 81696 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_70
timestamp 1679585382
transform 1 0 82368 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_77
timestamp 1679585382
transform 1 0 83040 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_84
timestamp 1679585382
transform 1 0 83712 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_91
timestamp 1679585382
transform 1 0 84384 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_98
timestamp 1679585382
transform 1 0 85056 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_105
timestamp 1679585382
transform 1 0 85728 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_112
timestamp 1679585382
transform 1 0 86400 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_119
timestamp 1679585382
transform 1 0 87072 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_126
timestamp 1679585382
transform 1 0 87744 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_133
timestamp 1679585382
transform 1 0 88416 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_140
timestamp 1679585382
transform 1 0 89088 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_147
timestamp 1679585382
transform 1 0 89760 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_154
timestamp 1679585382
transform 1 0 90432 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_161
timestamp 1679585382
transform 1 0 91104 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_168
timestamp 1679585382
transform 1 0 91776 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_175
timestamp 1679585382
transform 1 0 92448 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_182
timestamp 1679585382
transform 1 0 93120 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_189
timestamp 1679585382
transform 1 0 93792 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_196
timestamp 1679585382
transform 1 0 94464 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_203
timestamp 1679585382
transform 1 0 95136 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_210
timestamp 1679585382
transform 1 0 95808 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_217
timestamp 1679585382
transform 1 0 96480 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_224
timestamp 1679585382
transform 1 0 97152 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_231
timestamp 1679585382
transform 1 0 97824 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_238
timestamp 1679585382
transform 1 0 98496 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_245
timestamp 1679585382
transform 1 0 99168 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_252
timestamp 1679585382
transform 1 0 99840 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_259
timestamp 1679585382
transform 1 0 100512 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_266
timestamp 1679585382
transform 1 0 101184 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_273
timestamp 1679585382
transform 1 0 101856 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_280
timestamp 1679585382
transform 1 0 102528 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_287
timestamp 1679585382
transform 1 0 103200 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_294
timestamp 1679585382
transform 1 0 103872 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_301
timestamp 1679585382
transform 1 0 104544 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_308
timestamp 1679585382
transform 1 0 105216 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_315
timestamp 1679585382
transform 1 0 105888 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_322
timestamp 1679585382
transform 1 0 106560 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_329
timestamp 1679585382
transform 1 0 107232 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_336
timestamp 1679585382
transform 1 0 107904 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_343
timestamp 1679585382
transform 1 0 108576 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_350
timestamp 1679585382
transform 1 0 109248 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_357
timestamp 1679585382
transform 1 0 109920 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_364
timestamp 1679585382
transform 1 0 110592 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_371
timestamp 1679585382
transform 1 0 111264 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_378
timestamp 1679585382
transform 1 0 111936 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_385
timestamp 1679585382
transform 1 0 112608 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_392
timestamp 1679585382
transform 1 0 113280 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_399
timestamp 1679585382
transform 1 0 113952 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_406
timestamp 1679585382
transform 1 0 114624 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_413
timestamp 1679585382
transform 1 0 115296 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_420
timestamp 1679585382
transform 1 0 115968 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_427
timestamp 1679585382
transform 1 0 116640 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_434
timestamp 1679585382
transform 1 0 117312 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_441
timestamp 1679585382
transform 1 0 117984 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_448
timestamp 1679585382
transform 1 0 118656 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_455
timestamp 1679585382
transform 1 0 119328 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_462
timestamp 1679585382
transform 1 0 120000 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_469
timestamp 1679585382
transform 1 0 120672 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_476
timestamp 1679585382
transform 1 0 121344 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_483
timestamp 1679585382
transform 1 0 122016 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_490
timestamp 1679585382
transform 1 0 122688 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_497
timestamp 1679585382
transform 1 0 123360 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_504
timestamp 1679585382
transform 1 0 124032 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_511
timestamp 1679585382
transform 1 0 124704 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_518
timestamp 1679585382
transform 1 0 125376 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_525
timestamp 1679585382
transform 1 0 126048 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_532
timestamp 1679585382
transform 1 0 126720 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_539
timestamp 1679585382
transform 1 0 127392 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_546
timestamp 1679585382
transform 1 0 128064 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_553
timestamp 1679585382
transform 1 0 128736 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_560
timestamp 1679585382
transform 1 0 129408 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_567
timestamp 1679585382
transform 1 0 130080 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_574
timestamp 1679585382
transform 1 0 130752 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_581
timestamp 1679585382
transform 1 0 131424 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_588
timestamp 1679585382
transform 1 0 132096 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_595
timestamp 1679585382
transform 1 0 132768 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_602
timestamp 1679585382
transform 1 0 133440 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_609
timestamp 1679585382
transform 1 0 134112 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_616
timestamp 1679585382
transform 1 0 134784 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_623
timestamp 1679585382
transform 1 0 135456 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_630
timestamp 1679585382
transform 1 0 136128 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_637
timestamp 1679585382
transform 1 0 136800 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_644
timestamp 1679585382
transform 1 0 137472 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_651
timestamp 1679585382
transform 1 0 138144 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_658
timestamp 1679585382
transform 1 0 138816 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_665
timestamp 1679585382
transform 1 0 139488 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_672
timestamp 1679585382
transform 1 0 140160 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_679
timestamp 1679585382
transform 1 0 140832 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_686
timestamp 1679585382
transform 1 0 141504 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_693
timestamp 1679585382
transform 1 0 142176 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_700
timestamp 1679585382
transform 1 0 142848 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_707
timestamp 1679585382
transform 1 0 143520 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_714
timestamp 1679585382
transform 1 0 144192 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_721
timestamp 1679585382
transform 1 0 144864 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_728
timestamp 1679585382
transform 1 0 145536 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_735
timestamp 1679585382
transform 1 0 146208 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_742
timestamp 1679585382
transform 1 0 146880 0 -1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_29_749
timestamp 1679585382
transform 1 0 147552 0 -1 98280
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_756
timestamp 1677583258
transform 1 0 148224 0 -1 98280
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_0
timestamp 1679585382
transform 1 0 75648 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_7
timestamp 1679585382
transform 1 0 76320 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_14
timestamp 1679585382
transform 1 0 76992 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_21
timestamp 1679585382
transform 1 0 77664 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_28
timestamp 1679585382
transform 1 0 78336 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_35
timestamp 1679585382
transform 1 0 79008 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_42
timestamp 1679585382
transform 1 0 79680 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_49
timestamp 1679585382
transform 1 0 80352 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_56
timestamp 1679585382
transform 1 0 81024 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_63
timestamp 1679585382
transform 1 0 81696 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_70
timestamp 1679585382
transform 1 0 82368 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_77
timestamp 1679585382
transform 1 0 83040 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_84
timestamp 1679585382
transform 1 0 83712 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_91
timestamp 1679585382
transform 1 0 84384 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_98
timestamp 1679585382
transform 1 0 85056 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_105
timestamp 1679585382
transform 1 0 85728 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_112
timestamp 1679585382
transform 1 0 86400 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_119
timestamp 1679585382
transform 1 0 87072 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_126
timestamp 1679585382
transform 1 0 87744 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_133
timestamp 1679585382
transform 1 0 88416 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_140
timestamp 1679585382
transform 1 0 89088 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_147
timestamp 1679585382
transform 1 0 89760 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_154
timestamp 1679585382
transform 1 0 90432 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_161
timestamp 1679585382
transform 1 0 91104 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_168
timestamp 1679585382
transform 1 0 91776 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_175
timestamp 1679585382
transform 1 0 92448 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_182
timestamp 1679585382
transform 1 0 93120 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_189
timestamp 1679585382
transform 1 0 93792 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_196
timestamp 1679585382
transform 1 0 94464 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_203
timestamp 1679585382
transform 1 0 95136 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_210
timestamp 1679585382
transform 1 0 95808 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_217
timestamp 1679585382
transform 1 0 96480 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_224
timestamp 1679585382
transform 1 0 97152 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_231
timestamp 1679585382
transform 1 0 97824 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_238
timestamp 1679585382
transform 1 0 98496 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_245
timestamp 1679585382
transform 1 0 99168 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_252
timestamp 1679585382
transform 1 0 99840 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_259
timestamp 1679585382
transform 1 0 100512 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_266
timestamp 1679585382
transform 1 0 101184 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_273
timestamp 1679585382
transform 1 0 101856 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_280
timestamp 1679585382
transform 1 0 102528 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_287
timestamp 1679585382
transform 1 0 103200 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_294
timestamp 1679585382
transform 1 0 103872 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_301
timestamp 1679585382
transform 1 0 104544 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_308
timestamp 1679585382
transform 1 0 105216 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_315
timestamp 1679585382
transform 1 0 105888 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_322
timestamp 1679585382
transform 1 0 106560 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_329
timestamp 1679585382
transform 1 0 107232 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_336
timestamp 1679585382
transform 1 0 107904 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_343
timestamp 1679585382
transform 1 0 108576 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_350
timestamp 1679585382
transform 1 0 109248 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_357
timestamp 1679585382
transform 1 0 109920 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_364
timestamp 1679585382
transform 1 0 110592 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_371
timestamp 1679585382
transform 1 0 111264 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_378
timestamp 1679585382
transform 1 0 111936 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_385
timestamp 1679585382
transform 1 0 112608 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_392
timestamp 1679585382
transform 1 0 113280 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_399
timestamp 1679585382
transform 1 0 113952 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_406
timestamp 1679585382
transform 1 0 114624 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_413
timestamp 1679585382
transform 1 0 115296 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_420
timestamp 1679585382
transform 1 0 115968 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_427
timestamp 1679585382
transform 1 0 116640 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_434
timestamp 1679585382
transform 1 0 117312 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_441
timestamp 1679585382
transform 1 0 117984 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_448
timestamp 1679585382
transform 1 0 118656 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_455
timestamp 1679585382
transform 1 0 119328 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_462
timestamp 1679585382
transform 1 0 120000 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_469
timestamp 1679585382
transform 1 0 120672 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_476
timestamp 1679585382
transform 1 0 121344 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_483
timestamp 1679585382
transform 1 0 122016 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_490
timestamp 1679585382
transform 1 0 122688 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_497
timestamp 1679585382
transform 1 0 123360 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_504
timestamp 1679585382
transform 1 0 124032 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_511
timestamp 1679585382
transform 1 0 124704 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_518
timestamp 1679585382
transform 1 0 125376 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_525
timestamp 1679585382
transform 1 0 126048 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_532
timestamp 1679585382
transform 1 0 126720 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_539
timestamp 1679585382
transform 1 0 127392 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_546
timestamp 1679585382
transform 1 0 128064 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_553
timestamp 1679585382
transform 1 0 128736 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_560
timestamp 1679585382
transform 1 0 129408 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_567
timestamp 1679585382
transform 1 0 130080 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_574
timestamp 1679585382
transform 1 0 130752 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_581
timestamp 1679585382
transform 1 0 131424 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_588
timestamp 1679585382
transform 1 0 132096 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_595
timestamp 1679585382
transform 1 0 132768 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_602
timestamp 1679585382
transform 1 0 133440 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_609
timestamp 1679585382
transform 1 0 134112 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_616
timestamp 1679585382
transform 1 0 134784 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_623
timestamp 1679585382
transform 1 0 135456 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_630
timestamp 1679585382
transform 1 0 136128 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_637
timestamp 1679585382
transform 1 0 136800 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_644
timestamp 1679585382
transform 1 0 137472 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_651
timestamp 1679585382
transform 1 0 138144 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_658
timestamp 1679585382
transform 1 0 138816 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_665
timestamp 1679585382
transform 1 0 139488 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_672
timestamp 1679585382
transform 1 0 140160 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_679
timestamp 1679585382
transform 1 0 140832 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_686
timestamp 1679585382
transform 1 0 141504 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_693
timestamp 1679585382
transform 1 0 142176 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_700
timestamp 1679585382
transform 1 0 142848 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_707
timestamp 1679585382
transform 1 0 143520 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_714
timestamp 1679585382
transform 1 0 144192 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_721
timestamp 1679585382
transform 1 0 144864 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_728
timestamp 1679585382
transform 1 0 145536 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_735
timestamp 1679585382
transform 1 0 146208 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_742
timestamp 1679585382
transform 1 0 146880 0 1 98280
box -48 -56 720 834
use sg13g2_decap_8  FILLER_30_749
timestamp 1679585382
transform 1 0 147552 0 1 98280
box -48 -56 720 834
use sg13g2_fill_1  FILLER_30_756
timestamp 1677583258
transform 1 0 148224 0 1 98280
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_0
timestamp 1679585382
transform 1 0 75648 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_7
timestamp 1679585382
transform 1 0 76320 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_14
timestamp 1679585382
transform 1 0 76992 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_21
timestamp 1679585382
transform 1 0 77664 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_28
timestamp 1679585382
transform 1 0 78336 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_35
timestamp 1679585382
transform 1 0 79008 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_42
timestamp 1679585382
transform 1 0 79680 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_49
timestamp 1679585382
transform 1 0 80352 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_56
timestamp 1679585382
transform 1 0 81024 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_63
timestamp 1679585382
transform 1 0 81696 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_70
timestamp 1679585382
transform 1 0 82368 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_77
timestamp 1679585382
transform 1 0 83040 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_84
timestamp 1679585382
transform 1 0 83712 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_91
timestamp 1679585382
transform 1 0 84384 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_98
timestamp 1679585382
transform 1 0 85056 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_105
timestamp 1679585382
transform 1 0 85728 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_112
timestamp 1679585382
transform 1 0 86400 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_119
timestamp 1679585382
transform 1 0 87072 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_126
timestamp 1679585382
transform 1 0 87744 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_133
timestamp 1679585382
transform 1 0 88416 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_140
timestamp 1679585382
transform 1 0 89088 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_147
timestamp 1679585382
transform 1 0 89760 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_154
timestamp 1679585382
transform 1 0 90432 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_161
timestamp 1679585382
transform 1 0 91104 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_168
timestamp 1679585382
transform 1 0 91776 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_175
timestamp 1679585382
transform 1 0 92448 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_182
timestamp 1679585382
transform 1 0 93120 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_189
timestamp 1679585382
transform 1 0 93792 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_196
timestamp 1679585382
transform 1 0 94464 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_203
timestamp 1679585382
transform 1 0 95136 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_210
timestamp 1679585382
transform 1 0 95808 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_217
timestamp 1679585382
transform 1 0 96480 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_224
timestamp 1679585382
transform 1 0 97152 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_231
timestamp 1679585382
transform 1 0 97824 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_238
timestamp 1679585382
transform 1 0 98496 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_245
timestamp 1679585382
transform 1 0 99168 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_252
timestamp 1679585382
transform 1 0 99840 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_259
timestamp 1679585382
transform 1 0 100512 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_266
timestamp 1679585382
transform 1 0 101184 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_273
timestamp 1679585382
transform 1 0 101856 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_280
timestamp 1679585382
transform 1 0 102528 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_287
timestamp 1679585382
transform 1 0 103200 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_294
timestamp 1679585382
transform 1 0 103872 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_301
timestamp 1679585382
transform 1 0 104544 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_308
timestamp 1679585382
transform 1 0 105216 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_315
timestamp 1679585382
transform 1 0 105888 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_322
timestamp 1679585382
transform 1 0 106560 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_329
timestamp 1679585382
transform 1 0 107232 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_336
timestamp 1679585382
transform 1 0 107904 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_343
timestamp 1679585382
transform 1 0 108576 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_350
timestamp 1679585382
transform 1 0 109248 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_357
timestamp 1679585382
transform 1 0 109920 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_364
timestamp 1679585382
transform 1 0 110592 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_371
timestamp 1679585382
transform 1 0 111264 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_378
timestamp 1679585382
transform 1 0 111936 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_385
timestamp 1679585382
transform 1 0 112608 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_392
timestamp 1679585382
transform 1 0 113280 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_399
timestamp 1679585382
transform 1 0 113952 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_406
timestamp 1679585382
transform 1 0 114624 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_413
timestamp 1679585382
transform 1 0 115296 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_420
timestamp 1679585382
transform 1 0 115968 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_427
timestamp 1679585382
transform 1 0 116640 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_434
timestamp 1679585382
transform 1 0 117312 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_441
timestamp 1679585382
transform 1 0 117984 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_448
timestamp 1679585382
transform 1 0 118656 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_455
timestamp 1679585382
transform 1 0 119328 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_462
timestamp 1679585382
transform 1 0 120000 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_469
timestamp 1679585382
transform 1 0 120672 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_476
timestamp 1679585382
transform 1 0 121344 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_483
timestamp 1679585382
transform 1 0 122016 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_490
timestamp 1679585382
transform 1 0 122688 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_497
timestamp 1679585382
transform 1 0 123360 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_504
timestamp 1679585382
transform 1 0 124032 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_511
timestamp 1679585382
transform 1 0 124704 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_518
timestamp 1679585382
transform 1 0 125376 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_525
timestamp 1679585382
transform 1 0 126048 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_532
timestamp 1679585382
transform 1 0 126720 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_539
timestamp 1679585382
transform 1 0 127392 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_546
timestamp 1679585382
transform 1 0 128064 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_553
timestamp 1679585382
transform 1 0 128736 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_560
timestamp 1679585382
transform 1 0 129408 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_567
timestamp 1679585382
transform 1 0 130080 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_574
timestamp 1679585382
transform 1 0 130752 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_581
timestamp 1679585382
transform 1 0 131424 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_588
timestamp 1679585382
transform 1 0 132096 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_595
timestamp 1679585382
transform 1 0 132768 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_602
timestamp 1679585382
transform 1 0 133440 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_609
timestamp 1679585382
transform 1 0 134112 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_616
timestamp 1679585382
transform 1 0 134784 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_623
timestamp 1679585382
transform 1 0 135456 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_630
timestamp 1679585382
transform 1 0 136128 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_637
timestamp 1679585382
transform 1 0 136800 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_644
timestamp 1679585382
transform 1 0 137472 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_651
timestamp 1679585382
transform 1 0 138144 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_658
timestamp 1679585382
transform 1 0 138816 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_665
timestamp 1679585382
transform 1 0 139488 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_672
timestamp 1679585382
transform 1 0 140160 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_679
timestamp 1679585382
transform 1 0 140832 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_686
timestamp 1679585382
transform 1 0 141504 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_693
timestamp 1679585382
transform 1 0 142176 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_700
timestamp 1679585382
transform 1 0 142848 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_707
timestamp 1679585382
transform 1 0 143520 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_714
timestamp 1679585382
transform 1 0 144192 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_721
timestamp 1679585382
transform 1 0 144864 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_728
timestamp 1679585382
transform 1 0 145536 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_735
timestamp 1679585382
transform 1 0 146208 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_742
timestamp 1679585382
transform 1 0 146880 0 -1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_31_749
timestamp 1679585382
transform 1 0 147552 0 -1 99792
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_756
timestamp 1677583258
transform 1 0 148224 0 -1 99792
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_0
timestamp 1679585382
transform 1 0 75648 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_7
timestamp 1679585382
transform 1 0 76320 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_14
timestamp 1679585382
transform 1 0 76992 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_21
timestamp 1679585382
transform 1 0 77664 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_28
timestamp 1679585382
transform 1 0 78336 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_35
timestamp 1679585382
transform 1 0 79008 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_42
timestamp 1679585382
transform 1 0 79680 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_49
timestamp 1679585382
transform 1 0 80352 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_56
timestamp 1679585382
transform 1 0 81024 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_63
timestamp 1679585382
transform 1 0 81696 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_70
timestamp 1679585382
transform 1 0 82368 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_77
timestamp 1679585382
transform 1 0 83040 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_84
timestamp 1679585382
transform 1 0 83712 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_91
timestamp 1679585382
transform 1 0 84384 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_98
timestamp 1679585382
transform 1 0 85056 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_105
timestamp 1679585382
transform 1 0 85728 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_112
timestamp 1679585382
transform 1 0 86400 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_119
timestamp 1679585382
transform 1 0 87072 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_126
timestamp 1679585382
transform 1 0 87744 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_133
timestamp 1679585382
transform 1 0 88416 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_140
timestamp 1679585382
transform 1 0 89088 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_147
timestamp 1679585382
transform 1 0 89760 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_154
timestamp 1679585382
transform 1 0 90432 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_161
timestamp 1679585382
transform 1 0 91104 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_168
timestamp 1679585382
transform 1 0 91776 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_175
timestamp 1679585382
transform 1 0 92448 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_182
timestamp 1679585382
transform 1 0 93120 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_189
timestamp 1679585382
transform 1 0 93792 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_196
timestamp 1679585382
transform 1 0 94464 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_203
timestamp 1679585382
transform 1 0 95136 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_210
timestamp 1679585382
transform 1 0 95808 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_217
timestamp 1679585382
transform 1 0 96480 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_224
timestamp 1679585382
transform 1 0 97152 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_231
timestamp 1679585382
transform 1 0 97824 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_238
timestamp 1679585382
transform 1 0 98496 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_245
timestamp 1679585382
transform 1 0 99168 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_252
timestamp 1679585382
transform 1 0 99840 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_259
timestamp 1679585382
transform 1 0 100512 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_266
timestamp 1679585382
transform 1 0 101184 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_273
timestamp 1679585382
transform 1 0 101856 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_280
timestamp 1679585382
transform 1 0 102528 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_287
timestamp 1679585382
transform 1 0 103200 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_294
timestamp 1679585382
transform 1 0 103872 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_301
timestamp 1679585382
transform 1 0 104544 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_308
timestamp 1679585382
transform 1 0 105216 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_315
timestamp 1679585382
transform 1 0 105888 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_322
timestamp 1679585382
transform 1 0 106560 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_329
timestamp 1679585382
transform 1 0 107232 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_336
timestamp 1679585382
transform 1 0 107904 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_343
timestamp 1679585382
transform 1 0 108576 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_350
timestamp 1679585382
transform 1 0 109248 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_357
timestamp 1679585382
transform 1 0 109920 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_364
timestamp 1679585382
transform 1 0 110592 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_371
timestamp 1679585382
transform 1 0 111264 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_378
timestamp 1679585382
transform 1 0 111936 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_385
timestamp 1679585382
transform 1 0 112608 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_392
timestamp 1679585382
transform 1 0 113280 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_399
timestamp 1679585382
transform 1 0 113952 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_406
timestamp 1679585382
transform 1 0 114624 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_413
timestamp 1679585382
transform 1 0 115296 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_420
timestamp 1679585382
transform 1 0 115968 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_427
timestamp 1679585382
transform 1 0 116640 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_434
timestamp 1679585382
transform 1 0 117312 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_441
timestamp 1679585382
transform 1 0 117984 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_448
timestamp 1679585382
transform 1 0 118656 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_455
timestamp 1679585382
transform 1 0 119328 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_462
timestamp 1679585382
transform 1 0 120000 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_469
timestamp 1679585382
transform 1 0 120672 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_476
timestamp 1679585382
transform 1 0 121344 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_483
timestamp 1679585382
transform 1 0 122016 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_490
timestamp 1679585382
transform 1 0 122688 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_497
timestamp 1679585382
transform 1 0 123360 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_504
timestamp 1679585382
transform 1 0 124032 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_511
timestamp 1679585382
transform 1 0 124704 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_518
timestamp 1679585382
transform 1 0 125376 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_525
timestamp 1679585382
transform 1 0 126048 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_532
timestamp 1679585382
transform 1 0 126720 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_539
timestamp 1679585382
transform 1 0 127392 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_546
timestamp 1679585382
transform 1 0 128064 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_553
timestamp 1679585382
transform 1 0 128736 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_560
timestamp 1679585382
transform 1 0 129408 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_567
timestamp 1679585382
transform 1 0 130080 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_574
timestamp 1679585382
transform 1 0 130752 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_581
timestamp 1679585382
transform 1 0 131424 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_588
timestamp 1679585382
transform 1 0 132096 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_595
timestamp 1679585382
transform 1 0 132768 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_602
timestamp 1679585382
transform 1 0 133440 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_609
timestamp 1679585382
transform 1 0 134112 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_616
timestamp 1679585382
transform 1 0 134784 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_623
timestamp 1679585382
transform 1 0 135456 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_630
timestamp 1679585382
transform 1 0 136128 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_637
timestamp 1679585382
transform 1 0 136800 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_644
timestamp 1679585382
transform 1 0 137472 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_651
timestamp 1679585382
transform 1 0 138144 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_658
timestamp 1679585382
transform 1 0 138816 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_665
timestamp 1679585382
transform 1 0 139488 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_672
timestamp 1679585382
transform 1 0 140160 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_679
timestamp 1679585382
transform 1 0 140832 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_686
timestamp 1679585382
transform 1 0 141504 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_693
timestamp 1679585382
transform 1 0 142176 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_700
timestamp 1679585382
transform 1 0 142848 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_707
timestamp 1679585382
transform 1 0 143520 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_714
timestamp 1679585382
transform 1 0 144192 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_721
timestamp 1679585382
transform 1 0 144864 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_728
timestamp 1679585382
transform 1 0 145536 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_735
timestamp 1679585382
transform 1 0 146208 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_742
timestamp 1679585382
transform 1 0 146880 0 1 99792
box -48 -56 720 834
use sg13g2_decap_8  FILLER_32_749
timestamp 1679585382
transform 1 0 147552 0 1 99792
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_756
timestamp 1677583258
transform 1 0 148224 0 1 99792
box -48 -56 144 834
use sg13g2_decap_8  FILLER_33_0
timestamp 1679585382
transform 1 0 75648 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_7
timestamp 1679585382
transform 1 0 76320 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_14
timestamp 1679585382
transform 1 0 76992 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_21
timestamp 1679585382
transform 1 0 77664 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_28
timestamp 1679585382
transform 1 0 78336 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_35
timestamp 1679585382
transform 1 0 79008 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_42
timestamp 1679585382
transform 1 0 79680 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_49
timestamp 1679585382
transform 1 0 80352 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_56
timestamp 1679585382
transform 1 0 81024 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_63
timestamp 1679585382
transform 1 0 81696 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_70
timestamp 1679585382
transform 1 0 82368 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_77
timestamp 1679585382
transform 1 0 83040 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_84
timestamp 1679585382
transform 1 0 83712 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_91
timestamp 1679585382
transform 1 0 84384 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_98
timestamp 1679585382
transform 1 0 85056 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_105
timestamp 1679585382
transform 1 0 85728 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_112
timestamp 1679585382
transform 1 0 86400 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_119
timestamp 1679585382
transform 1 0 87072 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_126
timestamp 1679585382
transform 1 0 87744 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_133
timestamp 1679585382
transform 1 0 88416 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_140
timestamp 1679585382
transform 1 0 89088 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_147
timestamp 1679585382
transform 1 0 89760 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_154
timestamp 1679585382
transform 1 0 90432 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_161
timestamp 1679585382
transform 1 0 91104 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_168
timestamp 1679585382
transform 1 0 91776 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_175
timestamp 1679585382
transform 1 0 92448 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_182
timestamp 1679585382
transform 1 0 93120 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_189
timestamp 1679585382
transform 1 0 93792 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_196
timestamp 1679585382
transform 1 0 94464 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_203
timestamp 1679585382
transform 1 0 95136 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_210
timestamp 1679585382
transform 1 0 95808 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_217
timestamp 1679585382
transform 1 0 96480 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_224
timestamp 1679585382
transform 1 0 97152 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_231
timestamp 1679585382
transform 1 0 97824 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_238
timestamp 1679585382
transform 1 0 98496 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_245
timestamp 1679585382
transform 1 0 99168 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_252
timestamp 1679585382
transform 1 0 99840 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_259
timestamp 1679585382
transform 1 0 100512 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_266
timestamp 1679585382
transform 1 0 101184 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_273
timestamp 1679585382
transform 1 0 101856 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_280
timestamp 1679585382
transform 1 0 102528 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_287
timestamp 1679585382
transform 1 0 103200 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_294
timestamp 1679585382
transform 1 0 103872 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_301
timestamp 1679585382
transform 1 0 104544 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_308
timestamp 1679585382
transform 1 0 105216 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_315
timestamp 1679585382
transform 1 0 105888 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_322
timestamp 1679585382
transform 1 0 106560 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_329
timestamp 1679585382
transform 1 0 107232 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_336
timestamp 1679585382
transform 1 0 107904 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_343
timestamp 1679585382
transform 1 0 108576 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_350
timestamp 1679585382
transform 1 0 109248 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_357
timestamp 1679585382
transform 1 0 109920 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_364
timestamp 1679585382
transform 1 0 110592 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_371
timestamp 1679585382
transform 1 0 111264 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_378
timestamp 1679585382
transform 1 0 111936 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_385
timestamp 1679585382
transform 1 0 112608 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_392
timestamp 1679585382
transform 1 0 113280 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_399
timestamp 1679585382
transform 1 0 113952 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_406
timestamp 1679585382
transform 1 0 114624 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_413
timestamp 1679585382
transform 1 0 115296 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_420
timestamp 1679585382
transform 1 0 115968 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_427
timestamp 1679585382
transform 1 0 116640 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_434
timestamp 1679585382
transform 1 0 117312 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_441
timestamp 1679585382
transform 1 0 117984 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_448
timestamp 1679585382
transform 1 0 118656 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_455
timestamp 1679585382
transform 1 0 119328 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_462
timestamp 1679585382
transform 1 0 120000 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_469
timestamp 1679585382
transform 1 0 120672 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_476
timestamp 1679585382
transform 1 0 121344 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_483
timestamp 1679585382
transform 1 0 122016 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_490
timestamp 1679585382
transform 1 0 122688 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_497
timestamp 1679585382
transform 1 0 123360 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_504
timestamp 1679585382
transform 1 0 124032 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_511
timestamp 1679585382
transform 1 0 124704 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_518
timestamp 1679585382
transform 1 0 125376 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_525
timestamp 1679585382
transform 1 0 126048 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_532
timestamp 1679585382
transform 1 0 126720 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_539
timestamp 1679585382
transform 1 0 127392 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_546
timestamp 1679585382
transform 1 0 128064 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_553
timestamp 1679585382
transform 1 0 128736 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_560
timestamp 1679585382
transform 1 0 129408 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_567
timestamp 1679585382
transform 1 0 130080 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_574
timestamp 1679585382
transform 1 0 130752 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_581
timestamp 1679585382
transform 1 0 131424 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_588
timestamp 1679585382
transform 1 0 132096 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_595
timestamp 1679585382
transform 1 0 132768 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_602
timestamp 1679585382
transform 1 0 133440 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_609
timestamp 1679585382
transform 1 0 134112 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_616
timestamp 1679585382
transform 1 0 134784 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_623
timestamp 1679585382
transform 1 0 135456 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_630
timestamp 1679585382
transform 1 0 136128 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_637
timestamp 1679585382
transform 1 0 136800 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_644
timestamp 1679585382
transform 1 0 137472 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_651
timestamp 1679585382
transform 1 0 138144 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_658
timestamp 1679585382
transform 1 0 138816 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_665
timestamp 1679585382
transform 1 0 139488 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_672
timestamp 1679585382
transform 1 0 140160 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_679
timestamp 1679585382
transform 1 0 140832 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_686
timestamp 1679585382
transform 1 0 141504 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_693
timestamp 1679585382
transform 1 0 142176 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_700
timestamp 1679585382
transform 1 0 142848 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_707
timestamp 1679585382
transform 1 0 143520 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_714
timestamp 1679585382
transform 1 0 144192 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_721
timestamp 1679585382
transform 1 0 144864 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_728
timestamp 1679585382
transform 1 0 145536 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_735
timestamp 1679585382
transform 1 0 146208 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_742
timestamp 1679585382
transform 1 0 146880 0 -1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_749
timestamp 1679585382
transform 1 0 147552 0 -1 101304
box -48 -56 720 834
use sg13g2_fill_1  FILLER_33_756
timestamp 1677583258
transform 1 0 148224 0 -1 101304
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679585382
transform 1 0 75648 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_7
timestamp 1679585382
transform 1 0 76320 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_14
timestamp 1679585382
transform 1 0 76992 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_21
timestamp 1679585382
transform 1 0 77664 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_28
timestamp 1679585382
transform 1 0 78336 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_35
timestamp 1679585382
transform 1 0 79008 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_42
timestamp 1679585382
transform 1 0 79680 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_49
timestamp 1679585382
transform 1 0 80352 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_56
timestamp 1679585382
transform 1 0 81024 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_63
timestamp 1679585382
transform 1 0 81696 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_70
timestamp 1679585382
transform 1 0 82368 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_77
timestamp 1679585382
transform 1 0 83040 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_84
timestamp 1679585382
transform 1 0 83712 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_91
timestamp 1679585382
transform 1 0 84384 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_98
timestamp 1679585382
transform 1 0 85056 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_105
timestamp 1679585382
transform 1 0 85728 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_112
timestamp 1679585382
transform 1 0 86400 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_119
timestamp 1679585382
transform 1 0 87072 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_126
timestamp 1679585382
transform 1 0 87744 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_133
timestamp 1679585382
transform 1 0 88416 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_140
timestamp 1679585382
transform 1 0 89088 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_147
timestamp 1679585382
transform 1 0 89760 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_154
timestamp 1679585382
transform 1 0 90432 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_161
timestamp 1679585382
transform 1 0 91104 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_168
timestamp 1679585382
transform 1 0 91776 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_175
timestamp 1679585382
transform 1 0 92448 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_182
timestamp 1679585382
transform 1 0 93120 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_189
timestamp 1679585382
transform 1 0 93792 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_196
timestamp 1679585382
transform 1 0 94464 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_203
timestamp 1679585382
transform 1 0 95136 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_210
timestamp 1679585382
transform 1 0 95808 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_217
timestamp 1679585382
transform 1 0 96480 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_224
timestamp 1679585382
transform 1 0 97152 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_231
timestamp 1679585382
transform 1 0 97824 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_238
timestamp 1679585382
transform 1 0 98496 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_245
timestamp 1679585382
transform 1 0 99168 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_252
timestamp 1679585382
transform 1 0 99840 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_259
timestamp 1679585382
transform 1 0 100512 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_266
timestamp 1679585382
transform 1 0 101184 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_273
timestamp 1679585382
transform 1 0 101856 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_280
timestamp 1679585382
transform 1 0 102528 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_287
timestamp 1679585382
transform 1 0 103200 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_294
timestamp 1679585382
transform 1 0 103872 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_301
timestamp 1679585382
transform 1 0 104544 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_308
timestamp 1679585382
transform 1 0 105216 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_315
timestamp 1679585382
transform 1 0 105888 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_322
timestamp 1679585382
transform 1 0 106560 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_329
timestamp 1679585382
transform 1 0 107232 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_336
timestamp 1679585382
transform 1 0 107904 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_343
timestamp 1679585382
transform 1 0 108576 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_350
timestamp 1679585382
transform 1 0 109248 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_357
timestamp 1679585382
transform 1 0 109920 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_364
timestamp 1679585382
transform 1 0 110592 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_371
timestamp 1679585382
transform 1 0 111264 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_378
timestamp 1679585382
transform 1 0 111936 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_385
timestamp 1679585382
transform 1 0 112608 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_392
timestamp 1679585382
transform 1 0 113280 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_399
timestamp 1679585382
transform 1 0 113952 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_406
timestamp 1679585382
transform 1 0 114624 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_413
timestamp 1679585382
transform 1 0 115296 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_420
timestamp 1679585382
transform 1 0 115968 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_427
timestamp 1679585382
transform 1 0 116640 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_434
timestamp 1679585382
transform 1 0 117312 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_441
timestamp 1679585382
transform 1 0 117984 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_448
timestamp 1679585382
transform 1 0 118656 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_455
timestamp 1679585382
transform 1 0 119328 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_462
timestamp 1679585382
transform 1 0 120000 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_469
timestamp 1679585382
transform 1 0 120672 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_476
timestamp 1679585382
transform 1 0 121344 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_483
timestamp 1679585382
transform 1 0 122016 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_490
timestamp 1679585382
transform 1 0 122688 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_497
timestamp 1679585382
transform 1 0 123360 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_504
timestamp 1679585382
transform 1 0 124032 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_511
timestamp 1679585382
transform 1 0 124704 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_518
timestamp 1679585382
transform 1 0 125376 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_525
timestamp 1679585382
transform 1 0 126048 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_532
timestamp 1679585382
transform 1 0 126720 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_539
timestamp 1679585382
transform 1 0 127392 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_546
timestamp 1679585382
transform 1 0 128064 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_553
timestamp 1679585382
transform 1 0 128736 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_560
timestamp 1679585382
transform 1 0 129408 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_567
timestamp 1679585382
transform 1 0 130080 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_574
timestamp 1679585382
transform 1 0 130752 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_581
timestamp 1679585382
transform 1 0 131424 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_588
timestamp 1679585382
transform 1 0 132096 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_595
timestamp 1679585382
transform 1 0 132768 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_602
timestamp 1679585382
transform 1 0 133440 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_609
timestamp 1679585382
transform 1 0 134112 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_616
timestamp 1679585382
transform 1 0 134784 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_623
timestamp 1679585382
transform 1 0 135456 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_630
timestamp 1679585382
transform 1 0 136128 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_637
timestamp 1679585382
transform 1 0 136800 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_644
timestamp 1679585382
transform 1 0 137472 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_651
timestamp 1679585382
transform 1 0 138144 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_658
timestamp 1679585382
transform 1 0 138816 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_665
timestamp 1679585382
transform 1 0 139488 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_672
timestamp 1679585382
transform 1 0 140160 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_679
timestamp 1679585382
transform 1 0 140832 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_686
timestamp 1679585382
transform 1 0 141504 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_693
timestamp 1679585382
transform 1 0 142176 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_700
timestamp 1679585382
transform 1 0 142848 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_707
timestamp 1679585382
transform 1 0 143520 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_714
timestamp 1679585382
transform 1 0 144192 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_721
timestamp 1679585382
transform 1 0 144864 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_728
timestamp 1679585382
transform 1 0 145536 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_735
timestamp 1679585382
transform 1 0 146208 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_742
timestamp 1679585382
transform 1 0 146880 0 1 101304
box -48 -56 720 834
use sg13g2_decap_8  FILLER_34_749
timestamp 1679585382
transform 1 0 147552 0 1 101304
box -48 -56 720 834
use sg13g2_fill_1  FILLER_34_756
timestamp 1677583258
transform 1 0 148224 0 1 101304
box -48 -56 144 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679585382
transform 1 0 75648 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679585382
transform 1 0 76320 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_14
timestamp 1679585382
transform 1 0 76992 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_21
timestamp 1679585382
transform 1 0 77664 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_28
timestamp 1679585382
transform 1 0 78336 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_35
timestamp 1679585382
transform 1 0 79008 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_42
timestamp 1679585382
transform 1 0 79680 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_49
timestamp 1679585382
transform 1 0 80352 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_56
timestamp 1679585382
transform 1 0 81024 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_63
timestamp 1679585382
transform 1 0 81696 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_70
timestamp 1679585382
transform 1 0 82368 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_77
timestamp 1679585382
transform 1 0 83040 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_84
timestamp 1679585382
transform 1 0 83712 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_91
timestamp 1679585382
transform 1 0 84384 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_98
timestamp 1679585382
transform 1 0 85056 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_105
timestamp 1679585382
transform 1 0 85728 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_112
timestamp 1679585382
transform 1 0 86400 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_119
timestamp 1679585382
transform 1 0 87072 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_126
timestamp 1679585382
transform 1 0 87744 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_133
timestamp 1679585382
transform 1 0 88416 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_140
timestamp 1679585382
transform 1 0 89088 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_147
timestamp 1679585382
transform 1 0 89760 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_154
timestamp 1679585382
transform 1 0 90432 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_161
timestamp 1679585382
transform 1 0 91104 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_168
timestamp 1679585382
transform 1 0 91776 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_175
timestamp 1679585382
transform 1 0 92448 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_182
timestamp 1679585382
transform 1 0 93120 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_189
timestamp 1679585382
transform 1 0 93792 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_196
timestamp 1679585382
transform 1 0 94464 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_203
timestamp 1679585382
transform 1 0 95136 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_210
timestamp 1679585382
transform 1 0 95808 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_217
timestamp 1679585382
transform 1 0 96480 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_224
timestamp 1679585382
transform 1 0 97152 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_231
timestamp 1679585382
transform 1 0 97824 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_238
timestamp 1679585382
transform 1 0 98496 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_245
timestamp 1679585382
transform 1 0 99168 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_252
timestamp 1679585382
transform 1 0 99840 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_259
timestamp 1679585382
transform 1 0 100512 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_266
timestamp 1679585382
transform 1 0 101184 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_273
timestamp 1679585382
transform 1 0 101856 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_280
timestamp 1679585382
transform 1 0 102528 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_287
timestamp 1679585382
transform 1 0 103200 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_294
timestamp 1679585382
transform 1 0 103872 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_301
timestamp 1679585382
transform 1 0 104544 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_308
timestamp 1679585382
transform 1 0 105216 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_315
timestamp 1679585382
transform 1 0 105888 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_322
timestamp 1679585382
transform 1 0 106560 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_329
timestamp 1679585382
transform 1 0 107232 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_336
timestamp 1679585382
transform 1 0 107904 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_343
timestamp 1679585382
transform 1 0 108576 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_350
timestamp 1679585382
transform 1 0 109248 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_357
timestamp 1679585382
transform 1 0 109920 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_364
timestamp 1679585382
transform 1 0 110592 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_371
timestamp 1679585382
transform 1 0 111264 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_378
timestamp 1679585382
transform 1 0 111936 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_385
timestamp 1679585382
transform 1 0 112608 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_392
timestamp 1679585382
transform 1 0 113280 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_399
timestamp 1679585382
transform 1 0 113952 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_406
timestamp 1679585382
transform 1 0 114624 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_413
timestamp 1679585382
transform 1 0 115296 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_420
timestamp 1679585382
transform 1 0 115968 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_427
timestamp 1679585382
transform 1 0 116640 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_434
timestamp 1679585382
transform 1 0 117312 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_441
timestamp 1679585382
transform 1 0 117984 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_448
timestamp 1679585382
transform 1 0 118656 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_455
timestamp 1679585382
transform 1 0 119328 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_462
timestamp 1679585382
transform 1 0 120000 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_469
timestamp 1679585382
transform 1 0 120672 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_476
timestamp 1679585382
transform 1 0 121344 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_483
timestamp 1679585382
transform 1 0 122016 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_490
timestamp 1679585382
transform 1 0 122688 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_497
timestamp 1679585382
transform 1 0 123360 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_504
timestamp 1679585382
transform 1 0 124032 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_511
timestamp 1679585382
transform 1 0 124704 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_518
timestamp 1679585382
transform 1 0 125376 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_525
timestamp 1679585382
transform 1 0 126048 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_532
timestamp 1679585382
transform 1 0 126720 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_539
timestamp 1679585382
transform 1 0 127392 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_546
timestamp 1679585382
transform 1 0 128064 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_553
timestamp 1679585382
transform 1 0 128736 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_560
timestamp 1679585382
transform 1 0 129408 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_567
timestamp 1679585382
transform 1 0 130080 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_574
timestamp 1679585382
transform 1 0 130752 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_581
timestamp 1679585382
transform 1 0 131424 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_588
timestamp 1679585382
transform 1 0 132096 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_595
timestamp 1679585382
transform 1 0 132768 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_602
timestamp 1679585382
transform 1 0 133440 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_609
timestamp 1679585382
transform 1 0 134112 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_616
timestamp 1679585382
transform 1 0 134784 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_623
timestamp 1679585382
transform 1 0 135456 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_630
timestamp 1679585382
transform 1 0 136128 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_637
timestamp 1679585382
transform 1 0 136800 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_644
timestamp 1679585382
transform 1 0 137472 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_651
timestamp 1679585382
transform 1 0 138144 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_658
timestamp 1679585382
transform 1 0 138816 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_665
timestamp 1679585382
transform 1 0 139488 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_672
timestamp 1679585382
transform 1 0 140160 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_679
timestamp 1679585382
transform 1 0 140832 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_686
timestamp 1679585382
transform 1 0 141504 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_693
timestamp 1679585382
transform 1 0 142176 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_700
timestamp 1679585382
transform 1 0 142848 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_707
timestamp 1679585382
transform 1 0 143520 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_714
timestamp 1679585382
transform 1 0 144192 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_721
timestamp 1679585382
transform 1 0 144864 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_728
timestamp 1679585382
transform 1 0 145536 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_735
timestamp 1679585382
transform 1 0 146208 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_742
timestamp 1679585382
transform 1 0 146880 0 -1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_749
timestamp 1679585382
transform 1 0 147552 0 -1 102816
box -48 -56 720 834
use sg13g2_fill_1  FILLER_35_756
timestamp 1677583258
transform 1 0 148224 0 -1 102816
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679585382
transform 1 0 75648 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679585382
transform 1 0 76320 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_14
timestamp 1679585382
transform 1 0 76992 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_21
timestamp 1679585382
transform 1 0 77664 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_28
timestamp 1679585382
transform 1 0 78336 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_35
timestamp 1679585382
transform 1 0 79008 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_42
timestamp 1679585382
transform 1 0 79680 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_49
timestamp 1679585382
transform 1 0 80352 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_56
timestamp 1679585382
transform 1 0 81024 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_63
timestamp 1679585382
transform 1 0 81696 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_70
timestamp 1679585382
transform 1 0 82368 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_77
timestamp 1679585382
transform 1 0 83040 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_84
timestamp 1679585382
transform 1 0 83712 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_91
timestamp 1679585382
transform 1 0 84384 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_98
timestamp 1679585382
transform 1 0 85056 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_105
timestamp 1679585382
transform 1 0 85728 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_112
timestamp 1679585382
transform 1 0 86400 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_119
timestamp 1679585382
transform 1 0 87072 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_126
timestamp 1679585382
transform 1 0 87744 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_133
timestamp 1679585382
transform 1 0 88416 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_140
timestamp 1679585382
transform 1 0 89088 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_147
timestamp 1679585382
transform 1 0 89760 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_154
timestamp 1679585382
transform 1 0 90432 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_161
timestamp 1679585382
transform 1 0 91104 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_168
timestamp 1679585382
transform 1 0 91776 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_175
timestamp 1679585382
transform 1 0 92448 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_182
timestamp 1679585382
transform 1 0 93120 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_189
timestamp 1679585382
transform 1 0 93792 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_196
timestamp 1679585382
transform 1 0 94464 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_203
timestamp 1679585382
transform 1 0 95136 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_210
timestamp 1679585382
transform 1 0 95808 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_217
timestamp 1679585382
transform 1 0 96480 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_224
timestamp 1679585382
transform 1 0 97152 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_231
timestamp 1679585382
transform 1 0 97824 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_238
timestamp 1679585382
transform 1 0 98496 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_245
timestamp 1679585382
transform 1 0 99168 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_252
timestamp 1679585382
transform 1 0 99840 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_259
timestamp 1679585382
transform 1 0 100512 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_266
timestamp 1679585382
transform 1 0 101184 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_273
timestamp 1679585382
transform 1 0 101856 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_280
timestamp 1679585382
transform 1 0 102528 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_287
timestamp 1679585382
transform 1 0 103200 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_294
timestamp 1679585382
transform 1 0 103872 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_301
timestamp 1679585382
transform 1 0 104544 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_308
timestamp 1679585382
transform 1 0 105216 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_315
timestamp 1679585382
transform 1 0 105888 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_322
timestamp 1679585382
transform 1 0 106560 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_329
timestamp 1679585382
transform 1 0 107232 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_336
timestamp 1679585382
transform 1 0 107904 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_343
timestamp 1679585382
transform 1 0 108576 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_350
timestamp 1679585382
transform 1 0 109248 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_357
timestamp 1679585382
transform 1 0 109920 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_364
timestamp 1679585382
transform 1 0 110592 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_371
timestamp 1679585382
transform 1 0 111264 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_378
timestamp 1679585382
transform 1 0 111936 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_385
timestamp 1679585382
transform 1 0 112608 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_392
timestamp 1679585382
transform 1 0 113280 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_399
timestamp 1679585382
transform 1 0 113952 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_406
timestamp 1679585382
transform 1 0 114624 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_413
timestamp 1679585382
transform 1 0 115296 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_420
timestamp 1679585382
transform 1 0 115968 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_427
timestamp 1679585382
transform 1 0 116640 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_434
timestamp 1679585382
transform 1 0 117312 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_441
timestamp 1679585382
transform 1 0 117984 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_448
timestamp 1679585382
transform 1 0 118656 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_455
timestamp 1679585382
transform 1 0 119328 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_462
timestamp 1679585382
transform 1 0 120000 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_469
timestamp 1679585382
transform 1 0 120672 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_476
timestamp 1679585382
transform 1 0 121344 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_483
timestamp 1679585382
transform 1 0 122016 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_490
timestamp 1679585382
transform 1 0 122688 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_497
timestamp 1679585382
transform 1 0 123360 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_504
timestamp 1679585382
transform 1 0 124032 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_511
timestamp 1679585382
transform 1 0 124704 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_518
timestamp 1679585382
transform 1 0 125376 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_525
timestamp 1679585382
transform 1 0 126048 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_532
timestamp 1679585382
transform 1 0 126720 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_539
timestamp 1679585382
transform 1 0 127392 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_546
timestamp 1679585382
transform 1 0 128064 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_553
timestamp 1679585382
transform 1 0 128736 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_560
timestamp 1679585382
transform 1 0 129408 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_567
timestamp 1679585382
transform 1 0 130080 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_574
timestamp 1679585382
transform 1 0 130752 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_581
timestamp 1679585382
transform 1 0 131424 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_588
timestamp 1679585382
transform 1 0 132096 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_595
timestamp 1679585382
transform 1 0 132768 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_602
timestamp 1679585382
transform 1 0 133440 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_609
timestamp 1679585382
transform 1 0 134112 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_616
timestamp 1679585382
transform 1 0 134784 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_623
timestamp 1679585382
transform 1 0 135456 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_630
timestamp 1679585382
transform 1 0 136128 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_637
timestamp 1679585382
transform 1 0 136800 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_644
timestamp 1679585382
transform 1 0 137472 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_651
timestamp 1679585382
transform 1 0 138144 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_658
timestamp 1679585382
transform 1 0 138816 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_665
timestamp 1679585382
transform 1 0 139488 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_672
timestamp 1679585382
transform 1 0 140160 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_679
timestamp 1679585382
transform 1 0 140832 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_686
timestamp 1679585382
transform 1 0 141504 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_693
timestamp 1679585382
transform 1 0 142176 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_700
timestamp 1679585382
transform 1 0 142848 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_707
timestamp 1679585382
transform 1 0 143520 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_714
timestamp 1679585382
transform 1 0 144192 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_721
timestamp 1679585382
transform 1 0 144864 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_728
timestamp 1679585382
transform 1 0 145536 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_735
timestamp 1679585382
transform 1 0 146208 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_742
timestamp 1679585382
transform 1 0 146880 0 1 102816
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_749
timestamp 1679585382
transform 1 0 147552 0 1 102816
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_756
timestamp 1677583258
transform 1 0 148224 0 1 102816
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_0
timestamp 1679585382
transform 1 0 75648 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_7
timestamp 1679585382
transform 1 0 76320 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_14
timestamp 1679585382
transform 1 0 76992 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_21
timestamp 1679585382
transform 1 0 77664 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_28
timestamp 1679585382
transform 1 0 78336 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_35
timestamp 1679585382
transform 1 0 79008 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_42
timestamp 1679585382
transform 1 0 79680 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_49
timestamp 1679585382
transform 1 0 80352 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_56
timestamp 1679585382
transform 1 0 81024 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_63
timestamp 1679585382
transform 1 0 81696 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_70
timestamp 1679585382
transform 1 0 82368 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_77
timestamp 1679585382
transform 1 0 83040 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_84
timestamp 1679585382
transform 1 0 83712 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_91
timestamp 1679585382
transform 1 0 84384 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_98
timestamp 1679585382
transform 1 0 85056 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_105
timestamp 1679585382
transform 1 0 85728 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_112
timestamp 1679585382
transform 1 0 86400 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_119
timestamp 1679585382
transform 1 0 87072 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_126
timestamp 1679585382
transform 1 0 87744 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_133
timestamp 1679585382
transform 1 0 88416 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_140
timestamp 1679585382
transform 1 0 89088 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_147
timestamp 1679585382
transform 1 0 89760 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_154
timestamp 1679585382
transform 1 0 90432 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_161
timestamp 1679585382
transform 1 0 91104 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_168
timestamp 1679585382
transform 1 0 91776 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_175
timestamp 1679585382
transform 1 0 92448 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_182
timestamp 1679585382
transform 1 0 93120 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_189
timestamp 1679585382
transform 1 0 93792 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_196
timestamp 1679585382
transform 1 0 94464 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_203
timestamp 1679585382
transform 1 0 95136 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_210
timestamp 1679585382
transform 1 0 95808 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_217
timestamp 1679585382
transform 1 0 96480 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_224
timestamp 1679585382
transform 1 0 97152 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_231
timestamp 1679585382
transform 1 0 97824 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_238
timestamp 1679585382
transform 1 0 98496 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_245
timestamp 1679585382
transform 1 0 99168 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_252
timestamp 1679585382
transform 1 0 99840 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_259
timestamp 1679585382
transform 1 0 100512 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_266
timestamp 1679585382
transform 1 0 101184 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_273
timestamp 1679585382
transform 1 0 101856 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_280
timestamp 1679585382
transform 1 0 102528 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_287
timestamp 1679585382
transform 1 0 103200 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_294
timestamp 1679585382
transform 1 0 103872 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_301
timestamp 1679585382
transform 1 0 104544 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_308
timestamp 1679585382
transform 1 0 105216 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_315
timestamp 1679585382
transform 1 0 105888 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_322
timestamp 1679585382
transform 1 0 106560 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_329
timestamp 1679585382
transform 1 0 107232 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_336
timestamp 1679585382
transform 1 0 107904 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_343
timestamp 1679585382
transform 1 0 108576 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_350
timestamp 1679585382
transform 1 0 109248 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_357
timestamp 1679585382
transform 1 0 109920 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_364
timestamp 1679585382
transform 1 0 110592 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_371
timestamp 1679585382
transform 1 0 111264 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_378
timestamp 1679585382
transform 1 0 111936 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_385
timestamp 1679585382
transform 1 0 112608 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_392
timestamp 1679585382
transform 1 0 113280 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_399
timestamp 1679585382
transform 1 0 113952 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_406
timestamp 1679585382
transform 1 0 114624 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_413
timestamp 1679585382
transform 1 0 115296 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_420
timestamp 1679585382
transform 1 0 115968 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_427
timestamp 1679585382
transform 1 0 116640 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_434
timestamp 1679585382
transform 1 0 117312 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_441
timestamp 1679585382
transform 1 0 117984 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_448
timestamp 1679585382
transform 1 0 118656 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_455
timestamp 1679585382
transform 1 0 119328 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_462
timestamp 1679585382
transform 1 0 120000 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_469
timestamp 1679585382
transform 1 0 120672 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_476
timestamp 1679585382
transform 1 0 121344 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_483
timestamp 1679585382
transform 1 0 122016 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_490
timestamp 1679585382
transform 1 0 122688 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_497
timestamp 1679585382
transform 1 0 123360 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_504
timestamp 1679585382
transform 1 0 124032 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_511
timestamp 1679585382
transform 1 0 124704 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_518
timestamp 1679585382
transform 1 0 125376 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_525
timestamp 1679585382
transform 1 0 126048 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_532
timestamp 1679585382
transform 1 0 126720 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_539
timestamp 1679585382
transform 1 0 127392 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_546
timestamp 1679585382
transform 1 0 128064 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_553
timestamp 1679585382
transform 1 0 128736 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_560
timestamp 1679585382
transform 1 0 129408 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_567
timestamp 1679585382
transform 1 0 130080 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_574
timestamp 1679585382
transform 1 0 130752 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_581
timestamp 1679585382
transform 1 0 131424 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_588
timestamp 1679585382
transform 1 0 132096 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_595
timestamp 1679585382
transform 1 0 132768 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_602
timestamp 1679585382
transform 1 0 133440 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_609
timestamp 1679585382
transform 1 0 134112 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_616
timestamp 1679585382
transform 1 0 134784 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_623
timestamp 1679585382
transform 1 0 135456 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_630
timestamp 1679585382
transform 1 0 136128 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_637
timestamp 1679585382
transform 1 0 136800 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_644
timestamp 1679585382
transform 1 0 137472 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_651
timestamp 1679585382
transform 1 0 138144 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_658
timestamp 1679585382
transform 1 0 138816 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_665
timestamp 1679585382
transform 1 0 139488 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_672
timestamp 1679585382
transform 1 0 140160 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_679
timestamp 1679585382
transform 1 0 140832 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_686
timestamp 1679585382
transform 1 0 141504 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_693
timestamp 1679585382
transform 1 0 142176 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_700
timestamp 1679585382
transform 1 0 142848 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_707
timestamp 1679585382
transform 1 0 143520 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_714
timestamp 1679585382
transform 1 0 144192 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_721
timestamp 1679585382
transform 1 0 144864 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_728
timestamp 1679585382
transform 1 0 145536 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_735
timestamp 1679585382
transform 1 0 146208 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_742
timestamp 1679585382
transform 1 0 146880 0 -1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_37_749
timestamp 1679585382
transform 1 0 147552 0 -1 104328
box -48 -56 720 834
use sg13g2_fill_1  FILLER_37_756
timestamp 1677583258
transform 1 0 148224 0 -1 104328
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679585382
transform 1 0 75648 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_7
timestamp 1679585382
transform 1 0 76320 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_14
timestamp 1679585382
transform 1 0 76992 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_21
timestamp 1679585382
transform 1 0 77664 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_28
timestamp 1679585382
transform 1 0 78336 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_35
timestamp 1679585382
transform 1 0 79008 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_42
timestamp 1679585382
transform 1 0 79680 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_49
timestamp 1679585382
transform 1 0 80352 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_56
timestamp 1679585382
transform 1 0 81024 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_63
timestamp 1679585382
transform 1 0 81696 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_70
timestamp 1679585382
transform 1 0 82368 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_77
timestamp 1679585382
transform 1 0 83040 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_84
timestamp 1679585382
transform 1 0 83712 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_91
timestamp 1679585382
transform 1 0 84384 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_98
timestamp 1679585382
transform 1 0 85056 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_105
timestamp 1679585382
transform 1 0 85728 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_112
timestamp 1679585382
transform 1 0 86400 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_119
timestamp 1679585382
transform 1 0 87072 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_126
timestamp 1679585382
transform 1 0 87744 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_133
timestamp 1679585382
transform 1 0 88416 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_140
timestamp 1679585382
transform 1 0 89088 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_147
timestamp 1679585382
transform 1 0 89760 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_154
timestamp 1679585382
transform 1 0 90432 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_161
timestamp 1679585382
transform 1 0 91104 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_168
timestamp 1679585382
transform 1 0 91776 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_175
timestamp 1679585382
transform 1 0 92448 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_182
timestamp 1679585382
transform 1 0 93120 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_189
timestamp 1679585382
transform 1 0 93792 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_196
timestamp 1679585382
transform 1 0 94464 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_203
timestamp 1679585382
transform 1 0 95136 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_210
timestamp 1679585382
transform 1 0 95808 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_217
timestamp 1679585382
transform 1 0 96480 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_224
timestamp 1679585382
transform 1 0 97152 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_231
timestamp 1679585382
transform 1 0 97824 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_238
timestamp 1679585382
transform 1 0 98496 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_245
timestamp 1679585382
transform 1 0 99168 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_252
timestamp 1679585382
transform 1 0 99840 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_259
timestamp 1679585382
transform 1 0 100512 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_266
timestamp 1679585382
transform 1 0 101184 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_273
timestamp 1679585382
transform 1 0 101856 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_280
timestamp 1679585382
transform 1 0 102528 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_287
timestamp 1679585382
transform 1 0 103200 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_294
timestamp 1679585382
transform 1 0 103872 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_301
timestamp 1679585382
transform 1 0 104544 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_308
timestamp 1679585382
transform 1 0 105216 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_315
timestamp 1679585382
transform 1 0 105888 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_322
timestamp 1679585382
transform 1 0 106560 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_329
timestamp 1679585382
transform 1 0 107232 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_336
timestamp 1679585382
transform 1 0 107904 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_343
timestamp 1679585382
transform 1 0 108576 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_350
timestamp 1679585382
transform 1 0 109248 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_357
timestamp 1679585382
transform 1 0 109920 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_364
timestamp 1679585382
transform 1 0 110592 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_371
timestamp 1679585382
transform 1 0 111264 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_378
timestamp 1679585382
transform 1 0 111936 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_385
timestamp 1679585382
transform 1 0 112608 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_392
timestamp 1679585382
transform 1 0 113280 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_399
timestamp 1679585382
transform 1 0 113952 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_406
timestamp 1679585382
transform 1 0 114624 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_413
timestamp 1679585382
transform 1 0 115296 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_420
timestamp 1679585382
transform 1 0 115968 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_427
timestamp 1679585382
transform 1 0 116640 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_434
timestamp 1679585382
transform 1 0 117312 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_441
timestamp 1679585382
transform 1 0 117984 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_448
timestamp 1679585382
transform 1 0 118656 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_455
timestamp 1679585382
transform 1 0 119328 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_462
timestamp 1679585382
transform 1 0 120000 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_469
timestamp 1679585382
transform 1 0 120672 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_476
timestamp 1679585382
transform 1 0 121344 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_483
timestamp 1679585382
transform 1 0 122016 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_490
timestamp 1679585382
transform 1 0 122688 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_497
timestamp 1679585382
transform 1 0 123360 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_504
timestamp 1679585382
transform 1 0 124032 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_511
timestamp 1679585382
transform 1 0 124704 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_518
timestamp 1679585382
transform 1 0 125376 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_525
timestamp 1679585382
transform 1 0 126048 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_532
timestamp 1679585382
transform 1 0 126720 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_539
timestamp 1679585382
transform 1 0 127392 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_546
timestamp 1679585382
transform 1 0 128064 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_553
timestamp 1679585382
transform 1 0 128736 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_560
timestamp 1679585382
transform 1 0 129408 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_567
timestamp 1679585382
transform 1 0 130080 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_574
timestamp 1679585382
transform 1 0 130752 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_581
timestamp 1679585382
transform 1 0 131424 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_588
timestamp 1679585382
transform 1 0 132096 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_595
timestamp 1679585382
transform 1 0 132768 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_602
timestamp 1679585382
transform 1 0 133440 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_609
timestamp 1679585382
transform 1 0 134112 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_616
timestamp 1679585382
transform 1 0 134784 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_623
timestamp 1679585382
transform 1 0 135456 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_630
timestamp 1679585382
transform 1 0 136128 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_637
timestamp 1679585382
transform 1 0 136800 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_644
timestamp 1679585382
transform 1 0 137472 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_651
timestamp 1679585382
transform 1 0 138144 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_658
timestamp 1679585382
transform 1 0 138816 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_665
timestamp 1679585382
transform 1 0 139488 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_672
timestamp 1679585382
transform 1 0 140160 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_679
timestamp 1679585382
transform 1 0 140832 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_686
timestamp 1679585382
transform 1 0 141504 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_693
timestamp 1679585382
transform 1 0 142176 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_700
timestamp 1679585382
transform 1 0 142848 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_707
timestamp 1679585382
transform 1 0 143520 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_714
timestamp 1679585382
transform 1 0 144192 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_721
timestamp 1679585382
transform 1 0 144864 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_728
timestamp 1679585382
transform 1 0 145536 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_735
timestamp 1679585382
transform 1 0 146208 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_742
timestamp 1679585382
transform 1 0 146880 0 1 104328
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_749
timestamp 1679585382
transform 1 0 147552 0 1 104328
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_756
timestamp 1677583258
transform 1 0 148224 0 1 104328
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_0
timestamp 1679585382
transform 1 0 75648 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_7
timestamp 1679585382
transform 1 0 76320 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_14
timestamp 1679585382
transform 1 0 76992 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_21
timestamp 1679585382
transform 1 0 77664 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_28
timestamp 1679585382
transform 1 0 78336 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_35
timestamp 1679585382
transform 1 0 79008 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_42
timestamp 1679585382
transform 1 0 79680 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_49
timestamp 1679585382
transform 1 0 80352 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_56
timestamp 1679585382
transform 1 0 81024 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_63
timestamp 1679585382
transform 1 0 81696 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_70
timestamp 1679585382
transform 1 0 82368 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_77
timestamp 1679585382
transform 1 0 83040 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_84
timestamp 1679585382
transform 1 0 83712 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_91
timestamp 1679585382
transform 1 0 84384 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_98
timestamp 1679585382
transform 1 0 85056 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_105
timestamp 1679585382
transform 1 0 85728 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_112
timestamp 1679585382
transform 1 0 86400 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_119
timestamp 1679585382
transform 1 0 87072 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_126
timestamp 1679585382
transform 1 0 87744 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_133
timestamp 1679585382
transform 1 0 88416 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_140
timestamp 1679585382
transform 1 0 89088 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_147
timestamp 1679585382
transform 1 0 89760 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_154
timestamp 1679585382
transform 1 0 90432 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_161
timestamp 1679585382
transform 1 0 91104 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_168
timestamp 1679585382
transform 1 0 91776 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_175
timestamp 1679585382
transform 1 0 92448 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_182
timestamp 1679585382
transform 1 0 93120 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_189
timestamp 1679585382
transform 1 0 93792 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_196
timestamp 1679585382
transform 1 0 94464 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_203
timestamp 1679585382
transform 1 0 95136 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_210
timestamp 1679585382
transform 1 0 95808 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_217
timestamp 1679585382
transform 1 0 96480 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_224
timestamp 1679585382
transform 1 0 97152 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_231
timestamp 1679585382
transform 1 0 97824 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_238
timestamp 1679585382
transform 1 0 98496 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_245
timestamp 1679585382
transform 1 0 99168 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_252
timestamp 1679585382
transform 1 0 99840 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_259
timestamp 1679585382
transform 1 0 100512 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_266
timestamp 1679585382
transform 1 0 101184 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_273
timestamp 1679585382
transform 1 0 101856 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_280
timestamp 1679585382
transform 1 0 102528 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_287
timestamp 1679585382
transform 1 0 103200 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_294
timestamp 1679585382
transform 1 0 103872 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_301
timestamp 1679585382
transform 1 0 104544 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_308
timestamp 1679585382
transform 1 0 105216 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_315
timestamp 1679585382
transform 1 0 105888 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_322
timestamp 1679585382
transform 1 0 106560 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_329
timestamp 1679585382
transform 1 0 107232 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_336
timestamp 1679585382
transform 1 0 107904 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_343
timestamp 1679585382
transform 1 0 108576 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_350
timestamp 1679585382
transform 1 0 109248 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_357
timestamp 1679585382
transform 1 0 109920 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_364
timestamp 1679585382
transform 1 0 110592 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_371
timestamp 1679585382
transform 1 0 111264 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_378
timestamp 1679585382
transform 1 0 111936 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_385
timestamp 1679585382
transform 1 0 112608 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_392
timestamp 1679585382
transform 1 0 113280 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_399
timestamp 1679585382
transform 1 0 113952 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_406
timestamp 1679585382
transform 1 0 114624 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_413
timestamp 1679585382
transform 1 0 115296 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_420
timestamp 1679585382
transform 1 0 115968 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_427
timestamp 1679585382
transform 1 0 116640 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_434
timestamp 1679585382
transform 1 0 117312 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_441
timestamp 1679585382
transform 1 0 117984 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_448
timestamp 1679585382
transform 1 0 118656 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_455
timestamp 1679585382
transform 1 0 119328 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_462
timestamp 1679585382
transform 1 0 120000 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_469
timestamp 1679585382
transform 1 0 120672 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_476
timestamp 1679585382
transform 1 0 121344 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_483
timestamp 1679585382
transform 1 0 122016 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_490
timestamp 1679585382
transform 1 0 122688 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_497
timestamp 1679585382
transform 1 0 123360 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_504
timestamp 1679585382
transform 1 0 124032 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_511
timestamp 1679585382
transform 1 0 124704 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_518
timestamp 1679585382
transform 1 0 125376 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_525
timestamp 1679585382
transform 1 0 126048 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_532
timestamp 1679585382
transform 1 0 126720 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_539
timestamp 1679585382
transform 1 0 127392 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_546
timestamp 1679585382
transform 1 0 128064 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_553
timestamp 1679585382
transform 1 0 128736 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_560
timestamp 1679585382
transform 1 0 129408 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_567
timestamp 1679585382
transform 1 0 130080 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_574
timestamp 1679585382
transform 1 0 130752 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_581
timestamp 1679585382
transform 1 0 131424 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_588
timestamp 1679585382
transform 1 0 132096 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_595
timestamp 1679585382
transform 1 0 132768 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_602
timestamp 1679585382
transform 1 0 133440 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_609
timestamp 1679585382
transform 1 0 134112 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_616
timestamp 1679585382
transform 1 0 134784 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_623
timestamp 1679585382
transform 1 0 135456 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_630
timestamp 1679585382
transform 1 0 136128 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_637
timestamp 1679585382
transform 1 0 136800 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_644
timestamp 1679585382
transform 1 0 137472 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_651
timestamp 1679585382
transform 1 0 138144 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_658
timestamp 1679585382
transform 1 0 138816 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_665
timestamp 1679585382
transform 1 0 139488 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_672
timestamp 1679585382
transform 1 0 140160 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_679
timestamp 1679585382
transform 1 0 140832 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_686
timestamp 1679585382
transform 1 0 141504 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_693
timestamp 1679585382
transform 1 0 142176 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_700
timestamp 1679585382
transform 1 0 142848 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_707
timestamp 1679585382
transform 1 0 143520 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_714
timestamp 1679585382
transform 1 0 144192 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_721
timestamp 1679585382
transform 1 0 144864 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_728
timestamp 1679585382
transform 1 0 145536 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_735
timestamp 1679585382
transform 1 0 146208 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_742
timestamp 1679585382
transform 1 0 146880 0 -1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_39_749
timestamp 1679585382
transform 1 0 147552 0 -1 105840
box -48 -56 720 834
use sg13g2_fill_1  FILLER_39_756
timestamp 1677583258
transform 1 0 148224 0 -1 105840
box -48 -56 144 834
use sg13g2_decap_8  FILLER_40_0
timestamp 1679585382
transform 1 0 75648 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_7
timestamp 1679585382
transform 1 0 76320 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_14
timestamp 1679585382
transform 1 0 76992 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_21
timestamp 1679585382
transform 1 0 77664 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_28
timestamp 1679585382
transform 1 0 78336 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_35
timestamp 1679585382
transform 1 0 79008 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_42
timestamp 1679585382
transform 1 0 79680 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_49
timestamp 1679585382
transform 1 0 80352 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_56
timestamp 1679585382
transform 1 0 81024 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_63
timestamp 1679585382
transform 1 0 81696 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_70
timestamp 1679585382
transform 1 0 82368 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_77
timestamp 1679585382
transform 1 0 83040 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_84
timestamp 1679585382
transform 1 0 83712 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_91
timestamp 1679585382
transform 1 0 84384 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_98
timestamp 1679585382
transform 1 0 85056 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_105
timestamp 1679585382
transform 1 0 85728 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_112
timestamp 1679585382
transform 1 0 86400 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_119
timestamp 1679585382
transform 1 0 87072 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_126
timestamp 1679585382
transform 1 0 87744 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_133
timestamp 1679585382
transform 1 0 88416 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_140
timestamp 1679585382
transform 1 0 89088 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_147
timestamp 1679585382
transform 1 0 89760 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_154
timestamp 1679585382
transform 1 0 90432 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_161
timestamp 1679585382
transform 1 0 91104 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_168
timestamp 1679585382
transform 1 0 91776 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_175
timestamp 1679585382
transform 1 0 92448 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_182
timestamp 1679585382
transform 1 0 93120 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_189
timestamp 1679585382
transform 1 0 93792 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_196
timestamp 1679585382
transform 1 0 94464 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_203
timestamp 1679585382
transform 1 0 95136 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_210
timestamp 1679585382
transform 1 0 95808 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_217
timestamp 1679585382
transform 1 0 96480 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_224
timestamp 1679585382
transform 1 0 97152 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_231
timestamp 1679585382
transform 1 0 97824 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_238
timestamp 1679585382
transform 1 0 98496 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_245
timestamp 1679585382
transform 1 0 99168 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_252
timestamp 1679585382
transform 1 0 99840 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_259
timestamp 1679585382
transform 1 0 100512 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_266
timestamp 1679585382
transform 1 0 101184 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_273
timestamp 1679585382
transform 1 0 101856 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_280
timestamp 1679585382
transform 1 0 102528 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_287
timestamp 1679585382
transform 1 0 103200 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_294
timestamp 1679585382
transform 1 0 103872 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_301
timestamp 1679585382
transform 1 0 104544 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_308
timestamp 1679585382
transform 1 0 105216 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_315
timestamp 1679585382
transform 1 0 105888 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_322
timestamp 1679585382
transform 1 0 106560 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_329
timestamp 1679585382
transform 1 0 107232 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_336
timestamp 1679585382
transform 1 0 107904 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_343
timestamp 1679585382
transform 1 0 108576 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_350
timestamp 1679585382
transform 1 0 109248 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_357
timestamp 1679585382
transform 1 0 109920 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_364
timestamp 1679585382
transform 1 0 110592 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_371
timestamp 1679585382
transform 1 0 111264 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_378
timestamp 1679585382
transform 1 0 111936 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_385
timestamp 1679585382
transform 1 0 112608 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_392
timestamp 1679585382
transform 1 0 113280 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_399
timestamp 1679585382
transform 1 0 113952 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_406
timestamp 1679585382
transform 1 0 114624 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_413
timestamp 1679585382
transform 1 0 115296 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_420
timestamp 1679585382
transform 1 0 115968 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_427
timestamp 1679585382
transform 1 0 116640 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_434
timestamp 1679585382
transform 1 0 117312 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_441
timestamp 1679585382
transform 1 0 117984 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_448
timestamp 1679585382
transform 1 0 118656 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_455
timestamp 1679585382
transform 1 0 119328 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_462
timestamp 1679585382
transform 1 0 120000 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_469
timestamp 1679585382
transform 1 0 120672 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_476
timestamp 1679585382
transform 1 0 121344 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_483
timestamp 1679585382
transform 1 0 122016 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_490
timestamp 1679585382
transform 1 0 122688 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_497
timestamp 1679585382
transform 1 0 123360 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_504
timestamp 1679585382
transform 1 0 124032 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_511
timestamp 1679585382
transform 1 0 124704 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_518
timestamp 1679585382
transform 1 0 125376 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_525
timestamp 1679585382
transform 1 0 126048 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_532
timestamp 1679585382
transform 1 0 126720 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_539
timestamp 1679585382
transform 1 0 127392 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_546
timestamp 1679585382
transform 1 0 128064 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_553
timestamp 1679585382
transform 1 0 128736 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_560
timestamp 1679585382
transform 1 0 129408 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_567
timestamp 1679585382
transform 1 0 130080 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_574
timestamp 1679585382
transform 1 0 130752 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_581
timestamp 1679585382
transform 1 0 131424 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_588
timestamp 1679585382
transform 1 0 132096 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_595
timestamp 1679585382
transform 1 0 132768 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_602
timestamp 1679585382
transform 1 0 133440 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_609
timestamp 1679585382
transform 1 0 134112 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_616
timestamp 1679585382
transform 1 0 134784 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_623
timestamp 1679585382
transform 1 0 135456 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_630
timestamp 1679585382
transform 1 0 136128 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_637
timestamp 1679585382
transform 1 0 136800 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_644
timestamp 1679585382
transform 1 0 137472 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_651
timestamp 1679585382
transform 1 0 138144 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_658
timestamp 1679585382
transform 1 0 138816 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_665
timestamp 1679585382
transform 1 0 139488 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_672
timestamp 1679585382
transform 1 0 140160 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_679
timestamp 1679585382
transform 1 0 140832 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_686
timestamp 1679585382
transform 1 0 141504 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_693
timestamp 1679585382
transform 1 0 142176 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_700
timestamp 1679585382
transform 1 0 142848 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_707
timestamp 1679585382
transform 1 0 143520 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_714
timestamp 1679585382
transform 1 0 144192 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_721
timestamp 1679585382
transform 1 0 144864 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_728
timestamp 1679585382
transform 1 0 145536 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_735
timestamp 1679585382
transform 1 0 146208 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_742
timestamp 1679585382
transform 1 0 146880 0 1 105840
box -48 -56 720 834
use sg13g2_decap_8  FILLER_40_749
timestamp 1679585382
transform 1 0 147552 0 1 105840
box -48 -56 720 834
use sg13g2_fill_1  FILLER_40_756
timestamp 1677583258
transform 1 0 148224 0 1 105840
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679585382
transform 1 0 75648 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_7
timestamp 1679585382
transform 1 0 76320 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_14
timestamp 1679585382
transform 1 0 76992 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_21
timestamp 1679585382
transform 1 0 77664 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679585382
transform 1 0 78336 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679585382
transform 1 0 79008 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_42
timestamp 1679585382
transform 1 0 79680 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_49
timestamp 1679585382
transform 1 0 80352 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_56
timestamp 1679585382
transform 1 0 81024 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_63
timestamp 1679585382
transform 1 0 81696 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_70
timestamp 1679585382
transform 1 0 82368 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_77
timestamp 1679585382
transform 1 0 83040 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_84
timestamp 1679585382
transform 1 0 83712 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_91
timestamp 1679585382
transform 1 0 84384 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_98
timestamp 1679585382
transform 1 0 85056 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_105
timestamp 1679585382
transform 1 0 85728 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_112
timestamp 1679585382
transform 1 0 86400 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_119
timestamp 1679585382
transform 1 0 87072 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_126
timestamp 1679585382
transform 1 0 87744 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_133
timestamp 1679585382
transform 1 0 88416 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_140
timestamp 1679585382
transform 1 0 89088 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_147
timestamp 1679585382
transform 1 0 89760 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_154
timestamp 1679585382
transform 1 0 90432 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679585382
transform 1 0 91104 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_168
timestamp 1679585382
transform 1 0 91776 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_175
timestamp 1679585382
transform 1 0 92448 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_182
timestamp 1679585382
transform 1 0 93120 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_189
timestamp 1679585382
transform 1 0 93792 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_196
timestamp 1679585382
transform 1 0 94464 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_203
timestamp 1679585382
transform 1 0 95136 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_210
timestamp 1679585382
transform 1 0 95808 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_217
timestamp 1679585382
transform 1 0 96480 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_224
timestamp 1679585382
transform 1 0 97152 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_231
timestamp 1679585382
transform 1 0 97824 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_238
timestamp 1679585382
transform 1 0 98496 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_245
timestamp 1679585382
transform 1 0 99168 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_252
timestamp 1679585382
transform 1 0 99840 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_259
timestamp 1679585382
transform 1 0 100512 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_266
timestamp 1679585382
transform 1 0 101184 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_273
timestamp 1679585382
transform 1 0 101856 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_280
timestamp 1679585382
transform 1 0 102528 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_287
timestamp 1679585382
transform 1 0 103200 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_294
timestamp 1679585382
transform 1 0 103872 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_301
timestamp 1679585382
transform 1 0 104544 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_308
timestamp 1679585382
transform 1 0 105216 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_315
timestamp 1679585382
transform 1 0 105888 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_322
timestamp 1679585382
transform 1 0 106560 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_329
timestamp 1679585382
transform 1 0 107232 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_336
timestamp 1679585382
transform 1 0 107904 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_343
timestamp 1679585382
transform 1 0 108576 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_350
timestamp 1679585382
transform 1 0 109248 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_357
timestamp 1679585382
transform 1 0 109920 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_364
timestamp 1679585382
transform 1 0 110592 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_371
timestamp 1679585382
transform 1 0 111264 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_378
timestamp 1679585382
transform 1 0 111936 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_385
timestamp 1679585382
transform 1 0 112608 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_392
timestamp 1679585382
transform 1 0 113280 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_399
timestamp 1679585382
transform 1 0 113952 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_406
timestamp 1679585382
transform 1 0 114624 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_413
timestamp 1679585382
transform 1 0 115296 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_420
timestamp 1679585382
transform 1 0 115968 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_427
timestamp 1679585382
transform 1 0 116640 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_434
timestamp 1679585382
transform 1 0 117312 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_441
timestamp 1679585382
transform 1 0 117984 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_448
timestamp 1679585382
transform 1 0 118656 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_455
timestamp 1679585382
transform 1 0 119328 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_462
timestamp 1679585382
transform 1 0 120000 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_469
timestamp 1679585382
transform 1 0 120672 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_476
timestamp 1679585382
transform 1 0 121344 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_483
timestamp 1679585382
transform 1 0 122016 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_490
timestamp 1679585382
transform 1 0 122688 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_497
timestamp 1679585382
transform 1 0 123360 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_504
timestamp 1679585382
transform 1 0 124032 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_511
timestamp 1679585382
transform 1 0 124704 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_518
timestamp 1679585382
transform 1 0 125376 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_525
timestamp 1679585382
transform 1 0 126048 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_532
timestamp 1679585382
transform 1 0 126720 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_539
timestamp 1679585382
transform 1 0 127392 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_546
timestamp 1679585382
transform 1 0 128064 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_553
timestamp 1679585382
transform 1 0 128736 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_560
timestamp 1679585382
transform 1 0 129408 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_567
timestamp 1679585382
transform 1 0 130080 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_574
timestamp 1679585382
transform 1 0 130752 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_581
timestamp 1679585382
transform 1 0 131424 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_588
timestamp 1679585382
transform 1 0 132096 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_595
timestamp 1679585382
transform 1 0 132768 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_602
timestamp 1679585382
transform 1 0 133440 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_609
timestamp 1679585382
transform 1 0 134112 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_616
timestamp 1679585382
transform 1 0 134784 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_623
timestamp 1679585382
transform 1 0 135456 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_630
timestamp 1679585382
transform 1 0 136128 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_637
timestamp 1679585382
transform 1 0 136800 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_644
timestamp 1679585382
transform 1 0 137472 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_651
timestamp 1679585382
transform 1 0 138144 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_658
timestamp 1679585382
transform 1 0 138816 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_665
timestamp 1679585382
transform 1 0 139488 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_672
timestamp 1679585382
transform 1 0 140160 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_679
timestamp 1679585382
transform 1 0 140832 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_686
timestamp 1679585382
transform 1 0 141504 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_693
timestamp 1679585382
transform 1 0 142176 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_700
timestamp 1679585382
transform 1 0 142848 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_707
timestamp 1679585382
transform 1 0 143520 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_714
timestamp 1679585382
transform 1 0 144192 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_721
timestamp 1679585382
transform 1 0 144864 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_728
timestamp 1679585382
transform 1 0 145536 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_735
timestamp 1679585382
transform 1 0 146208 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_742
timestamp 1679585382
transform 1 0 146880 0 -1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_749
timestamp 1679585382
transform 1 0 147552 0 -1 107352
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_756
timestamp 1677583258
transform 1 0 148224 0 -1 107352
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_0
timestamp 1679585382
transform 1 0 75648 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_7
timestamp 1679585382
transform 1 0 76320 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_14
timestamp 1679585382
transform 1 0 76992 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_21
timestamp 1679585382
transform 1 0 77664 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_28
timestamp 1679585382
transform 1 0 78336 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_35
timestamp 1679585382
transform 1 0 79008 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_42
timestamp 1679585382
transform 1 0 79680 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_49
timestamp 1679585382
transform 1 0 80352 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_56
timestamp 1679585382
transform 1 0 81024 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_63
timestamp 1679585382
transform 1 0 81696 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_70
timestamp 1679585382
transform 1 0 82368 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_77
timestamp 1679585382
transform 1 0 83040 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_84
timestamp 1679585382
transform 1 0 83712 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_91
timestamp 1679585382
transform 1 0 84384 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_98
timestamp 1679585382
transform 1 0 85056 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_105
timestamp 1679585382
transform 1 0 85728 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_112
timestamp 1679585382
transform 1 0 86400 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_119
timestamp 1679585382
transform 1 0 87072 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_126
timestamp 1679585382
transform 1 0 87744 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_133
timestamp 1679585382
transform 1 0 88416 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_140
timestamp 1679585382
transform 1 0 89088 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_147
timestamp 1679585382
transform 1 0 89760 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_154
timestamp 1679585382
transform 1 0 90432 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_161
timestamp 1679585382
transform 1 0 91104 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_168
timestamp 1679585382
transform 1 0 91776 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_175
timestamp 1679585382
transform 1 0 92448 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_182
timestamp 1679585382
transform 1 0 93120 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_189
timestamp 1679585382
transform 1 0 93792 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_196
timestamp 1679585382
transform 1 0 94464 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_203
timestamp 1679585382
transform 1 0 95136 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_210
timestamp 1679585382
transform 1 0 95808 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_217
timestamp 1679585382
transform 1 0 96480 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_224
timestamp 1679585382
transform 1 0 97152 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_231
timestamp 1679585382
transform 1 0 97824 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_238
timestamp 1679585382
transform 1 0 98496 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_245
timestamp 1679585382
transform 1 0 99168 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_252
timestamp 1679585382
transform 1 0 99840 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_259
timestamp 1679585382
transform 1 0 100512 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_266
timestamp 1679585382
transform 1 0 101184 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_273
timestamp 1679585382
transform 1 0 101856 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_280
timestamp 1679585382
transform 1 0 102528 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_287
timestamp 1679585382
transform 1 0 103200 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_294
timestamp 1679585382
transform 1 0 103872 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_301
timestamp 1679585382
transform 1 0 104544 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_308
timestamp 1679585382
transform 1 0 105216 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_315
timestamp 1679585382
transform 1 0 105888 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_322
timestamp 1679585382
transform 1 0 106560 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_329
timestamp 1679585382
transform 1 0 107232 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_336
timestamp 1679585382
transform 1 0 107904 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_343
timestamp 1679585382
transform 1 0 108576 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_350
timestamp 1679585382
transform 1 0 109248 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_357
timestamp 1679585382
transform 1 0 109920 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_364
timestamp 1679585382
transform 1 0 110592 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_371
timestamp 1679585382
transform 1 0 111264 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_378
timestamp 1679585382
transform 1 0 111936 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_385
timestamp 1679585382
transform 1 0 112608 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_392
timestamp 1679585382
transform 1 0 113280 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_399
timestamp 1679585382
transform 1 0 113952 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_406
timestamp 1679585382
transform 1 0 114624 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_413
timestamp 1679585382
transform 1 0 115296 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_420
timestamp 1679585382
transform 1 0 115968 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_427
timestamp 1679585382
transform 1 0 116640 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_434
timestamp 1679585382
transform 1 0 117312 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_441
timestamp 1679585382
transform 1 0 117984 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_448
timestamp 1679585382
transform 1 0 118656 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_455
timestamp 1679585382
transform 1 0 119328 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_462
timestamp 1679585382
transform 1 0 120000 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_469
timestamp 1679585382
transform 1 0 120672 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_476
timestamp 1679585382
transform 1 0 121344 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_483
timestamp 1679585382
transform 1 0 122016 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_490
timestamp 1679585382
transform 1 0 122688 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_497
timestamp 1679585382
transform 1 0 123360 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_504
timestamp 1679585382
transform 1 0 124032 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_511
timestamp 1679585382
transform 1 0 124704 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_518
timestamp 1679585382
transform 1 0 125376 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_525
timestamp 1679585382
transform 1 0 126048 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_532
timestamp 1679585382
transform 1 0 126720 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_539
timestamp 1679585382
transform 1 0 127392 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_546
timestamp 1679585382
transform 1 0 128064 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_553
timestamp 1679585382
transform 1 0 128736 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_560
timestamp 1679585382
transform 1 0 129408 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_567
timestamp 1679585382
transform 1 0 130080 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_574
timestamp 1679585382
transform 1 0 130752 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_581
timestamp 1679585382
transform 1 0 131424 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_588
timestamp 1679585382
transform 1 0 132096 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_595
timestamp 1679585382
transform 1 0 132768 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_602
timestamp 1679585382
transform 1 0 133440 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_609
timestamp 1679585382
transform 1 0 134112 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_616
timestamp 1679585382
transform 1 0 134784 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_623
timestamp 1679585382
transform 1 0 135456 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_630
timestamp 1679585382
transform 1 0 136128 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_637
timestamp 1679585382
transform 1 0 136800 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_644
timestamp 1679585382
transform 1 0 137472 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_651
timestamp 1679585382
transform 1 0 138144 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_658
timestamp 1679585382
transform 1 0 138816 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_665
timestamp 1679585382
transform 1 0 139488 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_672
timestamp 1679585382
transform 1 0 140160 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_679
timestamp 1679585382
transform 1 0 140832 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_686
timestamp 1679585382
transform 1 0 141504 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_693
timestamp 1679585382
transform 1 0 142176 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_700
timestamp 1679585382
transform 1 0 142848 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_707
timestamp 1679585382
transform 1 0 143520 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_714
timestamp 1679585382
transform 1 0 144192 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_721
timestamp 1679585382
transform 1 0 144864 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_728
timestamp 1679585382
transform 1 0 145536 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_735
timestamp 1679585382
transform 1 0 146208 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_742
timestamp 1679585382
transform 1 0 146880 0 1 107352
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_749
timestamp 1679585382
transform 1 0 147552 0 1 107352
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_756
timestamp 1677583258
transform 1 0 148224 0 1 107352
box -48 -56 144 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679585382
transform 1 0 75648 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_7
timestamp 1679585382
transform 1 0 76320 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_14
timestamp 1679585382
transform 1 0 76992 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_21
timestamp 1679585382
transform 1 0 77664 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_28
timestamp 1679585382
transform 1 0 78336 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_35
timestamp 1679585382
transform 1 0 79008 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_42
timestamp 1679585382
transform 1 0 79680 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_49
timestamp 1679585382
transform 1 0 80352 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_56
timestamp 1679585382
transform 1 0 81024 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_63
timestamp 1679585382
transform 1 0 81696 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_70
timestamp 1679585382
transform 1 0 82368 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_77
timestamp 1679585382
transform 1 0 83040 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_84
timestamp 1679585382
transform 1 0 83712 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_91
timestamp 1679585382
transform 1 0 84384 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_98
timestamp 1679585382
transform 1 0 85056 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_105
timestamp 1679585382
transform 1 0 85728 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_112
timestamp 1679585382
transform 1 0 86400 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_119
timestamp 1679585382
transform 1 0 87072 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_126
timestamp 1679585382
transform 1 0 87744 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_133
timestamp 1679585382
transform 1 0 88416 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_140
timestamp 1679585382
transform 1 0 89088 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_147
timestamp 1679585382
transform 1 0 89760 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_154
timestamp 1679585382
transform 1 0 90432 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_161
timestamp 1679585382
transform 1 0 91104 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_168
timestamp 1679585382
transform 1 0 91776 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_175
timestamp 1679585382
transform 1 0 92448 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_182
timestamp 1679585382
transform 1 0 93120 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_189
timestamp 1679585382
transform 1 0 93792 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_196
timestamp 1679585382
transform 1 0 94464 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_203
timestamp 1679585382
transform 1 0 95136 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_210
timestamp 1679585382
transform 1 0 95808 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_217
timestamp 1679585382
transform 1 0 96480 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_224
timestamp 1679585382
transform 1 0 97152 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_231
timestamp 1679585382
transform 1 0 97824 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_238
timestamp 1679585382
transform 1 0 98496 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_245
timestamp 1679585382
transform 1 0 99168 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_252
timestamp 1679585382
transform 1 0 99840 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_259
timestamp 1679585382
transform 1 0 100512 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_266
timestamp 1679585382
transform 1 0 101184 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_273
timestamp 1679585382
transform 1 0 101856 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_280
timestamp 1679585382
transform 1 0 102528 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_287
timestamp 1679585382
transform 1 0 103200 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_294
timestamp 1679585382
transform 1 0 103872 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_301
timestamp 1679585382
transform 1 0 104544 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_308
timestamp 1679585382
transform 1 0 105216 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_315
timestamp 1679585382
transform 1 0 105888 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_322
timestamp 1679585382
transform 1 0 106560 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_329
timestamp 1679585382
transform 1 0 107232 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_336
timestamp 1679585382
transform 1 0 107904 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_343
timestamp 1679585382
transform 1 0 108576 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_350
timestamp 1679585382
transform 1 0 109248 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_357
timestamp 1679585382
transform 1 0 109920 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_364
timestamp 1679585382
transform 1 0 110592 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_371
timestamp 1679585382
transform 1 0 111264 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_378
timestamp 1679585382
transform 1 0 111936 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_385
timestamp 1679585382
transform 1 0 112608 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_392
timestamp 1679585382
transform 1 0 113280 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_399
timestamp 1679585382
transform 1 0 113952 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_406
timestamp 1679585382
transform 1 0 114624 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_413
timestamp 1679585382
transform 1 0 115296 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_420
timestamp 1679585382
transform 1 0 115968 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_427
timestamp 1679585382
transform 1 0 116640 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_434
timestamp 1679585382
transform 1 0 117312 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_441
timestamp 1679585382
transform 1 0 117984 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_448
timestamp 1679585382
transform 1 0 118656 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_455
timestamp 1679585382
transform 1 0 119328 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_462
timestamp 1679585382
transform 1 0 120000 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_469
timestamp 1679585382
transform 1 0 120672 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_476
timestamp 1679585382
transform 1 0 121344 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_483
timestamp 1679585382
transform 1 0 122016 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_490
timestamp 1679585382
transform 1 0 122688 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_497
timestamp 1679585382
transform 1 0 123360 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_504
timestamp 1679585382
transform 1 0 124032 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_511
timestamp 1679585382
transform 1 0 124704 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_518
timestamp 1679585382
transform 1 0 125376 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_525
timestamp 1679585382
transform 1 0 126048 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_532
timestamp 1679585382
transform 1 0 126720 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_539
timestamp 1679585382
transform 1 0 127392 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_546
timestamp 1679585382
transform 1 0 128064 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_553
timestamp 1679585382
transform 1 0 128736 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_560
timestamp 1679585382
transform 1 0 129408 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_567
timestamp 1679585382
transform 1 0 130080 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_574
timestamp 1679585382
transform 1 0 130752 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_581
timestamp 1679585382
transform 1 0 131424 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_588
timestamp 1679585382
transform 1 0 132096 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_595
timestamp 1679585382
transform 1 0 132768 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_602
timestamp 1679585382
transform 1 0 133440 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_609
timestamp 1679585382
transform 1 0 134112 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_616
timestamp 1679585382
transform 1 0 134784 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_623
timestamp 1679585382
transform 1 0 135456 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_630
timestamp 1679585382
transform 1 0 136128 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_637
timestamp 1679585382
transform 1 0 136800 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_644
timestamp 1679585382
transform 1 0 137472 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_651
timestamp 1679585382
transform 1 0 138144 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_658
timestamp 1679585382
transform 1 0 138816 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_665
timestamp 1679585382
transform 1 0 139488 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_672
timestamp 1679585382
transform 1 0 140160 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_679
timestamp 1679585382
transform 1 0 140832 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_686
timestamp 1679585382
transform 1 0 141504 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_693
timestamp 1679585382
transform 1 0 142176 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_700
timestamp 1679585382
transform 1 0 142848 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_707
timestamp 1679585382
transform 1 0 143520 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_714
timestamp 1679585382
transform 1 0 144192 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_721
timestamp 1679585382
transform 1 0 144864 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_728
timestamp 1679585382
transform 1 0 145536 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_735
timestamp 1679585382
transform 1 0 146208 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_742
timestamp 1679585382
transform 1 0 146880 0 -1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_43_749
timestamp 1679585382
transform 1 0 147552 0 -1 108864
box -48 -56 720 834
use sg13g2_fill_1  FILLER_43_756
timestamp 1677583258
transform 1 0 148224 0 -1 108864
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_0
timestamp 1679585382
transform 1 0 75648 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_7
timestamp 1679585382
transform 1 0 76320 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_14
timestamp 1679585382
transform 1 0 76992 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_21
timestamp 1679585382
transform 1 0 77664 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_28
timestamp 1679585382
transform 1 0 78336 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_35
timestamp 1679585382
transform 1 0 79008 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_42
timestamp 1679585382
transform 1 0 79680 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_49
timestamp 1679585382
transform 1 0 80352 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_56
timestamp 1679585382
transform 1 0 81024 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_63
timestamp 1679585382
transform 1 0 81696 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_70
timestamp 1679585382
transform 1 0 82368 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_77
timestamp 1679585382
transform 1 0 83040 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_84
timestamp 1679585382
transform 1 0 83712 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_91
timestamp 1679585382
transform 1 0 84384 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_98
timestamp 1679585382
transform 1 0 85056 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_105
timestamp 1679585382
transform 1 0 85728 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_112
timestamp 1679585382
transform 1 0 86400 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_119
timestamp 1679585382
transform 1 0 87072 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_126
timestamp 1679585382
transform 1 0 87744 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_133
timestamp 1679585382
transform 1 0 88416 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_140
timestamp 1679585382
transform 1 0 89088 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_147
timestamp 1679585382
transform 1 0 89760 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_154
timestamp 1679585382
transform 1 0 90432 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_161
timestamp 1679585382
transform 1 0 91104 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_168
timestamp 1679585382
transform 1 0 91776 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_175
timestamp 1679585382
transform 1 0 92448 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_182
timestamp 1679585382
transform 1 0 93120 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_189
timestamp 1679585382
transform 1 0 93792 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_196
timestamp 1679585382
transform 1 0 94464 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_203
timestamp 1679585382
transform 1 0 95136 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_210
timestamp 1679585382
transform 1 0 95808 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_217
timestamp 1679585382
transform 1 0 96480 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_224
timestamp 1679585382
transform 1 0 97152 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_231
timestamp 1679585382
transform 1 0 97824 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_238
timestamp 1679585382
transform 1 0 98496 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_245
timestamp 1679585382
transform 1 0 99168 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_252
timestamp 1679585382
transform 1 0 99840 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_259
timestamp 1679585382
transform 1 0 100512 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_266
timestamp 1679585382
transform 1 0 101184 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_273
timestamp 1679585382
transform 1 0 101856 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_280
timestamp 1679585382
transform 1 0 102528 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_287
timestamp 1679585382
transform 1 0 103200 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_294
timestamp 1679585382
transform 1 0 103872 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_301
timestamp 1679585382
transform 1 0 104544 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_308
timestamp 1679585382
transform 1 0 105216 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_315
timestamp 1679585382
transform 1 0 105888 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_322
timestamp 1679585382
transform 1 0 106560 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_329
timestamp 1679585382
transform 1 0 107232 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_336
timestamp 1679585382
transform 1 0 107904 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_343
timestamp 1679585382
transform 1 0 108576 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_350
timestamp 1679585382
transform 1 0 109248 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_357
timestamp 1679585382
transform 1 0 109920 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_364
timestamp 1679585382
transform 1 0 110592 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_371
timestamp 1679585382
transform 1 0 111264 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_378
timestamp 1679585382
transform 1 0 111936 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_385
timestamp 1679585382
transform 1 0 112608 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_392
timestamp 1679585382
transform 1 0 113280 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_399
timestamp 1679585382
transform 1 0 113952 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_406
timestamp 1679585382
transform 1 0 114624 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_413
timestamp 1679585382
transform 1 0 115296 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_420
timestamp 1679585382
transform 1 0 115968 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_427
timestamp 1679585382
transform 1 0 116640 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_434
timestamp 1679585382
transform 1 0 117312 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_441
timestamp 1679585382
transform 1 0 117984 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_448
timestamp 1679585382
transform 1 0 118656 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_455
timestamp 1679585382
transform 1 0 119328 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_462
timestamp 1679585382
transform 1 0 120000 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_469
timestamp 1679585382
transform 1 0 120672 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_476
timestamp 1679585382
transform 1 0 121344 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_483
timestamp 1679585382
transform 1 0 122016 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_490
timestamp 1679585382
transform 1 0 122688 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_497
timestamp 1679585382
transform 1 0 123360 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_504
timestamp 1679585382
transform 1 0 124032 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_511
timestamp 1679585382
transform 1 0 124704 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_518
timestamp 1679585382
transform 1 0 125376 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_525
timestamp 1679585382
transform 1 0 126048 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_532
timestamp 1679585382
transform 1 0 126720 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_539
timestamp 1679585382
transform 1 0 127392 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_546
timestamp 1679585382
transform 1 0 128064 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_553
timestamp 1679585382
transform 1 0 128736 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_560
timestamp 1679585382
transform 1 0 129408 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_567
timestamp 1679585382
transform 1 0 130080 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_574
timestamp 1679585382
transform 1 0 130752 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_581
timestamp 1679585382
transform 1 0 131424 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_588
timestamp 1679585382
transform 1 0 132096 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_595
timestamp 1679585382
transform 1 0 132768 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_602
timestamp 1679585382
transform 1 0 133440 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_609
timestamp 1679585382
transform 1 0 134112 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_616
timestamp 1679585382
transform 1 0 134784 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_623
timestamp 1679585382
transform 1 0 135456 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_630
timestamp 1679585382
transform 1 0 136128 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_637
timestamp 1679585382
transform 1 0 136800 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_644
timestamp 1679585382
transform 1 0 137472 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_651
timestamp 1679585382
transform 1 0 138144 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_658
timestamp 1679585382
transform 1 0 138816 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_665
timestamp 1679585382
transform 1 0 139488 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_672
timestamp 1679585382
transform 1 0 140160 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_679
timestamp 1679585382
transform 1 0 140832 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_686
timestamp 1679585382
transform 1 0 141504 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_693
timestamp 1679585382
transform 1 0 142176 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_700
timestamp 1679585382
transform 1 0 142848 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_707
timestamp 1679585382
transform 1 0 143520 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_714
timestamp 1679585382
transform 1 0 144192 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_721
timestamp 1679585382
transform 1 0 144864 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_728
timestamp 1679585382
transform 1 0 145536 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_735
timestamp 1679585382
transform 1 0 146208 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_742
timestamp 1679585382
transform 1 0 146880 0 1 108864
box -48 -56 720 834
use sg13g2_decap_8  FILLER_44_749
timestamp 1679585382
transform 1 0 147552 0 1 108864
box -48 -56 720 834
use sg13g2_fill_1  FILLER_44_756
timestamp 1677583258
transform 1 0 148224 0 1 108864
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679585382
transform 1 0 75648 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_7
timestamp 1679585382
transform 1 0 76320 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_14
timestamp 1679585382
transform 1 0 76992 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_21
timestamp 1679585382
transform 1 0 77664 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679585382
transform 1 0 78336 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679585382
transform 1 0 79008 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_42
timestamp 1679585382
transform 1 0 79680 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_49
timestamp 1679585382
transform 1 0 80352 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_56
timestamp 1679585382
transform 1 0 81024 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_63
timestamp 1679585382
transform 1 0 81696 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_70
timestamp 1679585382
transform 1 0 82368 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_77
timestamp 1679585382
transform 1 0 83040 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_84
timestamp 1679585382
transform 1 0 83712 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_91
timestamp 1679585382
transform 1 0 84384 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_98
timestamp 1679585382
transform 1 0 85056 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679585382
transform 1 0 85728 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_112
timestamp 1679585382
transform 1 0 86400 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_119
timestamp 1679585382
transform 1 0 87072 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_126
timestamp 1679585382
transform 1 0 87744 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_133
timestamp 1679585382
transform 1 0 88416 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_140
timestamp 1679585382
transform 1 0 89088 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_147
timestamp 1679585382
transform 1 0 89760 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_154
timestamp 1679585382
transform 1 0 90432 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_161
timestamp 1679585382
transform 1 0 91104 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_168
timestamp 1679585382
transform 1 0 91776 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_175
timestamp 1679585382
transform 1 0 92448 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_182
timestamp 1679585382
transform 1 0 93120 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_189
timestamp 1679585382
transform 1 0 93792 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_196
timestamp 1679585382
transform 1 0 94464 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_203
timestamp 1679585382
transform 1 0 95136 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_210
timestamp 1679585382
transform 1 0 95808 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_217
timestamp 1679585382
transform 1 0 96480 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_224
timestamp 1679585382
transform 1 0 97152 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_231
timestamp 1679585382
transform 1 0 97824 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_238
timestamp 1679585382
transform 1 0 98496 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_245
timestamp 1679585382
transform 1 0 99168 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_252
timestamp 1679585382
transform 1 0 99840 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_259
timestamp 1679585382
transform 1 0 100512 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_266
timestamp 1679585382
transform 1 0 101184 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_273
timestamp 1679585382
transform 1 0 101856 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_280
timestamp 1679585382
transform 1 0 102528 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_287
timestamp 1679585382
transform 1 0 103200 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_294
timestamp 1679585382
transform 1 0 103872 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_301
timestamp 1679585382
transform 1 0 104544 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_308
timestamp 1679585382
transform 1 0 105216 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_315
timestamp 1679585382
transform 1 0 105888 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_322
timestamp 1679585382
transform 1 0 106560 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_329
timestamp 1679585382
transform 1 0 107232 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_336
timestamp 1679585382
transform 1 0 107904 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_343
timestamp 1679585382
transform 1 0 108576 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_350
timestamp 1679585382
transform 1 0 109248 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_357
timestamp 1679585382
transform 1 0 109920 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_364
timestamp 1679585382
transform 1 0 110592 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_371
timestamp 1679585382
transform 1 0 111264 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_378
timestamp 1679585382
transform 1 0 111936 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_385
timestamp 1679585382
transform 1 0 112608 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_392
timestamp 1679585382
transform 1 0 113280 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_399
timestamp 1679585382
transform 1 0 113952 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_406
timestamp 1679585382
transform 1 0 114624 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_413
timestamp 1679585382
transform 1 0 115296 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_420
timestamp 1679585382
transform 1 0 115968 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_427
timestamp 1679585382
transform 1 0 116640 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_434
timestamp 1679585382
transform 1 0 117312 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_441
timestamp 1679585382
transform 1 0 117984 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_448
timestamp 1679585382
transform 1 0 118656 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_455
timestamp 1679585382
transform 1 0 119328 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_462
timestamp 1679585382
transform 1 0 120000 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_469
timestamp 1679585382
transform 1 0 120672 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_476
timestamp 1679585382
transform 1 0 121344 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_483
timestamp 1679585382
transform 1 0 122016 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_490
timestamp 1679585382
transform 1 0 122688 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_497
timestamp 1679585382
transform 1 0 123360 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_504
timestamp 1679585382
transform 1 0 124032 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_511
timestamp 1679585382
transform 1 0 124704 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_518
timestamp 1679585382
transform 1 0 125376 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_525
timestamp 1679585382
transform 1 0 126048 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_532
timestamp 1679585382
transform 1 0 126720 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_539
timestamp 1679585382
transform 1 0 127392 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_546
timestamp 1679585382
transform 1 0 128064 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_553
timestamp 1679585382
transform 1 0 128736 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_560
timestamp 1679585382
transform 1 0 129408 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_567
timestamp 1679585382
transform 1 0 130080 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_574
timestamp 1679585382
transform 1 0 130752 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_581
timestamp 1679585382
transform 1 0 131424 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_588
timestamp 1679585382
transform 1 0 132096 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_595
timestamp 1679585382
transform 1 0 132768 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_602
timestamp 1679585382
transform 1 0 133440 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_609
timestamp 1679585382
transform 1 0 134112 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_616
timestamp 1679585382
transform 1 0 134784 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_623
timestamp 1679585382
transform 1 0 135456 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_630
timestamp 1679585382
transform 1 0 136128 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_637
timestamp 1679585382
transform 1 0 136800 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_644
timestamp 1679585382
transform 1 0 137472 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_651
timestamp 1679585382
transform 1 0 138144 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_658
timestamp 1679585382
transform 1 0 138816 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_665
timestamp 1679585382
transform 1 0 139488 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_672
timestamp 1679585382
transform 1 0 140160 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_679
timestamp 1679585382
transform 1 0 140832 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_686
timestamp 1679585382
transform 1 0 141504 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_693
timestamp 1679585382
transform 1 0 142176 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_700
timestamp 1679585382
transform 1 0 142848 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_707
timestamp 1679585382
transform 1 0 143520 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_714
timestamp 1679585382
transform 1 0 144192 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_721
timestamp 1679585382
transform 1 0 144864 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_728
timestamp 1679585382
transform 1 0 145536 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_735
timestamp 1679585382
transform 1 0 146208 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_742
timestamp 1679585382
transform 1 0 146880 0 -1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_749
timestamp 1679585382
transform 1 0 147552 0 -1 110376
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_756
timestamp 1677583258
transform 1 0 148224 0 -1 110376
box -48 -56 144 834
use sg13g2_decap_8  FILLER_46_0
timestamp 1679585382
transform 1 0 75648 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_7
timestamp 1679585382
transform 1 0 76320 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_14
timestamp 1679585382
transform 1 0 76992 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_21
timestamp 1679585382
transform 1 0 77664 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_28
timestamp 1679585382
transform 1 0 78336 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_35
timestamp 1679585382
transform 1 0 79008 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_42
timestamp 1679585382
transform 1 0 79680 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_49
timestamp 1679585382
transform 1 0 80352 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_56
timestamp 1679585382
transform 1 0 81024 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_63
timestamp 1679585382
transform 1 0 81696 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_70
timestamp 1679585382
transform 1 0 82368 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_77
timestamp 1679585382
transform 1 0 83040 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_84
timestamp 1679585382
transform 1 0 83712 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_91
timestamp 1679585382
transform 1 0 84384 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_98
timestamp 1679585382
transform 1 0 85056 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_105
timestamp 1679585382
transform 1 0 85728 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_112
timestamp 1679585382
transform 1 0 86400 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_119
timestamp 1679585382
transform 1 0 87072 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_126
timestamp 1679585382
transform 1 0 87744 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_133
timestamp 1679585382
transform 1 0 88416 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_140
timestamp 1679585382
transform 1 0 89088 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_147
timestamp 1679585382
transform 1 0 89760 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_154
timestamp 1679585382
transform 1 0 90432 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_161
timestamp 1679585382
transform 1 0 91104 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_168
timestamp 1679585382
transform 1 0 91776 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_175
timestamp 1679585382
transform 1 0 92448 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_182
timestamp 1679585382
transform 1 0 93120 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_189
timestamp 1679585382
transform 1 0 93792 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_196
timestamp 1679585382
transform 1 0 94464 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_203
timestamp 1679585382
transform 1 0 95136 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_210
timestamp 1679585382
transform 1 0 95808 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_217
timestamp 1679585382
transform 1 0 96480 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_224
timestamp 1679585382
transform 1 0 97152 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_231
timestamp 1679585382
transform 1 0 97824 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_238
timestamp 1679585382
transform 1 0 98496 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_245
timestamp 1679585382
transform 1 0 99168 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_252
timestamp 1679585382
transform 1 0 99840 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_259
timestamp 1679585382
transform 1 0 100512 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_266
timestamp 1679585382
transform 1 0 101184 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_273
timestamp 1679585382
transform 1 0 101856 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_280
timestamp 1679585382
transform 1 0 102528 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_287
timestamp 1679585382
transform 1 0 103200 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_294
timestamp 1679585382
transform 1 0 103872 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_301
timestamp 1679585382
transform 1 0 104544 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_308
timestamp 1679585382
transform 1 0 105216 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_315
timestamp 1679585382
transform 1 0 105888 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_322
timestamp 1679585382
transform 1 0 106560 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_329
timestamp 1679585382
transform 1 0 107232 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_336
timestamp 1679585382
transform 1 0 107904 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_343
timestamp 1679585382
transform 1 0 108576 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_350
timestamp 1679585382
transform 1 0 109248 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_357
timestamp 1679585382
transform 1 0 109920 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_364
timestamp 1679585382
transform 1 0 110592 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_371
timestamp 1679585382
transform 1 0 111264 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_378
timestamp 1679585382
transform 1 0 111936 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_385
timestamp 1679585382
transform 1 0 112608 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_392
timestamp 1679585382
transform 1 0 113280 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_399
timestamp 1679585382
transform 1 0 113952 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_406
timestamp 1679585382
transform 1 0 114624 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_413
timestamp 1679585382
transform 1 0 115296 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_420
timestamp 1679585382
transform 1 0 115968 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_427
timestamp 1679585382
transform 1 0 116640 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_434
timestamp 1679585382
transform 1 0 117312 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_441
timestamp 1679585382
transform 1 0 117984 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_448
timestamp 1679585382
transform 1 0 118656 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_455
timestamp 1679585382
transform 1 0 119328 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_462
timestamp 1679585382
transform 1 0 120000 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_469
timestamp 1679585382
transform 1 0 120672 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_476
timestamp 1679585382
transform 1 0 121344 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_483
timestamp 1679585382
transform 1 0 122016 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_490
timestamp 1679585382
transform 1 0 122688 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_497
timestamp 1679585382
transform 1 0 123360 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_504
timestamp 1679585382
transform 1 0 124032 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_511
timestamp 1679585382
transform 1 0 124704 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_518
timestamp 1679585382
transform 1 0 125376 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_525
timestamp 1679585382
transform 1 0 126048 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_532
timestamp 1679585382
transform 1 0 126720 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_539
timestamp 1679585382
transform 1 0 127392 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_546
timestamp 1679585382
transform 1 0 128064 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_553
timestamp 1679585382
transform 1 0 128736 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_560
timestamp 1679585382
transform 1 0 129408 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_567
timestamp 1679585382
transform 1 0 130080 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_574
timestamp 1679585382
transform 1 0 130752 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_581
timestamp 1679585382
transform 1 0 131424 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_588
timestamp 1679585382
transform 1 0 132096 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_595
timestamp 1679585382
transform 1 0 132768 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_602
timestamp 1679585382
transform 1 0 133440 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_609
timestamp 1679585382
transform 1 0 134112 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_616
timestamp 1679585382
transform 1 0 134784 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_623
timestamp 1679585382
transform 1 0 135456 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_630
timestamp 1679585382
transform 1 0 136128 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_637
timestamp 1679585382
transform 1 0 136800 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_644
timestamp 1679585382
transform 1 0 137472 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_651
timestamp 1679585382
transform 1 0 138144 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_658
timestamp 1679585382
transform 1 0 138816 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_665
timestamp 1679585382
transform 1 0 139488 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_672
timestamp 1679585382
transform 1 0 140160 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_679
timestamp 1679585382
transform 1 0 140832 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_686
timestamp 1679585382
transform 1 0 141504 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_693
timestamp 1679585382
transform 1 0 142176 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_700
timestamp 1679585382
transform 1 0 142848 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_707
timestamp 1679585382
transform 1 0 143520 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_714
timestamp 1679585382
transform 1 0 144192 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_721
timestamp 1679585382
transform 1 0 144864 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_728
timestamp 1679585382
transform 1 0 145536 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_735
timestamp 1679585382
transform 1 0 146208 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_742
timestamp 1679585382
transform 1 0 146880 0 1 110376
box -48 -56 720 834
use sg13g2_decap_8  FILLER_46_749
timestamp 1679585382
transform 1 0 147552 0 1 110376
box -48 -56 720 834
use sg13g2_fill_1  FILLER_46_756
timestamp 1677583258
transform 1 0 148224 0 1 110376
box -48 -56 144 834
use sg13g2_decap_8  FILLER_47_0
timestamp 1679585382
transform 1 0 75648 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_7
timestamp 1679585382
transform 1 0 76320 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_14
timestamp 1679585382
transform 1 0 76992 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_21
timestamp 1679585382
transform 1 0 77664 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_28
timestamp 1679585382
transform 1 0 78336 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_35
timestamp 1679585382
transform 1 0 79008 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_42
timestamp 1679585382
transform 1 0 79680 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_49
timestamp 1679585382
transform 1 0 80352 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_56
timestamp 1679585382
transform 1 0 81024 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_63
timestamp 1679585382
transform 1 0 81696 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_70
timestamp 1679585382
transform 1 0 82368 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_77
timestamp 1679585382
transform 1 0 83040 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_84
timestamp 1679585382
transform 1 0 83712 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_91
timestamp 1679585382
transform 1 0 84384 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_98
timestamp 1679585382
transform 1 0 85056 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_105
timestamp 1679585382
transform 1 0 85728 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_112
timestamp 1679585382
transform 1 0 86400 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_119
timestamp 1679585382
transform 1 0 87072 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_126
timestamp 1679585382
transform 1 0 87744 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_133
timestamp 1679585382
transform 1 0 88416 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679585382
transform 1 0 89088 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_147
timestamp 1679585382
transform 1 0 89760 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_154
timestamp 1679585382
transform 1 0 90432 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_161
timestamp 1679585382
transform 1 0 91104 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_168
timestamp 1679585382
transform 1 0 91776 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_175
timestamp 1679585382
transform 1 0 92448 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_182
timestamp 1679585382
transform 1 0 93120 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_189
timestamp 1679585382
transform 1 0 93792 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_196
timestamp 1679585382
transform 1 0 94464 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_203
timestamp 1679585382
transform 1 0 95136 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_210
timestamp 1679585382
transform 1 0 95808 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_217
timestamp 1679585382
transform 1 0 96480 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_224
timestamp 1679585382
transform 1 0 97152 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_231
timestamp 1679585382
transform 1 0 97824 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_238
timestamp 1679585382
transform 1 0 98496 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_245
timestamp 1679585382
transform 1 0 99168 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_252
timestamp 1679585382
transform 1 0 99840 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_259
timestamp 1679585382
transform 1 0 100512 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_266
timestamp 1679585382
transform 1 0 101184 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_273
timestamp 1679585382
transform 1 0 101856 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_280
timestamp 1679585382
transform 1 0 102528 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_287
timestamp 1679585382
transform 1 0 103200 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_294
timestamp 1679585382
transform 1 0 103872 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_301
timestamp 1679585382
transform 1 0 104544 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_308
timestamp 1679585382
transform 1 0 105216 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_315
timestamp 1679585382
transform 1 0 105888 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_322
timestamp 1679585382
transform 1 0 106560 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_329
timestamp 1679585382
transform 1 0 107232 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_336
timestamp 1679585382
transform 1 0 107904 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_343
timestamp 1679585382
transform 1 0 108576 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_350
timestamp 1679585382
transform 1 0 109248 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_357
timestamp 1679585382
transform 1 0 109920 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_364
timestamp 1679585382
transform 1 0 110592 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_371
timestamp 1679585382
transform 1 0 111264 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_378
timestamp 1679585382
transform 1 0 111936 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_385
timestamp 1679585382
transform 1 0 112608 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_392
timestamp 1679585382
transform 1 0 113280 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_399
timestamp 1679585382
transform 1 0 113952 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_406
timestamp 1679585382
transform 1 0 114624 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_413
timestamp 1679585382
transform 1 0 115296 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_420
timestamp 1679585382
transform 1 0 115968 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_427
timestamp 1679585382
transform 1 0 116640 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_434
timestamp 1679585382
transform 1 0 117312 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_441
timestamp 1679585382
transform 1 0 117984 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_448
timestamp 1679585382
transform 1 0 118656 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_455
timestamp 1679585382
transform 1 0 119328 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_462
timestamp 1679585382
transform 1 0 120000 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_469
timestamp 1679585382
transform 1 0 120672 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_476
timestamp 1679585382
transform 1 0 121344 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_483
timestamp 1679585382
transform 1 0 122016 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_490
timestamp 1679585382
transform 1 0 122688 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_497
timestamp 1679585382
transform 1 0 123360 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_504
timestamp 1679585382
transform 1 0 124032 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_511
timestamp 1679585382
transform 1 0 124704 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_518
timestamp 1679585382
transform 1 0 125376 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_525
timestamp 1679585382
transform 1 0 126048 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_532
timestamp 1679585382
transform 1 0 126720 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_539
timestamp 1679585382
transform 1 0 127392 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_546
timestamp 1679585382
transform 1 0 128064 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_553
timestamp 1679585382
transform 1 0 128736 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_560
timestamp 1679585382
transform 1 0 129408 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_567
timestamp 1679585382
transform 1 0 130080 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_574
timestamp 1679585382
transform 1 0 130752 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_581
timestamp 1679585382
transform 1 0 131424 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_588
timestamp 1679585382
transform 1 0 132096 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_595
timestamp 1679585382
transform 1 0 132768 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_602
timestamp 1679585382
transform 1 0 133440 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_609
timestamp 1679585382
transform 1 0 134112 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_616
timestamp 1679585382
transform 1 0 134784 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_623
timestamp 1679585382
transform 1 0 135456 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_630
timestamp 1679585382
transform 1 0 136128 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_637
timestamp 1679585382
transform 1 0 136800 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_644
timestamp 1679585382
transform 1 0 137472 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_651
timestamp 1679585382
transform 1 0 138144 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_658
timestamp 1679585382
transform 1 0 138816 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_665
timestamp 1679585382
transform 1 0 139488 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_672
timestamp 1679585382
transform 1 0 140160 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_679
timestamp 1679585382
transform 1 0 140832 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_686
timestamp 1679585382
transform 1 0 141504 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_693
timestamp 1679585382
transform 1 0 142176 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_700
timestamp 1679585382
transform 1 0 142848 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_707
timestamp 1679585382
transform 1 0 143520 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_714
timestamp 1679585382
transform 1 0 144192 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_721
timestamp 1679585382
transform 1 0 144864 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_728
timestamp 1679585382
transform 1 0 145536 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_735
timestamp 1679585382
transform 1 0 146208 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_742
timestamp 1679585382
transform 1 0 146880 0 -1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_47_749
timestamp 1679585382
transform 1 0 147552 0 -1 111888
box -48 -56 720 834
use sg13g2_fill_1  FILLER_47_756
timestamp 1677583258
transform 1 0 148224 0 -1 111888
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_0
timestamp 1679585382
transform 1 0 75648 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_7
timestamp 1679585382
transform 1 0 76320 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_14
timestamp 1679585382
transform 1 0 76992 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_21
timestamp 1679585382
transform 1 0 77664 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_28
timestamp 1679585382
transform 1 0 78336 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_35
timestamp 1679585382
transform 1 0 79008 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_42
timestamp 1679585382
transform 1 0 79680 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_49
timestamp 1679585382
transform 1 0 80352 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_56
timestamp 1679585382
transform 1 0 81024 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_63
timestamp 1679585382
transform 1 0 81696 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_70
timestamp 1679585382
transform 1 0 82368 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_77
timestamp 1679585382
transform 1 0 83040 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_84
timestamp 1679585382
transform 1 0 83712 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_91
timestamp 1679585382
transform 1 0 84384 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_98
timestamp 1679585382
transform 1 0 85056 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_105
timestamp 1679585382
transform 1 0 85728 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_112
timestamp 1679585382
transform 1 0 86400 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_119
timestamp 1679585382
transform 1 0 87072 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_126
timestamp 1679585382
transform 1 0 87744 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_133
timestamp 1679585382
transform 1 0 88416 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_140
timestamp 1679585382
transform 1 0 89088 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_147
timestamp 1679585382
transform 1 0 89760 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_154
timestamp 1679585382
transform 1 0 90432 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_161
timestamp 1679585382
transform 1 0 91104 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_168
timestamp 1679585382
transform 1 0 91776 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_175
timestamp 1679585382
transform 1 0 92448 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_182
timestamp 1679585382
transform 1 0 93120 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_189
timestamp 1679585382
transform 1 0 93792 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_196
timestamp 1679585382
transform 1 0 94464 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_203
timestamp 1679585382
transform 1 0 95136 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_210
timestamp 1679585382
transform 1 0 95808 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_217
timestamp 1679585382
transform 1 0 96480 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_224
timestamp 1679585382
transform 1 0 97152 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_231
timestamp 1679585382
transform 1 0 97824 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_238
timestamp 1679585382
transform 1 0 98496 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_245
timestamp 1679585382
transform 1 0 99168 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_252
timestamp 1679585382
transform 1 0 99840 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_259
timestamp 1679585382
transform 1 0 100512 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_266
timestamp 1679585382
transform 1 0 101184 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_273
timestamp 1679585382
transform 1 0 101856 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_280
timestamp 1679585382
transform 1 0 102528 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_287
timestamp 1679585382
transform 1 0 103200 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_294
timestamp 1679585382
transform 1 0 103872 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_301
timestamp 1679585382
transform 1 0 104544 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_308
timestamp 1679585382
transform 1 0 105216 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_315
timestamp 1679585382
transform 1 0 105888 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_322
timestamp 1679585382
transform 1 0 106560 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_329
timestamp 1679585382
transform 1 0 107232 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_336
timestamp 1679585382
transform 1 0 107904 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_343
timestamp 1679585382
transform 1 0 108576 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_350
timestamp 1679585382
transform 1 0 109248 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_357
timestamp 1679585382
transform 1 0 109920 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_364
timestamp 1679585382
transform 1 0 110592 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_371
timestamp 1679585382
transform 1 0 111264 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_378
timestamp 1679585382
transform 1 0 111936 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_385
timestamp 1679585382
transform 1 0 112608 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_392
timestamp 1679585382
transform 1 0 113280 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_399
timestamp 1679585382
transform 1 0 113952 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_406
timestamp 1679585382
transform 1 0 114624 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_413
timestamp 1679585382
transform 1 0 115296 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_420
timestamp 1679585382
transform 1 0 115968 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_427
timestamp 1679585382
transform 1 0 116640 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_434
timestamp 1679585382
transform 1 0 117312 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_441
timestamp 1679585382
transform 1 0 117984 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_448
timestamp 1679585382
transform 1 0 118656 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_455
timestamp 1679585382
transform 1 0 119328 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_462
timestamp 1679585382
transform 1 0 120000 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_469
timestamp 1679585382
transform 1 0 120672 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_476
timestamp 1679585382
transform 1 0 121344 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_483
timestamp 1679585382
transform 1 0 122016 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_490
timestamp 1679585382
transform 1 0 122688 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_497
timestamp 1679585382
transform 1 0 123360 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_504
timestamp 1679585382
transform 1 0 124032 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_511
timestamp 1679585382
transform 1 0 124704 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_518
timestamp 1679585382
transform 1 0 125376 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_525
timestamp 1679585382
transform 1 0 126048 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_532
timestamp 1679585382
transform 1 0 126720 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_539
timestamp 1679585382
transform 1 0 127392 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_546
timestamp 1679585382
transform 1 0 128064 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_553
timestamp 1679585382
transform 1 0 128736 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_560
timestamp 1679585382
transform 1 0 129408 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_567
timestamp 1679585382
transform 1 0 130080 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_574
timestamp 1679585382
transform 1 0 130752 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_581
timestamp 1679585382
transform 1 0 131424 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_588
timestamp 1679585382
transform 1 0 132096 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_595
timestamp 1679585382
transform 1 0 132768 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_602
timestamp 1679585382
transform 1 0 133440 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_609
timestamp 1679585382
transform 1 0 134112 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_616
timestamp 1679585382
transform 1 0 134784 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_623
timestamp 1679585382
transform 1 0 135456 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_630
timestamp 1679585382
transform 1 0 136128 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_637
timestamp 1679585382
transform 1 0 136800 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_644
timestamp 1679585382
transform 1 0 137472 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_651
timestamp 1679585382
transform 1 0 138144 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_658
timestamp 1679585382
transform 1 0 138816 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_665
timestamp 1679585382
transform 1 0 139488 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_672
timestamp 1679585382
transform 1 0 140160 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_679
timestamp 1679585382
transform 1 0 140832 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_686
timestamp 1679585382
transform 1 0 141504 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_693
timestamp 1679585382
transform 1 0 142176 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_700
timestamp 1679585382
transform 1 0 142848 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_707
timestamp 1679585382
transform 1 0 143520 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_714
timestamp 1679585382
transform 1 0 144192 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_721
timestamp 1679585382
transform 1 0 144864 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_728
timestamp 1679585382
transform 1 0 145536 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_735
timestamp 1679585382
transform 1 0 146208 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_742
timestamp 1679585382
transform 1 0 146880 0 1 111888
box -48 -56 720 834
use sg13g2_decap_8  FILLER_48_749
timestamp 1679585382
transform 1 0 147552 0 1 111888
box -48 -56 720 834
use sg13g2_fill_1  FILLER_48_756
timestamp 1677583258
transform 1 0 148224 0 1 111888
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_0
timestamp 1679585382
transform 1 0 75648 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_7
timestamp 1679585382
transform 1 0 76320 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_14
timestamp 1679585382
transform 1 0 76992 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679585382
transform 1 0 77664 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_28
timestamp 1679585382
transform 1 0 78336 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_35
timestamp 1679585382
transform 1 0 79008 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_42
timestamp 1679585382
transform 1 0 79680 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_49
timestamp 1679585382
transform 1 0 80352 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_56
timestamp 1679585382
transform 1 0 81024 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_63
timestamp 1679585382
transform 1 0 81696 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_70
timestamp 1679585382
transform 1 0 82368 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_77
timestamp 1679585382
transform 1 0 83040 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_84
timestamp 1679585382
transform 1 0 83712 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_91
timestamp 1679585382
transform 1 0 84384 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_98
timestamp 1679585382
transform 1 0 85056 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_105
timestamp 1679585382
transform 1 0 85728 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_112
timestamp 1679585382
transform 1 0 86400 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_119
timestamp 1679585382
transform 1 0 87072 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_126
timestamp 1679585382
transform 1 0 87744 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_133
timestamp 1679585382
transform 1 0 88416 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_140
timestamp 1679585382
transform 1 0 89088 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_147
timestamp 1679585382
transform 1 0 89760 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_154
timestamp 1679585382
transform 1 0 90432 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_161
timestamp 1679585382
transform 1 0 91104 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_168
timestamp 1679585382
transform 1 0 91776 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_175
timestamp 1679585382
transform 1 0 92448 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_182
timestamp 1679585382
transform 1 0 93120 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_189
timestamp 1679585382
transform 1 0 93792 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_196
timestamp 1679585382
transform 1 0 94464 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_203
timestamp 1679585382
transform 1 0 95136 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_210
timestamp 1679585382
transform 1 0 95808 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_217
timestamp 1679585382
transform 1 0 96480 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_224
timestamp 1679585382
transform 1 0 97152 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_231
timestamp 1679585382
transform 1 0 97824 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_238
timestamp 1679585382
transform 1 0 98496 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_245
timestamp 1679585382
transform 1 0 99168 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_252
timestamp 1679585382
transform 1 0 99840 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_259
timestamp 1679585382
transform 1 0 100512 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_266
timestamp 1679585382
transform 1 0 101184 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_273
timestamp 1679585382
transform 1 0 101856 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_280
timestamp 1679585382
transform 1 0 102528 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_287
timestamp 1679585382
transform 1 0 103200 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_294
timestamp 1679585382
transform 1 0 103872 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_301
timestamp 1679585382
transform 1 0 104544 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_308
timestamp 1679585382
transform 1 0 105216 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_315
timestamp 1679585382
transform 1 0 105888 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_322
timestamp 1679585382
transform 1 0 106560 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_329
timestamp 1679585382
transform 1 0 107232 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_336
timestamp 1679585382
transform 1 0 107904 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_343
timestamp 1679585382
transform 1 0 108576 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_350
timestamp 1679585382
transform 1 0 109248 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_357
timestamp 1679585382
transform 1 0 109920 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_364
timestamp 1679585382
transform 1 0 110592 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_371
timestamp 1679585382
transform 1 0 111264 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_378
timestamp 1679585382
transform 1 0 111936 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_385
timestamp 1679585382
transform 1 0 112608 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_392
timestamp 1679585382
transform 1 0 113280 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_399
timestamp 1679585382
transform 1 0 113952 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_406
timestamp 1679585382
transform 1 0 114624 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_413
timestamp 1679585382
transform 1 0 115296 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_420
timestamp 1679585382
transform 1 0 115968 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_427
timestamp 1679585382
transform 1 0 116640 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_434
timestamp 1679585382
transform 1 0 117312 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_441
timestamp 1679585382
transform 1 0 117984 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_448
timestamp 1679585382
transform 1 0 118656 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_455
timestamp 1679585382
transform 1 0 119328 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_462
timestamp 1679585382
transform 1 0 120000 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_469
timestamp 1679585382
transform 1 0 120672 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_476
timestamp 1679585382
transform 1 0 121344 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_483
timestamp 1679585382
transform 1 0 122016 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_490
timestamp 1679585382
transform 1 0 122688 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_497
timestamp 1679585382
transform 1 0 123360 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_504
timestamp 1679585382
transform 1 0 124032 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_511
timestamp 1679585382
transform 1 0 124704 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_518
timestamp 1679585382
transform 1 0 125376 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_525
timestamp 1679585382
transform 1 0 126048 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_532
timestamp 1679585382
transform 1 0 126720 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_539
timestamp 1679585382
transform 1 0 127392 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_546
timestamp 1679585382
transform 1 0 128064 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_553
timestamp 1679585382
transform 1 0 128736 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_560
timestamp 1679585382
transform 1 0 129408 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_567
timestamp 1679585382
transform 1 0 130080 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_574
timestamp 1679585382
transform 1 0 130752 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_581
timestamp 1679585382
transform 1 0 131424 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_588
timestamp 1679585382
transform 1 0 132096 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_595
timestamp 1679585382
transform 1 0 132768 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_602
timestamp 1679585382
transform 1 0 133440 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_609
timestamp 1679585382
transform 1 0 134112 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_616
timestamp 1679585382
transform 1 0 134784 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_623
timestamp 1679585382
transform 1 0 135456 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_630
timestamp 1679585382
transform 1 0 136128 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_637
timestamp 1679585382
transform 1 0 136800 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_644
timestamp 1679585382
transform 1 0 137472 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_651
timestamp 1679585382
transform 1 0 138144 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_658
timestamp 1679585382
transform 1 0 138816 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_665
timestamp 1679585382
transform 1 0 139488 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_672
timestamp 1679585382
transform 1 0 140160 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_679
timestamp 1679585382
transform 1 0 140832 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_686
timestamp 1679585382
transform 1 0 141504 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_693
timestamp 1679585382
transform 1 0 142176 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_700
timestamp 1679585382
transform 1 0 142848 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_707
timestamp 1679585382
transform 1 0 143520 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_714
timestamp 1679585382
transform 1 0 144192 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_721
timestamp 1679585382
transform 1 0 144864 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_728
timestamp 1679585382
transform 1 0 145536 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_735
timestamp 1679585382
transform 1 0 146208 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_742
timestamp 1679585382
transform 1 0 146880 0 -1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_749
timestamp 1679585382
transform 1 0 147552 0 -1 113400
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_756
timestamp 1677583258
transform 1 0 148224 0 -1 113400
box -48 -56 144 834
use sg13g2_decap_8  FILLER_50_0
timestamp 1679585382
transform 1 0 75648 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_7
timestamp 1679585382
transform 1 0 76320 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_14
timestamp 1679585382
transform 1 0 76992 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_21
timestamp 1679585382
transform 1 0 77664 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_28
timestamp 1679585382
transform 1 0 78336 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_35
timestamp 1679585382
transform 1 0 79008 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_42
timestamp 1679585382
transform 1 0 79680 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_49
timestamp 1679585382
transform 1 0 80352 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_56
timestamp 1679585382
transform 1 0 81024 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_63
timestamp 1679585382
transform 1 0 81696 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_70
timestamp 1679585382
transform 1 0 82368 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_77
timestamp 1679585382
transform 1 0 83040 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_84
timestamp 1679585382
transform 1 0 83712 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_91
timestamp 1679585382
transform 1 0 84384 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_98
timestamp 1679585382
transform 1 0 85056 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_105
timestamp 1679585382
transform 1 0 85728 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_112
timestamp 1679585382
transform 1 0 86400 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_119
timestamp 1679585382
transform 1 0 87072 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_126
timestamp 1679585382
transform 1 0 87744 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_133
timestamp 1679585382
transform 1 0 88416 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_140
timestamp 1679585382
transform 1 0 89088 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_147
timestamp 1679585382
transform 1 0 89760 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_154
timestamp 1679585382
transform 1 0 90432 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_161
timestamp 1679585382
transform 1 0 91104 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_168
timestamp 1679585382
transform 1 0 91776 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_175
timestamp 1679585382
transform 1 0 92448 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_182
timestamp 1679585382
transform 1 0 93120 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_189
timestamp 1679585382
transform 1 0 93792 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_196
timestamp 1679585382
transform 1 0 94464 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_203
timestamp 1679585382
transform 1 0 95136 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_210
timestamp 1679585382
transform 1 0 95808 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_217
timestamp 1679585382
transform 1 0 96480 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_224
timestamp 1679585382
transform 1 0 97152 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_231
timestamp 1679585382
transform 1 0 97824 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_238
timestamp 1679585382
transform 1 0 98496 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_245
timestamp 1679585382
transform 1 0 99168 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_252
timestamp 1679585382
transform 1 0 99840 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_259
timestamp 1679585382
transform 1 0 100512 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_266
timestamp 1679585382
transform 1 0 101184 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_273
timestamp 1679585382
transform 1 0 101856 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_280
timestamp 1679585382
transform 1 0 102528 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_287
timestamp 1679585382
transform 1 0 103200 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_294
timestamp 1679585382
transform 1 0 103872 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_301
timestamp 1679585382
transform 1 0 104544 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_308
timestamp 1679585382
transform 1 0 105216 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_315
timestamp 1679585382
transform 1 0 105888 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_322
timestamp 1679585382
transform 1 0 106560 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_329
timestamp 1679585382
transform 1 0 107232 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_336
timestamp 1679585382
transform 1 0 107904 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_343
timestamp 1679585382
transform 1 0 108576 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_350
timestamp 1679585382
transform 1 0 109248 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_357
timestamp 1679585382
transform 1 0 109920 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_364
timestamp 1679585382
transform 1 0 110592 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_371
timestamp 1679585382
transform 1 0 111264 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_378
timestamp 1679585382
transform 1 0 111936 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_385
timestamp 1679585382
transform 1 0 112608 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_392
timestamp 1679585382
transform 1 0 113280 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_399
timestamp 1679585382
transform 1 0 113952 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_406
timestamp 1679585382
transform 1 0 114624 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_413
timestamp 1679585382
transform 1 0 115296 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_420
timestamp 1679585382
transform 1 0 115968 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_427
timestamp 1679585382
transform 1 0 116640 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_434
timestamp 1679585382
transform 1 0 117312 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_441
timestamp 1679585382
transform 1 0 117984 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_448
timestamp 1679585382
transform 1 0 118656 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_455
timestamp 1679585382
transform 1 0 119328 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_462
timestamp 1679585382
transform 1 0 120000 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_469
timestamp 1679585382
transform 1 0 120672 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_476
timestamp 1679585382
transform 1 0 121344 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_483
timestamp 1679585382
transform 1 0 122016 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_490
timestamp 1679585382
transform 1 0 122688 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_497
timestamp 1679585382
transform 1 0 123360 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_504
timestamp 1679585382
transform 1 0 124032 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_511
timestamp 1679585382
transform 1 0 124704 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_518
timestamp 1679585382
transform 1 0 125376 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_525
timestamp 1679585382
transform 1 0 126048 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_532
timestamp 1679585382
transform 1 0 126720 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_539
timestamp 1679585382
transform 1 0 127392 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_546
timestamp 1679585382
transform 1 0 128064 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_553
timestamp 1679585382
transform 1 0 128736 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_560
timestamp 1679585382
transform 1 0 129408 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_567
timestamp 1679585382
transform 1 0 130080 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_574
timestamp 1679585382
transform 1 0 130752 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_581
timestamp 1679585382
transform 1 0 131424 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_588
timestamp 1679585382
transform 1 0 132096 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_595
timestamp 1679585382
transform 1 0 132768 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_602
timestamp 1679585382
transform 1 0 133440 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_609
timestamp 1679585382
transform 1 0 134112 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_616
timestamp 1679585382
transform 1 0 134784 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_623
timestamp 1679585382
transform 1 0 135456 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_630
timestamp 1679585382
transform 1 0 136128 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_637
timestamp 1679585382
transform 1 0 136800 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_644
timestamp 1679585382
transform 1 0 137472 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_651
timestamp 1679585382
transform 1 0 138144 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_658
timestamp 1679585382
transform 1 0 138816 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_665
timestamp 1679585382
transform 1 0 139488 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_672
timestamp 1679585382
transform 1 0 140160 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_679
timestamp 1679585382
transform 1 0 140832 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_686
timestamp 1679585382
transform 1 0 141504 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_693
timestamp 1679585382
transform 1 0 142176 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_700
timestamp 1679585382
transform 1 0 142848 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_707
timestamp 1679585382
transform 1 0 143520 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_714
timestamp 1679585382
transform 1 0 144192 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_721
timestamp 1679585382
transform 1 0 144864 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_728
timestamp 1679585382
transform 1 0 145536 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_735
timestamp 1679585382
transform 1 0 146208 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_742
timestamp 1679585382
transform 1 0 146880 0 1 113400
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_749
timestamp 1679585382
transform 1 0 147552 0 1 113400
box -48 -56 720 834
use sg13g2_fill_1  FILLER_50_756
timestamp 1677583258
transform 1 0 148224 0 1 113400
box -48 -56 144 834
use sg13g2_decap_8  FILLER_51_0
timestamp 1679585382
transform 1 0 75648 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_7
timestamp 1679585382
transform 1 0 76320 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_14
timestamp 1679585382
transform 1 0 76992 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_21
timestamp 1679585382
transform 1 0 77664 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_28
timestamp 1679585382
transform 1 0 78336 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_35
timestamp 1679585382
transform 1 0 79008 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_42
timestamp 1679585382
transform 1 0 79680 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_49
timestamp 1679585382
transform 1 0 80352 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_56
timestamp 1679585382
transform 1 0 81024 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_63
timestamp 1679585382
transform 1 0 81696 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_70
timestamp 1679585382
transform 1 0 82368 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_77
timestamp 1679585382
transform 1 0 83040 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_84
timestamp 1679585382
transform 1 0 83712 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_91
timestamp 1679585382
transform 1 0 84384 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_98
timestamp 1679585382
transform 1 0 85056 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_105
timestamp 1679585382
transform 1 0 85728 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_112
timestamp 1679585382
transform 1 0 86400 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_119
timestamp 1679585382
transform 1 0 87072 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_126
timestamp 1679585382
transform 1 0 87744 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_133
timestamp 1679585382
transform 1 0 88416 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_140
timestamp 1679585382
transform 1 0 89088 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_147
timestamp 1679585382
transform 1 0 89760 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_154
timestamp 1679585382
transform 1 0 90432 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_161
timestamp 1679585382
transform 1 0 91104 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_168
timestamp 1679585382
transform 1 0 91776 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_175
timestamp 1679585382
transform 1 0 92448 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_182
timestamp 1679585382
transform 1 0 93120 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_189
timestamp 1679585382
transform 1 0 93792 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_196
timestamp 1679585382
transform 1 0 94464 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_203
timestamp 1679585382
transform 1 0 95136 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_210
timestamp 1679585382
transform 1 0 95808 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_217
timestamp 1679585382
transform 1 0 96480 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_224
timestamp 1679585382
transform 1 0 97152 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_231
timestamp 1679585382
transform 1 0 97824 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_238
timestamp 1679585382
transform 1 0 98496 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_245
timestamp 1679585382
transform 1 0 99168 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_252
timestamp 1679585382
transform 1 0 99840 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_259
timestamp 1679585382
transform 1 0 100512 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_266
timestamp 1679585382
transform 1 0 101184 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_273
timestamp 1679585382
transform 1 0 101856 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_280
timestamp 1679585382
transform 1 0 102528 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_287
timestamp 1679585382
transform 1 0 103200 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_294
timestamp 1679585382
transform 1 0 103872 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_301
timestamp 1679585382
transform 1 0 104544 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_308
timestamp 1679585382
transform 1 0 105216 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_315
timestamp 1679585382
transform 1 0 105888 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_322
timestamp 1679585382
transform 1 0 106560 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_329
timestamp 1679585382
transform 1 0 107232 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_336
timestamp 1679585382
transform 1 0 107904 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_343
timestamp 1679585382
transform 1 0 108576 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_350
timestamp 1679585382
transform 1 0 109248 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_357
timestamp 1679585382
transform 1 0 109920 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_364
timestamp 1679585382
transform 1 0 110592 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_371
timestamp 1679585382
transform 1 0 111264 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_378
timestamp 1679585382
transform 1 0 111936 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_385
timestamp 1679585382
transform 1 0 112608 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_392
timestamp 1679585382
transform 1 0 113280 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_399
timestamp 1679585382
transform 1 0 113952 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_406
timestamp 1679585382
transform 1 0 114624 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_413
timestamp 1679585382
transform 1 0 115296 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_420
timestamp 1679585382
transform 1 0 115968 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_427
timestamp 1679585382
transform 1 0 116640 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_434
timestamp 1679585382
transform 1 0 117312 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_441
timestamp 1679585382
transform 1 0 117984 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_448
timestamp 1679585382
transform 1 0 118656 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_455
timestamp 1679585382
transform 1 0 119328 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_462
timestamp 1679585382
transform 1 0 120000 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_469
timestamp 1679585382
transform 1 0 120672 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_476
timestamp 1679585382
transform 1 0 121344 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_483
timestamp 1679585382
transform 1 0 122016 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_490
timestamp 1679585382
transform 1 0 122688 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_497
timestamp 1679585382
transform 1 0 123360 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_504
timestamp 1679585382
transform 1 0 124032 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_511
timestamp 1679585382
transform 1 0 124704 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_518
timestamp 1679585382
transform 1 0 125376 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_525
timestamp 1679585382
transform 1 0 126048 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_532
timestamp 1679585382
transform 1 0 126720 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_539
timestamp 1679585382
transform 1 0 127392 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_546
timestamp 1679585382
transform 1 0 128064 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_553
timestamp 1679585382
transform 1 0 128736 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_560
timestamp 1679585382
transform 1 0 129408 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_567
timestamp 1679585382
transform 1 0 130080 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_574
timestamp 1679585382
transform 1 0 130752 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_581
timestamp 1679585382
transform 1 0 131424 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_588
timestamp 1679585382
transform 1 0 132096 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_595
timestamp 1679585382
transform 1 0 132768 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_602
timestamp 1679585382
transform 1 0 133440 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_609
timestamp 1679585382
transform 1 0 134112 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_616
timestamp 1679585382
transform 1 0 134784 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_623
timestamp 1679585382
transform 1 0 135456 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_630
timestamp 1679585382
transform 1 0 136128 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_637
timestamp 1679585382
transform 1 0 136800 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_644
timestamp 1679585382
transform 1 0 137472 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_651
timestamp 1679585382
transform 1 0 138144 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_658
timestamp 1679585382
transform 1 0 138816 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_665
timestamp 1679585382
transform 1 0 139488 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_672
timestamp 1679585382
transform 1 0 140160 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_679
timestamp 1679585382
transform 1 0 140832 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_686
timestamp 1679585382
transform 1 0 141504 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_693
timestamp 1679585382
transform 1 0 142176 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_700
timestamp 1679585382
transform 1 0 142848 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_707
timestamp 1679585382
transform 1 0 143520 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_714
timestamp 1679585382
transform 1 0 144192 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_721
timestamp 1679585382
transform 1 0 144864 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_728
timestamp 1679585382
transform 1 0 145536 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_735
timestamp 1679585382
transform 1 0 146208 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_742
timestamp 1679585382
transform 1 0 146880 0 -1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_51_749
timestamp 1679585382
transform 1 0 147552 0 -1 114912
box -48 -56 720 834
use sg13g2_fill_1  FILLER_51_756
timestamp 1677583258
transform 1 0 148224 0 -1 114912
box -48 -56 144 834
use sg13g2_decap_8  FILLER_52_0
timestamp 1679585382
transform 1 0 75648 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_7
timestamp 1679585382
transform 1 0 76320 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_14
timestamp 1679585382
transform 1 0 76992 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_21
timestamp 1679585382
transform 1 0 77664 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_28
timestamp 1679585382
transform 1 0 78336 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_35
timestamp 1679585382
transform 1 0 79008 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_42
timestamp 1679585382
transform 1 0 79680 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_49
timestamp 1679585382
transform 1 0 80352 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_56
timestamp 1679585382
transform 1 0 81024 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_63
timestamp 1679585382
transform 1 0 81696 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_70
timestamp 1679585382
transform 1 0 82368 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_77
timestamp 1679585382
transform 1 0 83040 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_84
timestamp 1679585382
transform 1 0 83712 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_91
timestamp 1679585382
transform 1 0 84384 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_98
timestamp 1679585382
transform 1 0 85056 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_105
timestamp 1679585382
transform 1 0 85728 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_112
timestamp 1679585382
transform 1 0 86400 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_119
timestamp 1679585382
transform 1 0 87072 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_126
timestamp 1679585382
transform 1 0 87744 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_133
timestamp 1679585382
transform 1 0 88416 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_140
timestamp 1679585382
transform 1 0 89088 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_147
timestamp 1679585382
transform 1 0 89760 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_154
timestamp 1679585382
transform 1 0 90432 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_161
timestamp 1679585382
transform 1 0 91104 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_168
timestamp 1679585382
transform 1 0 91776 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_175
timestamp 1679585382
transform 1 0 92448 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_182
timestamp 1679585382
transform 1 0 93120 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_189
timestamp 1679585382
transform 1 0 93792 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_196
timestamp 1679585382
transform 1 0 94464 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_203
timestamp 1679585382
transform 1 0 95136 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_210
timestamp 1679585382
transform 1 0 95808 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_217
timestamp 1679585382
transform 1 0 96480 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_224
timestamp 1679585382
transform 1 0 97152 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_231
timestamp 1679585382
transform 1 0 97824 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_238
timestamp 1679585382
transform 1 0 98496 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_245
timestamp 1679585382
transform 1 0 99168 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_252
timestamp 1679585382
transform 1 0 99840 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_259
timestamp 1679585382
transform 1 0 100512 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_266
timestamp 1679585382
transform 1 0 101184 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_273
timestamp 1679585382
transform 1 0 101856 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_280
timestamp 1679585382
transform 1 0 102528 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_287
timestamp 1679585382
transform 1 0 103200 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_294
timestamp 1679585382
transform 1 0 103872 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_301
timestamp 1679585382
transform 1 0 104544 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_308
timestamp 1679585382
transform 1 0 105216 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_315
timestamp 1679585382
transform 1 0 105888 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_322
timestamp 1679585382
transform 1 0 106560 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_329
timestamp 1679585382
transform 1 0 107232 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_336
timestamp 1679585382
transform 1 0 107904 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_343
timestamp 1679585382
transform 1 0 108576 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_350
timestamp 1679585382
transform 1 0 109248 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_357
timestamp 1679585382
transform 1 0 109920 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_364
timestamp 1679585382
transform 1 0 110592 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_371
timestamp 1679585382
transform 1 0 111264 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_378
timestamp 1679585382
transform 1 0 111936 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_385
timestamp 1679585382
transform 1 0 112608 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_392
timestamp 1679585382
transform 1 0 113280 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_399
timestamp 1679585382
transform 1 0 113952 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_406
timestamp 1679585382
transform 1 0 114624 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_413
timestamp 1679585382
transform 1 0 115296 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_420
timestamp 1679585382
transform 1 0 115968 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_427
timestamp 1679585382
transform 1 0 116640 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_434
timestamp 1679585382
transform 1 0 117312 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_441
timestamp 1679585382
transform 1 0 117984 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_448
timestamp 1679585382
transform 1 0 118656 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_455
timestamp 1679585382
transform 1 0 119328 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_462
timestamp 1679585382
transform 1 0 120000 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_469
timestamp 1679585382
transform 1 0 120672 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_476
timestamp 1679585382
transform 1 0 121344 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_483
timestamp 1679585382
transform 1 0 122016 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_490
timestamp 1679585382
transform 1 0 122688 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_497
timestamp 1679585382
transform 1 0 123360 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_504
timestamp 1679585382
transform 1 0 124032 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_511
timestamp 1679585382
transform 1 0 124704 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_518
timestamp 1679585382
transform 1 0 125376 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_525
timestamp 1679585382
transform 1 0 126048 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_532
timestamp 1679585382
transform 1 0 126720 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_539
timestamp 1679585382
transform 1 0 127392 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_546
timestamp 1679585382
transform 1 0 128064 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_553
timestamp 1679585382
transform 1 0 128736 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_560
timestamp 1679585382
transform 1 0 129408 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_567
timestamp 1679585382
transform 1 0 130080 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_574
timestamp 1679585382
transform 1 0 130752 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_581
timestamp 1679585382
transform 1 0 131424 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_588
timestamp 1679585382
transform 1 0 132096 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_595
timestamp 1679585382
transform 1 0 132768 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_602
timestamp 1679585382
transform 1 0 133440 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_609
timestamp 1679585382
transform 1 0 134112 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_616
timestamp 1679585382
transform 1 0 134784 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_623
timestamp 1679585382
transform 1 0 135456 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_630
timestamp 1679585382
transform 1 0 136128 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_637
timestamp 1679585382
transform 1 0 136800 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_644
timestamp 1679585382
transform 1 0 137472 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_651
timestamp 1679585382
transform 1 0 138144 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_658
timestamp 1679585382
transform 1 0 138816 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_665
timestamp 1679585382
transform 1 0 139488 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_672
timestamp 1679585382
transform 1 0 140160 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_679
timestamp 1679585382
transform 1 0 140832 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_686
timestamp 1679585382
transform 1 0 141504 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_693
timestamp 1679585382
transform 1 0 142176 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_700
timestamp 1679585382
transform 1 0 142848 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_707
timestamp 1679585382
transform 1 0 143520 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_714
timestamp 1679585382
transform 1 0 144192 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_721
timestamp 1679585382
transform 1 0 144864 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_728
timestamp 1679585382
transform 1 0 145536 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_735
timestamp 1679585382
transform 1 0 146208 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_742
timestamp 1679585382
transform 1 0 146880 0 1 114912
box -48 -56 720 834
use sg13g2_decap_8  FILLER_52_749
timestamp 1679585382
transform 1 0 147552 0 1 114912
box -48 -56 720 834
use sg13g2_fill_1  FILLER_52_756
timestamp 1677583258
transform 1 0 148224 0 1 114912
box -48 -56 144 834
use sg13g2_decap_8  FILLER_53_0
timestamp 1679585382
transform 1 0 75648 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_7
timestamp 1679585382
transform 1 0 76320 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_14
timestamp 1679585382
transform 1 0 76992 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_21
timestamp 1679585382
transform 1 0 77664 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_28
timestamp 1679585382
transform 1 0 78336 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_35
timestamp 1679585382
transform 1 0 79008 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_42
timestamp 1679585382
transform 1 0 79680 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_49
timestamp 1679585382
transform 1 0 80352 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_56
timestamp 1679585382
transform 1 0 81024 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_63
timestamp 1679585382
transform 1 0 81696 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_70
timestamp 1679585382
transform 1 0 82368 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_77
timestamp 1679585382
transform 1 0 83040 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_84
timestamp 1679585382
transform 1 0 83712 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_91
timestamp 1679585382
transform 1 0 84384 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_98
timestamp 1679585382
transform 1 0 85056 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_105
timestamp 1679585382
transform 1 0 85728 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_112
timestamp 1679585382
transform 1 0 86400 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_119
timestamp 1679585382
transform 1 0 87072 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_126
timestamp 1679585382
transform 1 0 87744 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_133
timestamp 1679585382
transform 1 0 88416 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_140
timestamp 1679585382
transform 1 0 89088 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_147
timestamp 1679585382
transform 1 0 89760 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_154
timestamp 1679585382
transform 1 0 90432 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_161
timestamp 1679585382
transform 1 0 91104 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_168
timestamp 1679585382
transform 1 0 91776 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_175
timestamp 1679585382
transform 1 0 92448 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_182
timestamp 1679585382
transform 1 0 93120 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_189
timestamp 1679585382
transform 1 0 93792 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_196
timestamp 1679585382
transform 1 0 94464 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_203
timestamp 1679585382
transform 1 0 95136 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_210
timestamp 1679585382
transform 1 0 95808 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_217
timestamp 1679585382
transform 1 0 96480 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_224
timestamp 1679585382
transform 1 0 97152 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_231
timestamp 1679585382
transform 1 0 97824 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_238
timestamp 1679585382
transform 1 0 98496 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_245
timestamp 1679585382
transform 1 0 99168 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_252
timestamp 1679585382
transform 1 0 99840 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_259
timestamp 1679585382
transform 1 0 100512 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_266
timestamp 1679585382
transform 1 0 101184 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_273
timestamp 1679585382
transform 1 0 101856 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_280
timestamp 1679585382
transform 1 0 102528 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_287
timestamp 1679585382
transform 1 0 103200 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_294
timestamp 1679585382
transform 1 0 103872 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_301
timestamp 1679585382
transform 1 0 104544 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_308
timestamp 1679585382
transform 1 0 105216 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_315
timestamp 1679585382
transform 1 0 105888 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_322
timestamp 1679585382
transform 1 0 106560 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_329
timestamp 1679585382
transform 1 0 107232 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_336
timestamp 1679585382
transform 1 0 107904 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_343
timestamp 1679585382
transform 1 0 108576 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_350
timestamp 1679585382
transform 1 0 109248 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_357
timestamp 1679585382
transform 1 0 109920 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_364
timestamp 1679585382
transform 1 0 110592 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_371
timestamp 1679585382
transform 1 0 111264 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_378
timestamp 1679585382
transform 1 0 111936 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_385
timestamp 1679585382
transform 1 0 112608 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_392
timestamp 1679585382
transform 1 0 113280 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_399
timestamp 1679585382
transform 1 0 113952 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_406
timestamp 1679585382
transform 1 0 114624 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_413
timestamp 1679585382
transform 1 0 115296 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_420
timestamp 1679585382
transform 1 0 115968 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_427
timestamp 1679585382
transform 1 0 116640 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_434
timestamp 1679585382
transform 1 0 117312 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_441
timestamp 1679585382
transform 1 0 117984 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_448
timestamp 1679585382
transform 1 0 118656 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_455
timestamp 1679585382
transform 1 0 119328 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_462
timestamp 1679585382
transform 1 0 120000 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_469
timestamp 1679585382
transform 1 0 120672 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_476
timestamp 1679585382
transform 1 0 121344 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_483
timestamp 1679585382
transform 1 0 122016 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_490
timestamp 1679585382
transform 1 0 122688 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_497
timestamp 1679585382
transform 1 0 123360 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_504
timestamp 1679585382
transform 1 0 124032 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_511
timestamp 1679585382
transform 1 0 124704 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_518
timestamp 1679585382
transform 1 0 125376 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_525
timestamp 1679585382
transform 1 0 126048 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_532
timestamp 1679585382
transform 1 0 126720 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_539
timestamp 1679585382
transform 1 0 127392 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_546
timestamp 1679585382
transform 1 0 128064 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_553
timestamp 1679585382
transform 1 0 128736 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_560
timestamp 1679585382
transform 1 0 129408 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_567
timestamp 1679585382
transform 1 0 130080 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_574
timestamp 1679585382
transform 1 0 130752 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_581
timestamp 1679585382
transform 1 0 131424 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_588
timestamp 1679585382
transform 1 0 132096 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_595
timestamp 1679585382
transform 1 0 132768 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_602
timestamp 1679585382
transform 1 0 133440 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_609
timestamp 1679585382
transform 1 0 134112 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_616
timestamp 1679585382
transform 1 0 134784 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_623
timestamp 1679585382
transform 1 0 135456 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_630
timestamp 1679585382
transform 1 0 136128 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_637
timestamp 1679585382
transform 1 0 136800 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_644
timestamp 1679585382
transform 1 0 137472 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_651
timestamp 1679585382
transform 1 0 138144 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_658
timestamp 1679585382
transform 1 0 138816 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_665
timestamp 1679585382
transform 1 0 139488 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_672
timestamp 1679585382
transform 1 0 140160 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_679
timestamp 1679585382
transform 1 0 140832 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_686
timestamp 1679585382
transform 1 0 141504 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_693
timestamp 1679585382
transform 1 0 142176 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_700
timestamp 1679585382
transform 1 0 142848 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_707
timestamp 1679585382
transform 1 0 143520 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_714
timestamp 1679585382
transform 1 0 144192 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_721
timestamp 1679585382
transform 1 0 144864 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_728
timestamp 1679585382
transform 1 0 145536 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_735
timestamp 1679585382
transform 1 0 146208 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_742
timestamp 1679585382
transform 1 0 146880 0 -1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_749
timestamp 1679585382
transform 1 0 147552 0 -1 116424
box -48 -56 720 834
use sg13g2_fill_1  FILLER_53_756
timestamp 1677583258
transform 1 0 148224 0 -1 116424
box -48 -56 144 834
use sg13g2_decap_8  FILLER_54_0
timestamp 1679585382
transform 1 0 75648 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_7
timestamp 1679585382
transform 1 0 76320 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_14
timestamp 1679585382
transform 1 0 76992 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_21
timestamp 1679585382
transform 1 0 77664 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_28
timestamp 1679585382
transform 1 0 78336 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_35
timestamp 1679585382
transform 1 0 79008 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_42
timestamp 1679585382
transform 1 0 79680 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_49
timestamp 1679585382
transform 1 0 80352 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_56
timestamp 1679585382
transform 1 0 81024 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_63
timestamp 1679585382
transform 1 0 81696 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_70
timestamp 1679585382
transform 1 0 82368 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_77
timestamp 1679585382
transform 1 0 83040 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_84
timestamp 1679585382
transform 1 0 83712 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_91
timestamp 1679585382
transform 1 0 84384 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_98
timestamp 1679585382
transform 1 0 85056 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_105
timestamp 1679585382
transform 1 0 85728 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_112
timestamp 1679585382
transform 1 0 86400 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_119
timestamp 1679585382
transform 1 0 87072 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_126
timestamp 1679585382
transform 1 0 87744 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_133
timestamp 1679585382
transform 1 0 88416 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_140
timestamp 1679585382
transform 1 0 89088 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_147
timestamp 1679585382
transform 1 0 89760 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_154
timestamp 1679585382
transform 1 0 90432 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_161
timestamp 1679585382
transform 1 0 91104 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_168
timestamp 1679585382
transform 1 0 91776 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_175
timestamp 1679585382
transform 1 0 92448 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_182
timestamp 1679585382
transform 1 0 93120 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_189
timestamp 1679585382
transform 1 0 93792 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_196
timestamp 1679585382
transform 1 0 94464 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_203
timestamp 1679585382
transform 1 0 95136 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_210
timestamp 1679585382
transform 1 0 95808 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_217
timestamp 1679585382
transform 1 0 96480 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_224
timestamp 1679585382
transform 1 0 97152 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_231
timestamp 1679585382
transform 1 0 97824 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_238
timestamp 1679585382
transform 1 0 98496 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_245
timestamp 1679585382
transform 1 0 99168 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_252
timestamp 1679585382
transform 1 0 99840 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_259
timestamp 1679585382
transform 1 0 100512 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_266
timestamp 1679585382
transform 1 0 101184 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_273
timestamp 1679585382
transform 1 0 101856 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_280
timestamp 1679585382
transform 1 0 102528 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_287
timestamp 1679585382
transform 1 0 103200 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_294
timestamp 1679585382
transform 1 0 103872 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_301
timestamp 1679585382
transform 1 0 104544 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_308
timestamp 1679585382
transform 1 0 105216 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_315
timestamp 1679585382
transform 1 0 105888 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_322
timestamp 1679585382
transform 1 0 106560 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_329
timestamp 1679585382
transform 1 0 107232 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_336
timestamp 1679585382
transform 1 0 107904 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_343
timestamp 1679585382
transform 1 0 108576 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_350
timestamp 1679585382
transform 1 0 109248 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_357
timestamp 1679585382
transform 1 0 109920 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_364
timestamp 1679585382
transform 1 0 110592 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_371
timestamp 1679585382
transform 1 0 111264 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_378
timestamp 1679585382
transform 1 0 111936 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_385
timestamp 1679585382
transform 1 0 112608 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_392
timestamp 1679585382
transform 1 0 113280 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_399
timestamp 1679585382
transform 1 0 113952 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_406
timestamp 1679585382
transform 1 0 114624 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_413
timestamp 1679585382
transform 1 0 115296 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_420
timestamp 1679585382
transform 1 0 115968 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_427
timestamp 1679585382
transform 1 0 116640 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_434
timestamp 1679585382
transform 1 0 117312 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_441
timestamp 1679585382
transform 1 0 117984 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_448
timestamp 1679585382
transform 1 0 118656 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_455
timestamp 1679585382
transform 1 0 119328 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_462
timestamp 1679585382
transform 1 0 120000 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_469
timestamp 1679585382
transform 1 0 120672 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_476
timestamp 1679585382
transform 1 0 121344 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_483
timestamp 1679585382
transform 1 0 122016 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_490
timestamp 1679585382
transform 1 0 122688 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_497
timestamp 1679585382
transform 1 0 123360 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_504
timestamp 1679585382
transform 1 0 124032 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_511
timestamp 1679585382
transform 1 0 124704 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_518
timestamp 1679585382
transform 1 0 125376 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_525
timestamp 1679585382
transform 1 0 126048 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_532
timestamp 1679585382
transform 1 0 126720 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_539
timestamp 1679585382
transform 1 0 127392 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_546
timestamp 1679585382
transform 1 0 128064 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_553
timestamp 1679585382
transform 1 0 128736 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_560
timestamp 1679585382
transform 1 0 129408 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_567
timestamp 1679585382
transform 1 0 130080 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_574
timestamp 1679585382
transform 1 0 130752 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_581
timestamp 1679585382
transform 1 0 131424 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_588
timestamp 1679585382
transform 1 0 132096 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_595
timestamp 1679585382
transform 1 0 132768 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_602
timestamp 1679585382
transform 1 0 133440 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_609
timestamp 1679585382
transform 1 0 134112 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_616
timestamp 1679585382
transform 1 0 134784 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_623
timestamp 1679585382
transform 1 0 135456 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_630
timestamp 1679585382
transform 1 0 136128 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_637
timestamp 1679585382
transform 1 0 136800 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_644
timestamp 1679585382
transform 1 0 137472 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_651
timestamp 1679585382
transform 1 0 138144 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_658
timestamp 1679585382
transform 1 0 138816 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_665
timestamp 1679585382
transform 1 0 139488 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_672
timestamp 1679585382
transform 1 0 140160 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_679
timestamp 1679585382
transform 1 0 140832 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_686
timestamp 1679585382
transform 1 0 141504 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_693
timestamp 1679585382
transform 1 0 142176 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_700
timestamp 1679585382
transform 1 0 142848 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_707
timestamp 1679585382
transform 1 0 143520 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_714
timestamp 1679585382
transform 1 0 144192 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_721
timestamp 1679585382
transform 1 0 144864 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_728
timestamp 1679585382
transform 1 0 145536 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_735
timestamp 1679585382
transform 1 0 146208 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_742
timestamp 1679585382
transform 1 0 146880 0 1 116424
box -48 -56 720 834
use sg13g2_decap_8  FILLER_54_749
timestamp 1679585382
transform 1 0 147552 0 1 116424
box -48 -56 720 834
use sg13g2_fill_1  FILLER_54_756
timestamp 1677583258
transform 1 0 148224 0 1 116424
box -48 -56 144 834
use sg13g2_decap_8  FILLER_55_0
timestamp 1679585382
transform 1 0 75648 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_7
timestamp 1679585382
transform 1 0 76320 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_14
timestamp 1679585382
transform 1 0 76992 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_21
timestamp 1679585382
transform 1 0 77664 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_28
timestamp 1679585382
transform 1 0 78336 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_35
timestamp 1679585382
transform 1 0 79008 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_42
timestamp 1679585382
transform 1 0 79680 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_49
timestamp 1679585382
transform 1 0 80352 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_56
timestamp 1679585382
transform 1 0 81024 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_63
timestamp 1679585382
transform 1 0 81696 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_70
timestamp 1679585382
transform 1 0 82368 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_77
timestamp 1679585382
transform 1 0 83040 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_84
timestamp 1679585382
transform 1 0 83712 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_91
timestamp 1679585382
transform 1 0 84384 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_98
timestamp 1679585382
transform 1 0 85056 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_105
timestamp 1679585382
transform 1 0 85728 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_112
timestamp 1679585382
transform 1 0 86400 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_119
timestamp 1679585382
transform 1 0 87072 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_126
timestamp 1679585382
transform 1 0 87744 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_133
timestamp 1679585382
transform 1 0 88416 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_140
timestamp 1679585382
transform 1 0 89088 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_147
timestamp 1679585382
transform 1 0 89760 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_154
timestamp 1679585382
transform 1 0 90432 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_161
timestamp 1679585382
transform 1 0 91104 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_168
timestamp 1679585382
transform 1 0 91776 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_175
timestamp 1679585382
transform 1 0 92448 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_182
timestamp 1679585382
transform 1 0 93120 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_189
timestamp 1679585382
transform 1 0 93792 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_196
timestamp 1679585382
transform 1 0 94464 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_203
timestamp 1679585382
transform 1 0 95136 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_210
timestamp 1679585382
transform 1 0 95808 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_217
timestamp 1679585382
transform 1 0 96480 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_224
timestamp 1679585382
transform 1 0 97152 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_231
timestamp 1679585382
transform 1 0 97824 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_238
timestamp 1679585382
transform 1 0 98496 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_245
timestamp 1679585382
transform 1 0 99168 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_252
timestamp 1679585382
transform 1 0 99840 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_259
timestamp 1679585382
transform 1 0 100512 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_266
timestamp 1679585382
transform 1 0 101184 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_273
timestamp 1679585382
transform 1 0 101856 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_280
timestamp 1679585382
transform 1 0 102528 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_287
timestamp 1679585382
transform 1 0 103200 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_294
timestamp 1679585382
transform 1 0 103872 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_301
timestamp 1679585382
transform 1 0 104544 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_308
timestamp 1679585382
transform 1 0 105216 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_315
timestamp 1679585382
transform 1 0 105888 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_322
timestamp 1679585382
transform 1 0 106560 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_329
timestamp 1679585382
transform 1 0 107232 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_336
timestamp 1679585382
transform 1 0 107904 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_343
timestamp 1679585382
transform 1 0 108576 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_350
timestamp 1679585382
transform 1 0 109248 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_357
timestamp 1679585382
transform 1 0 109920 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_364
timestamp 1679585382
transform 1 0 110592 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_371
timestamp 1679585382
transform 1 0 111264 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_378
timestamp 1679585382
transform 1 0 111936 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_385
timestamp 1679585382
transform 1 0 112608 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_392
timestamp 1679585382
transform 1 0 113280 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_399
timestamp 1679585382
transform 1 0 113952 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_406
timestamp 1679585382
transform 1 0 114624 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_413
timestamp 1679585382
transform 1 0 115296 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_420
timestamp 1679585382
transform 1 0 115968 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_427
timestamp 1679585382
transform 1 0 116640 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_434
timestamp 1679585382
transform 1 0 117312 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_441
timestamp 1679585382
transform 1 0 117984 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_448
timestamp 1679585382
transform 1 0 118656 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_455
timestamp 1679585382
transform 1 0 119328 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_462
timestamp 1679585382
transform 1 0 120000 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_469
timestamp 1679585382
transform 1 0 120672 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_476
timestamp 1679585382
transform 1 0 121344 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_483
timestamp 1679585382
transform 1 0 122016 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_490
timestamp 1679585382
transform 1 0 122688 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_497
timestamp 1679585382
transform 1 0 123360 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_504
timestamp 1679585382
transform 1 0 124032 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_511
timestamp 1679585382
transform 1 0 124704 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_518
timestamp 1679585382
transform 1 0 125376 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_525
timestamp 1679585382
transform 1 0 126048 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_532
timestamp 1679585382
transform 1 0 126720 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_539
timestamp 1679585382
transform 1 0 127392 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_546
timestamp 1679585382
transform 1 0 128064 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_553
timestamp 1679585382
transform 1 0 128736 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_560
timestamp 1679585382
transform 1 0 129408 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_567
timestamp 1679585382
transform 1 0 130080 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_574
timestamp 1679585382
transform 1 0 130752 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_581
timestamp 1679585382
transform 1 0 131424 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_588
timestamp 1679585382
transform 1 0 132096 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_595
timestamp 1679585382
transform 1 0 132768 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_602
timestamp 1679585382
transform 1 0 133440 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_609
timestamp 1679585382
transform 1 0 134112 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_616
timestamp 1679585382
transform 1 0 134784 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_623
timestamp 1679585382
transform 1 0 135456 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_630
timestamp 1679585382
transform 1 0 136128 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_637
timestamp 1679585382
transform 1 0 136800 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_644
timestamp 1679585382
transform 1 0 137472 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_651
timestamp 1679585382
transform 1 0 138144 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_658
timestamp 1679585382
transform 1 0 138816 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_665
timestamp 1679585382
transform 1 0 139488 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_672
timestamp 1679585382
transform 1 0 140160 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_679
timestamp 1679585382
transform 1 0 140832 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_686
timestamp 1679585382
transform 1 0 141504 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_693
timestamp 1679585382
transform 1 0 142176 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_700
timestamp 1679585382
transform 1 0 142848 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_707
timestamp 1679585382
transform 1 0 143520 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_714
timestamp 1679585382
transform 1 0 144192 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_721
timestamp 1679585382
transform 1 0 144864 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_728
timestamp 1679585382
transform 1 0 145536 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_735
timestamp 1679585382
transform 1 0 146208 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_742
timestamp 1679585382
transform 1 0 146880 0 -1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_749
timestamp 1679585382
transform 1 0 147552 0 -1 117936
box -48 -56 720 834
use sg13g2_fill_1  FILLER_55_756
timestamp 1677583258
transform 1 0 148224 0 -1 117936
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_0
timestamp 1679585382
transform 1 0 75648 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_7
timestamp 1679585382
transform 1 0 76320 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_14
timestamp 1679585382
transform 1 0 76992 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_21
timestamp 1679585382
transform 1 0 77664 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_28
timestamp 1679585382
transform 1 0 78336 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_35
timestamp 1679585382
transform 1 0 79008 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_42
timestamp 1679585382
transform 1 0 79680 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_49
timestamp 1679585382
transform 1 0 80352 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_56
timestamp 1679585382
transform 1 0 81024 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_63
timestamp 1679585382
transform 1 0 81696 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_70
timestamp 1679585382
transform 1 0 82368 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_77
timestamp 1679585382
transform 1 0 83040 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_84
timestamp 1679585382
transform 1 0 83712 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_91
timestamp 1679585382
transform 1 0 84384 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_98
timestamp 1679585382
transform 1 0 85056 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_105
timestamp 1679585382
transform 1 0 85728 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_112
timestamp 1679585382
transform 1 0 86400 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_119
timestamp 1679585382
transform 1 0 87072 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_126
timestamp 1679585382
transform 1 0 87744 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_133
timestamp 1679585382
transform 1 0 88416 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_140
timestamp 1679585382
transform 1 0 89088 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_147
timestamp 1679585382
transform 1 0 89760 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_154
timestamp 1679585382
transform 1 0 90432 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_161
timestamp 1679585382
transform 1 0 91104 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_168
timestamp 1679585382
transform 1 0 91776 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_175
timestamp 1679585382
transform 1 0 92448 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_182
timestamp 1679585382
transform 1 0 93120 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_189
timestamp 1679585382
transform 1 0 93792 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_196
timestamp 1679585382
transform 1 0 94464 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_203
timestamp 1679585382
transform 1 0 95136 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_210
timestamp 1679585382
transform 1 0 95808 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_217
timestamp 1679585382
transform 1 0 96480 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_224
timestamp 1679585382
transform 1 0 97152 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_231
timestamp 1679585382
transform 1 0 97824 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_238
timestamp 1679585382
transform 1 0 98496 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_245
timestamp 1679585382
transform 1 0 99168 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_252
timestamp 1679585382
transform 1 0 99840 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_259
timestamp 1679585382
transform 1 0 100512 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_266
timestamp 1679585382
transform 1 0 101184 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_273
timestamp 1679585382
transform 1 0 101856 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_280
timestamp 1679585382
transform 1 0 102528 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_287
timestamp 1679585382
transform 1 0 103200 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_294
timestamp 1679585382
transform 1 0 103872 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_301
timestamp 1679585382
transform 1 0 104544 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_308
timestamp 1679585382
transform 1 0 105216 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_315
timestamp 1679585382
transform 1 0 105888 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_322
timestamp 1679585382
transform 1 0 106560 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_329
timestamp 1679585382
transform 1 0 107232 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_336
timestamp 1679585382
transform 1 0 107904 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_343
timestamp 1679585382
transform 1 0 108576 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_350
timestamp 1679585382
transform 1 0 109248 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_357
timestamp 1679585382
transform 1 0 109920 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_364
timestamp 1679585382
transform 1 0 110592 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_371
timestamp 1679585382
transform 1 0 111264 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_378
timestamp 1679585382
transform 1 0 111936 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_385
timestamp 1679585382
transform 1 0 112608 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_392
timestamp 1679585382
transform 1 0 113280 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_399
timestamp 1679585382
transform 1 0 113952 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_406
timestamp 1679585382
transform 1 0 114624 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_413
timestamp 1679585382
transform 1 0 115296 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_420
timestamp 1679585382
transform 1 0 115968 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_427
timestamp 1679585382
transform 1 0 116640 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_434
timestamp 1679585382
transform 1 0 117312 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_441
timestamp 1679585382
transform 1 0 117984 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_448
timestamp 1679585382
transform 1 0 118656 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_455
timestamp 1679585382
transform 1 0 119328 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_462
timestamp 1679585382
transform 1 0 120000 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_469
timestamp 1679585382
transform 1 0 120672 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_476
timestamp 1679585382
transform 1 0 121344 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_483
timestamp 1679585382
transform 1 0 122016 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_490
timestamp 1679585382
transform 1 0 122688 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_497
timestamp 1679585382
transform 1 0 123360 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_504
timestamp 1679585382
transform 1 0 124032 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_511
timestamp 1679585382
transform 1 0 124704 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_518
timestamp 1679585382
transform 1 0 125376 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_525
timestamp 1679585382
transform 1 0 126048 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_532
timestamp 1679585382
transform 1 0 126720 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_539
timestamp 1679585382
transform 1 0 127392 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_546
timestamp 1679585382
transform 1 0 128064 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_553
timestamp 1679585382
transform 1 0 128736 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_560
timestamp 1679585382
transform 1 0 129408 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_567
timestamp 1679585382
transform 1 0 130080 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_574
timestamp 1679585382
transform 1 0 130752 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_581
timestamp 1679585382
transform 1 0 131424 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_588
timestamp 1679585382
transform 1 0 132096 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_595
timestamp 1679585382
transform 1 0 132768 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_602
timestamp 1679585382
transform 1 0 133440 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_609
timestamp 1679585382
transform 1 0 134112 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_616
timestamp 1679585382
transform 1 0 134784 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_623
timestamp 1679585382
transform 1 0 135456 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_630
timestamp 1679585382
transform 1 0 136128 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_637
timestamp 1679585382
transform 1 0 136800 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_644
timestamp 1679585382
transform 1 0 137472 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_651
timestamp 1679585382
transform 1 0 138144 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_658
timestamp 1679585382
transform 1 0 138816 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_665
timestamp 1679585382
transform 1 0 139488 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_672
timestamp 1679585382
transform 1 0 140160 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_679
timestamp 1679585382
transform 1 0 140832 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_686
timestamp 1679585382
transform 1 0 141504 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_693
timestamp 1679585382
transform 1 0 142176 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_700
timestamp 1679585382
transform 1 0 142848 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_707
timestamp 1679585382
transform 1 0 143520 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_714
timestamp 1679585382
transform 1 0 144192 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_721
timestamp 1679585382
transform 1 0 144864 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_728
timestamp 1679585382
transform 1 0 145536 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_735
timestamp 1679585382
transform 1 0 146208 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_742
timestamp 1679585382
transform 1 0 146880 0 1 117936
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_749
timestamp 1679585382
transform 1 0 147552 0 1 117936
box -48 -56 720 834
use sg13g2_fill_1  FILLER_56_756
timestamp 1677583258
transform 1 0 148224 0 1 117936
box -48 -56 144 834
use sg13g2_decap_8  FILLER_57_0
timestamp 1679585382
transform 1 0 75648 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_7
timestamp 1679585382
transform 1 0 76320 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_14
timestamp 1679585382
transform 1 0 76992 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_21
timestamp 1679585382
transform 1 0 77664 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_28
timestamp 1679585382
transform 1 0 78336 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_35
timestamp 1679585382
transform 1 0 79008 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_42
timestamp 1679585382
transform 1 0 79680 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_49
timestamp 1679585382
transform 1 0 80352 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_56
timestamp 1679585382
transform 1 0 81024 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_63
timestamp 1679585382
transform 1 0 81696 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_70
timestamp 1679585382
transform 1 0 82368 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_77
timestamp 1679585382
transform 1 0 83040 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_84
timestamp 1679585382
transform 1 0 83712 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_91
timestamp 1679585382
transform 1 0 84384 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_98
timestamp 1679585382
transform 1 0 85056 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_105
timestamp 1679585382
transform 1 0 85728 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_112
timestamp 1679585382
transform 1 0 86400 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_119
timestamp 1679585382
transform 1 0 87072 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_126
timestamp 1679585382
transform 1 0 87744 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_133
timestamp 1679585382
transform 1 0 88416 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_140
timestamp 1679585382
transform 1 0 89088 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_147
timestamp 1679585382
transform 1 0 89760 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_154
timestamp 1679585382
transform 1 0 90432 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_161
timestamp 1679585382
transform 1 0 91104 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_168
timestamp 1679585382
transform 1 0 91776 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_175
timestamp 1679585382
transform 1 0 92448 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_182
timestamp 1679585382
transform 1 0 93120 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_189
timestamp 1679585382
transform 1 0 93792 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_196
timestamp 1679585382
transform 1 0 94464 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_203
timestamp 1679585382
transform 1 0 95136 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_210
timestamp 1679585382
transform 1 0 95808 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_217
timestamp 1679585382
transform 1 0 96480 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_224
timestamp 1679585382
transform 1 0 97152 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_231
timestamp 1679585382
transform 1 0 97824 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_238
timestamp 1679585382
transform 1 0 98496 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_245
timestamp 1679585382
transform 1 0 99168 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_252
timestamp 1679585382
transform 1 0 99840 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_259
timestamp 1679585382
transform 1 0 100512 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_266
timestamp 1679585382
transform 1 0 101184 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_273
timestamp 1679585382
transform 1 0 101856 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_280
timestamp 1679585382
transform 1 0 102528 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_287
timestamp 1679585382
transform 1 0 103200 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_294
timestamp 1679585382
transform 1 0 103872 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_301
timestamp 1679585382
transform 1 0 104544 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_308
timestamp 1679585382
transform 1 0 105216 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_315
timestamp 1679585382
transform 1 0 105888 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_322
timestamp 1679585382
transform 1 0 106560 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_329
timestamp 1679585382
transform 1 0 107232 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_336
timestamp 1679585382
transform 1 0 107904 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_343
timestamp 1679585382
transform 1 0 108576 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_350
timestamp 1679585382
transform 1 0 109248 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_357
timestamp 1679585382
transform 1 0 109920 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_364
timestamp 1679585382
transform 1 0 110592 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_371
timestamp 1679585382
transform 1 0 111264 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_378
timestamp 1679585382
transform 1 0 111936 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_385
timestamp 1679585382
transform 1 0 112608 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_392
timestamp 1679585382
transform 1 0 113280 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_399
timestamp 1679585382
transform 1 0 113952 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_406
timestamp 1679585382
transform 1 0 114624 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_413
timestamp 1679585382
transform 1 0 115296 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_420
timestamp 1679585382
transform 1 0 115968 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_427
timestamp 1679585382
transform 1 0 116640 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_434
timestamp 1679585382
transform 1 0 117312 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_441
timestamp 1679585382
transform 1 0 117984 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_448
timestamp 1679585382
transform 1 0 118656 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_455
timestamp 1679585382
transform 1 0 119328 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_462
timestamp 1679585382
transform 1 0 120000 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_469
timestamp 1679585382
transform 1 0 120672 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_476
timestamp 1679585382
transform 1 0 121344 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_483
timestamp 1679585382
transform 1 0 122016 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_490
timestamp 1679585382
transform 1 0 122688 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_497
timestamp 1679585382
transform 1 0 123360 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_504
timestamp 1679585382
transform 1 0 124032 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_511
timestamp 1679585382
transform 1 0 124704 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_518
timestamp 1679585382
transform 1 0 125376 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_525
timestamp 1679585382
transform 1 0 126048 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_532
timestamp 1679585382
transform 1 0 126720 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_539
timestamp 1679585382
transform 1 0 127392 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_546
timestamp 1679585382
transform 1 0 128064 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_553
timestamp 1679585382
transform 1 0 128736 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_560
timestamp 1679585382
transform 1 0 129408 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_567
timestamp 1679585382
transform 1 0 130080 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_574
timestamp 1679585382
transform 1 0 130752 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_581
timestamp 1679585382
transform 1 0 131424 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_588
timestamp 1679585382
transform 1 0 132096 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_595
timestamp 1679585382
transform 1 0 132768 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_602
timestamp 1679585382
transform 1 0 133440 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_609
timestamp 1679585382
transform 1 0 134112 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_616
timestamp 1679585382
transform 1 0 134784 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_623
timestamp 1679585382
transform 1 0 135456 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_630
timestamp 1679585382
transform 1 0 136128 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_637
timestamp 1679585382
transform 1 0 136800 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_644
timestamp 1679585382
transform 1 0 137472 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_651
timestamp 1679585382
transform 1 0 138144 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_658
timestamp 1679585382
transform 1 0 138816 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_665
timestamp 1679585382
transform 1 0 139488 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_672
timestamp 1679585382
transform 1 0 140160 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_679
timestamp 1679585382
transform 1 0 140832 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_686
timestamp 1679585382
transform 1 0 141504 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_693
timestamp 1679585382
transform 1 0 142176 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_700
timestamp 1679585382
transform 1 0 142848 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_707
timestamp 1679585382
transform 1 0 143520 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_714
timestamp 1679585382
transform 1 0 144192 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_721
timestamp 1679585382
transform 1 0 144864 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_728
timestamp 1679585382
transform 1 0 145536 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_735
timestamp 1679585382
transform 1 0 146208 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_742
timestamp 1679585382
transform 1 0 146880 0 -1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_57_749
timestamp 1679585382
transform 1 0 147552 0 -1 119448
box -48 -56 720 834
use sg13g2_fill_1  FILLER_57_756
timestamp 1677583258
transform 1 0 148224 0 -1 119448
box -48 -56 144 834
use sg13g2_decap_8  FILLER_58_0
timestamp 1679585382
transform 1 0 75648 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_7
timestamp 1679585382
transform 1 0 76320 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_14
timestamp 1679585382
transform 1 0 76992 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_21
timestamp 1679585382
transform 1 0 77664 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_28
timestamp 1679585382
transform 1 0 78336 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_35
timestamp 1679585382
transform 1 0 79008 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_42
timestamp 1679585382
transform 1 0 79680 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_49
timestamp 1679585382
transform 1 0 80352 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_56
timestamp 1679585382
transform 1 0 81024 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_63
timestamp 1679585382
transform 1 0 81696 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_70
timestamp 1679585382
transform 1 0 82368 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_77
timestamp 1679585382
transform 1 0 83040 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_84
timestamp 1679585382
transform 1 0 83712 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_91
timestamp 1679585382
transform 1 0 84384 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_98
timestamp 1679585382
transform 1 0 85056 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_105
timestamp 1679585382
transform 1 0 85728 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_112
timestamp 1679585382
transform 1 0 86400 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_119
timestamp 1679585382
transform 1 0 87072 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_126
timestamp 1679585382
transform 1 0 87744 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_133
timestamp 1679585382
transform 1 0 88416 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_140
timestamp 1679585382
transform 1 0 89088 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_147
timestamp 1679585382
transform 1 0 89760 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_154
timestamp 1679585382
transform 1 0 90432 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_161
timestamp 1679585382
transform 1 0 91104 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_168
timestamp 1679585382
transform 1 0 91776 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_175
timestamp 1679585382
transform 1 0 92448 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_182
timestamp 1679585382
transform 1 0 93120 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_189
timestamp 1679585382
transform 1 0 93792 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_196
timestamp 1679585382
transform 1 0 94464 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_203
timestamp 1679585382
transform 1 0 95136 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_210
timestamp 1679585382
transform 1 0 95808 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_217
timestamp 1679585382
transform 1 0 96480 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_224
timestamp 1679585382
transform 1 0 97152 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_231
timestamp 1679585382
transform 1 0 97824 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_238
timestamp 1679585382
transform 1 0 98496 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_245
timestamp 1679585382
transform 1 0 99168 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_252
timestamp 1679585382
transform 1 0 99840 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_259
timestamp 1679585382
transform 1 0 100512 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_266
timestamp 1679585382
transform 1 0 101184 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_273
timestamp 1679585382
transform 1 0 101856 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_280
timestamp 1679585382
transform 1 0 102528 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_287
timestamp 1679585382
transform 1 0 103200 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_294
timestamp 1679585382
transform 1 0 103872 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_301
timestamp 1679585382
transform 1 0 104544 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_308
timestamp 1679585382
transform 1 0 105216 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_315
timestamp 1679585382
transform 1 0 105888 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_322
timestamp 1679585382
transform 1 0 106560 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_329
timestamp 1679585382
transform 1 0 107232 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_336
timestamp 1679585382
transform 1 0 107904 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_343
timestamp 1679585382
transform 1 0 108576 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_350
timestamp 1679585382
transform 1 0 109248 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_357
timestamp 1679585382
transform 1 0 109920 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_364
timestamp 1679585382
transform 1 0 110592 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_371
timestamp 1679585382
transform 1 0 111264 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_378
timestamp 1679585382
transform 1 0 111936 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_385
timestamp 1679585382
transform 1 0 112608 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_392
timestamp 1679585382
transform 1 0 113280 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_399
timestamp 1679585382
transform 1 0 113952 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_406
timestamp 1679585382
transform 1 0 114624 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_413
timestamp 1679585382
transform 1 0 115296 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_420
timestamp 1679585382
transform 1 0 115968 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_427
timestamp 1679585382
transform 1 0 116640 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_434
timestamp 1679585382
transform 1 0 117312 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_441
timestamp 1679585382
transform 1 0 117984 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_448
timestamp 1679585382
transform 1 0 118656 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_455
timestamp 1679585382
transform 1 0 119328 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_462
timestamp 1679585382
transform 1 0 120000 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_469
timestamp 1679585382
transform 1 0 120672 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_476
timestamp 1679585382
transform 1 0 121344 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_483
timestamp 1679585382
transform 1 0 122016 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_490
timestamp 1679585382
transform 1 0 122688 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_497
timestamp 1679585382
transform 1 0 123360 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_504
timestamp 1679585382
transform 1 0 124032 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_511
timestamp 1679585382
transform 1 0 124704 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_518
timestamp 1679585382
transform 1 0 125376 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_525
timestamp 1679585382
transform 1 0 126048 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_532
timestamp 1679585382
transform 1 0 126720 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_539
timestamp 1679585382
transform 1 0 127392 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_546
timestamp 1679585382
transform 1 0 128064 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_553
timestamp 1679585382
transform 1 0 128736 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_560
timestamp 1679585382
transform 1 0 129408 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_567
timestamp 1679585382
transform 1 0 130080 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_574
timestamp 1679585382
transform 1 0 130752 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_581
timestamp 1679585382
transform 1 0 131424 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_588
timestamp 1679585382
transform 1 0 132096 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_595
timestamp 1679585382
transform 1 0 132768 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_602
timestamp 1679585382
transform 1 0 133440 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_609
timestamp 1679585382
transform 1 0 134112 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_616
timestamp 1679585382
transform 1 0 134784 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_623
timestamp 1679585382
transform 1 0 135456 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_630
timestamp 1679585382
transform 1 0 136128 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_637
timestamp 1679585382
transform 1 0 136800 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_644
timestamp 1679585382
transform 1 0 137472 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_651
timestamp 1679585382
transform 1 0 138144 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_658
timestamp 1679585382
transform 1 0 138816 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_665
timestamp 1679585382
transform 1 0 139488 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_672
timestamp 1679585382
transform 1 0 140160 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_679
timestamp 1679585382
transform 1 0 140832 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_686
timestamp 1679585382
transform 1 0 141504 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_693
timestamp 1679585382
transform 1 0 142176 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_700
timestamp 1679585382
transform 1 0 142848 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_707
timestamp 1679585382
transform 1 0 143520 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_714
timestamp 1679585382
transform 1 0 144192 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_721
timestamp 1679585382
transform 1 0 144864 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_728
timestamp 1679585382
transform 1 0 145536 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_735
timestamp 1679585382
transform 1 0 146208 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_742
timestamp 1679585382
transform 1 0 146880 0 1 119448
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_749
timestamp 1679585382
transform 1 0 147552 0 1 119448
box -48 -56 720 834
use sg13g2_fill_1  FILLER_58_756
timestamp 1677583258
transform 1 0 148224 0 1 119448
box -48 -56 144 834
use sg13g2_decap_8  FILLER_59_0
timestamp 1679585382
transform 1 0 75648 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_7
timestamp 1679585382
transform 1 0 76320 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_14
timestamp 1679585382
transform 1 0 76992 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_21
timestamp 1679585382
transform 1 0 77664 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_28
timestamp 1679585382
transform 1 0 78336 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_35
timestamp 1679585382
transform 1 0 79008 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_42
timestamp 1679585382
transform 1 0 79680 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_49
timestamp 1679585382
transform 1 0 80352 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_56
timestamp 1679585382
transform 1 0 81024 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_63
timestamp 1679585382
transform 1 0 81696 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_70
timestamp 1679585382
transform 1 0 82368 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_77
timestamp 1679585382
transform 1 0 83040 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_84
timestamp 1679585382
transform 1 0 83712 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_91
timestamp 1679585382
transform 1 0 84384 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_98
timestamp 1679585382
transform 1 0 85056 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_105
timestamp 1679585382
transform 1 0 85728 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_112
timestamp 1679585382
transform 1 0 86400 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_119
timestamp 1679585382
transform 1 0 87072 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_126
timestamp 1679585382
transform 1 0 87744 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_133
timestamp 1679585382
transform 1 0 88416 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_140
timestamp 1679585382
transform 1 0 89088 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_147
timestamp 1679585382
transform 1 0 89760 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_154
timestamp 1679585382
transform 1 0 90432 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_161
timestamp 1679585382
transform 1 0 91104 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_168
timestamp 1679585382
transform 1 0 91776 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_175
timestamp 1679585382
transform 1 0 92448 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_182
timestamp 1679585382
transform 1 0 93120 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_189
timestamp 1679585382
transform 1 0 93792 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_196
timestamp 1679585382
transform 1 0 94464 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_203
timestamp 1679585382
transform 1 0 95136 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_210
timestamp 1679585382
transform 1 0 95808 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_217
timestamp 1679585382
transform 1 0 96480 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_224
timestamp 1679585382
transform 1 0 97152 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_231
timestamp 1679585382
transform 1 0 97824 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_238
timestamp 1679585382
transform 1 0 98496 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_245
timestamp 1679585382
transform 1 0 99168 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_252
timestamp 1679585382
transform 1 0 99840 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_259
timestamp 1679585382
transform 1 0 100512 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_266
timestamp 1679585382
transform 1 0 101184 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_273
timestamp 1679585382
transform 1 0 101856 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_280
timestamp 1679585382
transform 1 0 102528 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_287
timestamp 1679585382
transform 1 0 103200 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_294
timestamp 1679585382
transform 1 0 103872 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_301
timestamp 1679585382
transform 1 0 104544 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_308
timestamp 1679585382
transform 1 0 105216 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_315
timestamp 1679585382
transform 1 0 105888 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_322
timestamp 1679585382
transform 1 0 106560 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_329
timestamp 1679585382
transform 1 0 107232 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_336
timestamp 1679585382
transform 1 0 107904 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_343
timestamp 1679585382
transform 1 0 108576 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_350
timestamp 1679585382
transform 1 0 109248 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_357
timestamp 1679585382
transform 1 0 109920 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_364
timestamp 1679585382
transform 1 0 110592 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_371
timestamp 1679585382
transform 1 0 111264 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_378
timestamp 1679585382
transform 1 0 111936 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_385
timestamp 1679585382
transform 1 0 112608 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_392
timestamp 1679585382
transform 1 0 113280 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_399
timestamp 1679585382
transform 1 0 113952 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_406
timestamp 1679585382
transform 1 0 114624 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_413
timestamp 1679585382
transform 1 0 115296 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_420
timestamp 1679585382
transform 1 0 115968 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_427
timestamp 1679585382
transform 1 0 116640 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_434
timestamp 1679585382
transform 1 0 117312 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_441
timestamp 1679585382
transform 1 0 117984 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_448
timestamp 1679585382
transform 1 0 118656 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_455
timestamp 1679585382
transform 1 0 119328 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_462
timestamp 1679585382
transform 1 0 120000 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_469
timestamp 1679585382
transform 1 0 120672 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_476
timestamp 1679585382
transform 1 0 121344 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_483
timestamp 1679585382
transform 1 0 122016 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_490
timestamp 1679585382
transform 1 0 122688 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_497
timestamp 1679585382
transform 1 0 123360 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_504
timestamp 1679585382
transform 1 0 124032 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_511
timestamp 1679585382
transform 1 0 124704 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_518
timestamp 1679585382
transform 1 0 125376 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_525
timestamp 1679585382
transform 1 0 126048 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_532
timestamp 1679585382
transform 1 0 126720 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_539
timestamp 1679585382
transform 1 0 127392 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_546
timestamp 1679585382
transform 1 0 128064 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_553
timestamp 1679585382
transform 1 0 128736 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_560
timestamp 1679585382
transform 1 0 129408 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_567
timestamp 1679585382
transform 1 0 130080 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_574
timestamp 1679585382
transform 1 0 130752 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_581
timestamp 1679585382
transform 1 0 131424 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_588
timestamp 1679585382
transform 1 0 132096 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_595
timestamp 1679585382
transform 1 0 132768 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_602
timestamp 1679585382
transform 1 0 133440 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_609
timestamp 1679585382
transform 1 0 134112 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_616
timestamp 1679585382
transform 1 0 134784 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_623
timestamp 1679585382
transform 1 0 135456 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_630
timestamp 1679585382
transform 1 0 136128 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_637
timestamp 1679585382
transform 1 0 136800 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_644
timestamp 1679585382
transform 1 0 137472 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_651
timestamp 1679585382
transform 1 0 138144 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_658
timestamp 1679585382
transform 1 0 138816 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_665
timestamp 1679585382
transform 1 0 139488 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_672
timestamp 1679585382
transform 1 0 140160 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_679
timestamp 1679585382
transform 1 0 140832 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_686
timestamp 1679585382
transform 1 0 141504 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_693
timestamp 1679585382
transform 1 0 142176 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_700
timestamp 1679585382
transform 1 0 142848 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_707
timestamp 1679585382
transform 1 0 143520 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_714
timestamp 1679585382
transform 1 0 144192 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_721
timestamp 1679585382
transform 1 0 144864 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_728
timestamp 1679585382
transform 1 0 145536 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_735
timestamp 1679585382
transform 1 0 146208 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_742
timestamp 1679585382
transform 1 0 146880 0 -1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_749
timestamp 1679585382
transform 1 0 147552 0 -1 120960
box -48 -56 720 834
use sg13g2_fill_1  FILLER_59_756
timestamp 1677583258
transform 1 0 148224 0 -1 120960
box -48 -56 144 834
use sg13g2_decap_8  FILLER_60_0
timestamp 1679585382
transform 1 0 75648 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_7
timestamp 1679585382
transform 1 0 76320 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_14
timestamp 1679585382
transform 1 0 76992 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_21
timestamp 1679585382
transform 1 0 77664 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_28
timestamp 1679585382
transform 1 0 78336 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_35
timestamp 1679585382
transform 1 0 79008 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_42
timestamp 1679585382
transform 1 0 79680 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_49
timestamp 1679585382
transform 1 0 80352 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_56
timestamp 1679585382
transform 1 0 81024 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_63
timestamp 1679585382
transform 1 0 81696 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_70
timestamp 1679585382
transform 1 0 82368 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_77
timestamp 1679585382
transform 1 0 83040 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_84
timestamp 1679585382
transform 1 0 83712 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_91
timestamp 1679585382
transform 1 0 84384 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_98
timestamp 1679585382
transform 1 0 85056 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_105
timestamp 1679585382
transform 1 0 85728 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_112
timestamp 1679585382
transform 1 0 86400 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_119
timestamp 1679585382
transform 1 0 87072 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_126
timestamp 1679585382
transform 1 0 87744 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_133
timestamp 1679585382
transform 1 0 88416 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_140
timestamp 1679585382
transform 1 0 89088 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_147
timestamp 1679585382
transform 1 0 89760 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_154
timestamp 1679585382
transform 1 0 90432 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_161
timestamp 1679585382
transform 1 0 91104 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_168
timestamp 1679585382
transform 1 0 91776 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_175
timestamp 1679585382
transform 1 0 92448 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_182
timestamp 1679585382
transform 1 0 93120 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_189
timestamp 1679585382
transform 1 0 93792 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_196
timestamp 1679585382
transform 1 0 94464 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_203
timestamp 1679585382
transform 1 0 95136 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_210
timestamp 1679585382
transform 1 0 95808 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_217
timestamp 1679585382
transform 1 0 96480 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_224
timestamp 1679585382
transform 1 0 97152 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_231
timestamp 1679585382
transform 1 0 97824 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_238
timestamp 1679585382
transform 1 0 98496 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_245
timestamp 1679585382
transform 1 0 99168 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_252
timestamp 1679585382
transform 1 0 99840 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_259
timestamp 1679585382
transform 1 0 100512 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_266
timestamp 1679585382
transform 1 0 101184 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_273
timestamp 1679585382
transform 1 0 101856 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_280
timestamp 1679585382
transform 1 0 102528 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_287
timestamp 1679585382
transform 1 0 103200 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_294
timestamp 1679585382
transform 1 0 103872 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_301
timestamp 1679585382
transform 1 0 104544 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_308
timestamp 1679585382
transform 1 0 105216 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_315
timestamp 1679585382
transform 1 0 105888 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_322
timestamp 1679585382
transform 1 0 106560 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_329
timestamp 1679585382
transform 1 0 107232 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_336
timestamp 1679585382
transform 1 0 107904 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_343
timestamp 1679585382
transform 1 0 108576 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_350
timestamp 1679585382
transform 1 0 109248 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_357
timestamp 1679585382
transform 1 0 109920 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_364
timestamp 1679585382
transform 1 0 110592 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_371
timestamp 1679585382
transform 1 0 111264 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_378
timestamp 1679585382
transform 1 0 111936 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_385
timestamp 1679585382
transform 1 0 112608 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_392
timestamp 1679585382
transform 1 0 113280 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_399
timestamp 1679585382
transform 1 0 113952 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_406
timestamp 1679585382
transform 1 0 114624 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_413
timestamp 1679585382
transform 1 0 115296 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_420
timestamp 1679585382
transform 1 0 115968 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_427
timestamp 1679585382
transform 1 0 116640 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_434
timestamp 1679585382
transform 1 0 117312 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_441
timestamp 1679585382
transform 1 0 117984 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_448
timestamp 1679585382
transform 1 0 118656 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_455
timestamp 1679585382
transform 1 0 119328 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_462
timestamp 1679585382
transform 1 0 120000 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_469
timestamp 1679585382
transform 1 0 120672 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_476
timestamp 1679585382
transform 1 0 121344 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_483
timestamp 1679585382
transform 1 0 122016 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_490
timestamp 1679585382
transform 1 0 122688 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_497
timestamp 1679585382
transform 1 0 123360 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_504
timestamp 1679585382
transform 1 0 124032 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_511
timestamp 1679585382
transform 1 0 124704 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_518
timestamp 1679585382
transform 1 0 125376 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_525
timestamp 1679585382
transform 1 0 126048 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_532
timestamp 1679585382
transform 1 0 126720 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_539
timestamp 1679585382
transform 1 0 127392 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_546
timestamp 1679585382
transform 1 0 128064 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_553
timestamp 1679585382
transform 1 0 128736 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_560
timestamp 1679585382
transform 1 0 129408 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_567
timestamp 1679585382
transform 1 0 130080 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_574
timestamp 1679585382
transform 1 0 130752 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_581
timestamp 1679585382
transform 1 0 131424 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_588
timestamp 1679585382
transform 1 0 132096 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_595
timestamp 1679585382
transform 1 0 132768 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_602
timestamp 1679585382
transform 1 0 133440 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_609
timestamp 1679585382
transform 1 0 134112 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_616
timestamp 1679585382
transform 1 0 134784 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_623
timestamp 1679585382
transform 1 0 135456 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_630
timestamp 1679585382
transform 1 0 136128 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_637
timestamp 1679585382
transform 1 0 136800 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_644
timestamp 1679585382
transform 1 0 137472 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_651
timestamp 1679585382
transform 1 0 138144 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_658
timestamp 1679585382
transform 1 0 138816 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_665
timestamp 1679585382
transform 1 0 139488 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_672
timestamp 1679585382
transform 1 0 140160 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_679
timestamp 1679585382
transform 1 0 140832 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_686
timestamp 1679585382
transform 1 0 141504 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_693
timestamp 1679585382
transform 1 0 142176 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_700
timestamp 1679585382
transform 1 0 142848 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_707
timestamp 1679585382
transform 1 0 143520 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_714
timestamp 1679585382
transform 1 0 144192 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_721
timestamp 1679585382
transform 1 0 144864 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_728
timestamp 1679585382
transform 1 0 145536 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_735
timestamp 1679585382
transform 1 0 146208 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_742
timestamp 1679585382
transform 1 0 146880 0 1 120960
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_749
timestamp 1679585382
transform 1 0 147552 0 1 120960
box -48 -56 720 834
use sg13g2_fill_1  FILLER_60_756
timestamp 1677583258
transform 1 0 148224 0 1 120960
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_0
timestamp 1679585382
transform 1 0 75648 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_7
timestamp 1679585382
transform 1 0 76320 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_14
timestamp 1679585382
transform 1 0 76992 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_21
timestamp 1679585382
transform 1 0 77664 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_28
timestamp 1679585382
transform 1 0 78336 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_35
timestamp 1679585382
transform 1 0 79008 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_42
timestamp 1679585382
transform 1 0 79680 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_49
timestamp 1679585382
transform 1 0 80352 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_56
timestamp 1679585382
transform 1 0 81024 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_63
timestamp 1679585382
transform 1 0 81696 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_70
timestamp 1679585382
transform 1 0 82368 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_77
timestamp 1679585382
transform 1 0 83040 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_84
timestamp 1679585382
transform 1 0 83712 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_91
timestamp 1679585382
transform 1 0 84384 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_98
timestamp 1679585382
transform 1 0 85056 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_105
timestamp 1679585382
transform 1 0 85728 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_112
timestamp 1679585382
transform 1 0 86400 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_119
timestamp 1679585382
transform 1 0 87072 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_126
timestamp 1679585382
transform 1 0 87744 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_133
timestamp 1679585382
transform 1 0 88416 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_140
timestamp 1679585382
transform 1 0 89088 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_147
timestamp 1679585382
transform 1 0 89760 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_154
timestamp 1679585382
transform 1 0 90432 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_161
timestamp 1679585382
transform 1 0 91104 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_168
timestamp 1679585382
transform 1 0 91776 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_175
timestamp 1679585382
transform 1 0 92448 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_182
timestamp 1679585382
transform 1 0 93120 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_189
timestamp 1679585382
transform 1 0 93792 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_196
timestamp 1679585382
transform 1 0 94464 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_203
timestamp 1679585382
transform 1 0 95136 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_210
timestamp 1679585382
transform 1 0 95808 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_217
timestamp 1679585382
transform 1 0 96480 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_224
timestamp 1679585382
transform 1 0 97152 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_231
timestamp 1679585382
transform 1 0 97824 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_238
timestamp 1679585382
transform 1 0 98496 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_245
timestamp 1679585382
transform 1 0 99168 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_252
timestamp 1679585382
transform 1 0 99840 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_259
timestamp 1679585382
transform 1 0 100512 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_266
timestamp 1679585382
transform 1 0 101184 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_273
timestamp 1679585382
transform 1 0 101856 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_280
timestamp 1679585382
transform 1 0 102528 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_287
timestamp 1679585382
transform 1 0 103200 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_294
timestamp 1679585382
transform 1 0 103872 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_301
timestamp 1679585382
transform 1 0 104544 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_308
timestamp 1679585382
transform 1 0 105216 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_315
timestamp 1679585382
transform 1 0 105888 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_322
timestamp 1679585382
transform 1 0 106560 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_329
timestamp 1679585382
transform 1 0 107232 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_336
timestamp 1679585382
transform 1 0 107904 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_343
timestamp 1679585382
transform 1 0 108576 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_350
timestamp 1679585382
transform 1 0 109248 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_357
timestamp 1679585382
transform 1 0 109920 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_364
timestamp 1679585382
transform 1 0 110592 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_371
timestamp 1679585382
transform 1 0 111264 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_378
timestamp 1679585382
transform 1 0 111936 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_385
timestamp 1679585382
transform 1 0 112608 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_392
timestamp 1679585382
transform 1 0 113280 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_399
timestamp 1679585382
transform 1 0 113952 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_406
timestamp 1679585382
transform 1 0 114624 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_413
timestamp 1679585382
transform 1 0 115296 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_420
timestamp 1679585382
transform 1 0 115968 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_427
timestamp 1679585382
transform 1 0 116640 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_434
timestamp 1679585382
transform 1 0 117312 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_441
timestamp 1679585382
transform 1 0 117984 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_448
timestamp 1679585382
transform 1 0 118656 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_455
timestamp 1679585382
transform 1 0 119328 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_462
timestamp 1679585382
transform 1 0 120000 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_469
timestamp 1679585382
transform 1 0 120672 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_476
timestamp 1679585382
transform 1 0 121344 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_483
timestamp 1679585382
transform 1 0 122016 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_490
timestamp 1679585382
transform 1 0 122688 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_497
timestamp 1679585382
transform 1 0 123360 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_504
timestamp 1679585382
transform 1 0 124032 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_511
timestamp 1679585382
transform 1 0 124704 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_518
timestamp 1679585382
transform 1 0 125376 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_525
timestamp 1679585382
transform 1 0 126048 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_532
timestamp 1679585382
transform 1 0 126720 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_539
timestamp 1679585382
transform 1 0 127392 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_546
timestamp 1679585382
transform 1 0 128064 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_553
timestamp 1679585382
transform 1 0 128736 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_560
timestamp 1679585382
transform 1 0 129408 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_567
timestamp 1679585382
transform 1 0 130080 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_574
timestamp 1679585382
transform 1 0 130752 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_581
timestamp 1679585382
transform 1 0 131424 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_588
timestamp 1679585382
transform 1 0 132096 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_595
timestamp 1679585382
transform 1 0 132768 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_602
timestamp 1679585382
transform 1 0 133440 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_609
timestamp 1679585382
transform 1 0 134112 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_616
timestamp 1679585382
transform 1 0 134784 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_623
timestamp 1679585382
transform 1 0 135456 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_630
timestamp 1679585382
transform 1 0 136128 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_637
timestamp 1679585382
transform 1 0 136800 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_644
timestamp 1679585382
transform 1 0 137472 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_651
timestamp 1679585382
transform 1 0 138144 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_658
timestamp 1679585382
transform 1 0 138816 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_665
timestamp 1679585382
transform 1 0 139488 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_672
timestamp 1679585382
transform 1 0 140160 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_679
timestamp 1679585382
transform 1 0 140832 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_686
timestamp 1679585382
transform 1 0 141504 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_693
timestamp 1679585382
transform 1 0 142176 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_700
timestamp 1679585382
transform 1 0 142848 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_707
timestamp 1679585382
transform 1 0 143520 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_714
timestamp 1679585382
transform 1 0 144192 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_721
timestamp 1679585382
transform 1 0 144864 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_728
timestamp 1679585382
transform 1 0 145536 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_735
timestamp 1679585382
transform 1 0 146208 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_742
timestamp 1679585382
transform 1 0 146880 0 -1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_749
timestamp 1679585382
transform 1 0 147552 0 -1 122472
box -48 -56 720 834
use sg13g2_fill_1  FILLER_61_756
timestamp 1677583258
transform 1 0 148224 0 -1 122472
box -48 -56 144 834
use sg13g2_decap_8  FILLER_62_0
timestamp 1679585382
transform 1 0 75648 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_7
timestamp 1679585382
transform 1 0 76320 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_14
timestamp 1679585382
transform 1 0 76992 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_21
timestamp 1679585382
transform 1 0 77664 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_28
timestamp 1679585382
transform 1 0 78336 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_35
timestamp 1679585382
transform 1 0 79008 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_42
timestamp 1679585382
transform 1 0 79680 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_49
timestamp 1679585382
transform 1 0 80352 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_56
timestamp 1679585382
transform 1 0 81024 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_63
timestamp 1679585382
transform 1 0 81696 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_70
timestamp 1679585382
transform 1 0 82368 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_77
timestamp 1679585382
transform 1 0 83040 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_84
timestamp 1679585382
transform 1 0 83712 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_91
timestamp 1679585382
transform 1 0 84384 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_98
timestamp 1679585382
transform 1 0 85056 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_105
timestamp 1679585382
transform 1 0 85728 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_112
timestamp 1679585382
transform 1 0 86400 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_119
timestamp 1679585382
transform 1 0 87072 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_126
timestamp 1679585382
transform 1 0 87744 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_133
timestamp 1679585382
transform 1 0 88416 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_140
timestamp 1679585382
transform 1 0 89088 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_147
timestamp 1679585382
transform 1 0 89760 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_154
timestamp 1679585382
transform 1 0 90432 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_161
timestamp 1679585382
transform 1 0 91104 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_168
timestamp 1679585382
transform 1 0 91776 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_175
timestamp 1679585382
transform 1 0 92448 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_182
timestamp 1679585382
transform 1 0 93120 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_189
timestamp 1679585382
transform 1 0 93792 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_196
timestamp 1679585382
transform 1 0 94464 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_203
timestamp 1679585382
transform 1 0 95136 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_210
timestamp 1679585382
transform 1 0 95808 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_217
timestamp 1679585382
transform 1 0 96480 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_224
timestamp 1679585382
transform 1 0 97152 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_231
timestamp 1679585382
transform 1 0 97824 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_238
timestamp 1679585382
transform 1 0 98496 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_245
timestamp 1679585382
transform 1 0 99168 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_252
timestamp 1679585382
transform 1 0 99840 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_259
timestamp 1679585382
transform 1 0 100512 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_266
timestamp 1679585382
transform 1 0 101184 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_273
timestamp 1679585382
transform 1 0 101856 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_280
timestamp 1679585382
transform 1 0 102528 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_287
timestamp 1679585382
transform 1 0 103200 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_294
timestamp 1679585382
transform 1 0 103872 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_301
timestamp 1679585382
transform 1 0 104544 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_308
timestamp 1679585382
transform 1 0 105216 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_315
timestamp 1679585382
transform 1 0 105888 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_322
timestamp 1679585382
transform 1 0 106560 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_329
timestamp 1679585382
transform 1 0 107232 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_336
timestamp 1679585382
transform 1 0 107904 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_343
timestamp 1679585382
transform 1 0 108576 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_350
timestamp 1679585382
transform 1 0 109248 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_357
timestamp 1679585382
transform 1 0 109920 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_364
timestamp 1679585382
transform 1 0 110592 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_371
timestamp 1679585382
transform 1 0 111264 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_378
timestamp 1679585382
transform 1 0 111936 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_385
timestamp 1679585382
transform 1 0 112608 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_392
timestamp 1679585382
transform 1 0 113280 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_399
timestamp 1679585382
transform 1 0 113952 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_406
timestamp 1679585382
transform 1 0 114624 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_413
timestamp 1679585382
transform 1 0 115296 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_420
timestamp 1679585382
transform 1 0 115968 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_427
timestamp 1679585382
transform 1 0 116640 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_434
timestamp 1679585382
transform 1 0 117312 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_441
timestamp 1679585382
transform 1 0 117984 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_448
timestamp 1679585382
transform 1 0 118656 0 1 122472
box -48 -56 720 834
use sg13g2_fill_2  FILLER_62_455
timestamp 1677583704
transform 1 0 119328 0 1 122472
box -48 -56 240 834
use sg13g2_fill_1  FILLER_62_457
timestamp 1677583258
transform 1 0 119520 0 1 122472
box -48 -56 144 834
use sg13g2_decap_8  FILLER_62_462
timestamp 1679585382
transform 1 0 120000 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_469
timestamp 1679585382
transform 1 0 120672 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_476
timestamp 1679585382
transform 1 0 121344 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_483
timestamp 1679585382
transform 1 0 122016 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_490
timestamp 1679585382
transform 1 0 122688 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_497
timestamp 1679585382
transform 1 0 123360 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_504
timestamp 1679585382
transform 1 0 124032 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_511
timestamp 1679585382
transform 1 0 124704 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_518
timestamp 1679585382
transform 1 0 125376 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_525
timestamp 1679585382
transform 1 0 126048 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_532
timestamp 1679585382
transform 1 0 126720 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_539
timestamp 1679585382
transform 1 0 127392 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_546
timestamp 1679585382
transform 1 0 128064 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_553
timestamp 1679585382
transform 1 0 128736 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_560
timestamp 1679585382
transform 1 0 129408 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_567
timestamp 1679585382
transform 1 0 130080 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_574
timestamp 1679585382
transform 1 0 130752 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_581
timestamp 1679585382
transform 1 0 131424 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_588
timestamp 1679585382
transform 1 0 132096 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_595
timestamp 1679585382
transform 1 0 132768 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_602
timestamp 1679585382
transform 1 0 133440 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_609
timestamp 1679585382
transform 1 0 134112 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_616
timestamp 1679585382
transform 1 0 134784 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_623
timestamp 1679585382
transform 1 0 135456 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_630
timestamp 1679585382
transform 1 0 136128 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_637
timestamp 1679585382
transform 1 0 136800 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_644
timestamp 1679585382
transform 1 0 137472 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_651
timestamp 1679585382
transform 1 0 138144 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_658
timestamp 1679585382
transform 1 0 138816 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_665
timestamp 1679585382
transform 1 0 139488 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_672
timestamp 1679585382
transform 1 0 140160 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_679
timestamp 1679585382
transform 1 0 140832 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_686
timestamp 1679585382
transform 1 0 141504 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_693
timestamp 1679585382
transform 1 0 142176 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_700
timestamp 1679585382
transform 1 0 142848 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_707
timestamp 1679585382
transform 1 0 143520 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_714
timestamp 1679585382
transform 1 0 144192 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_721
timestamp 1679585382
transform 1 0 144864 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_728
timestamp 1679585382
transform 1 0 145536 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_735
timestamp 1679585382
transform 1 0 146208 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_742
timestamp 1679585382
transform 1 0 146880 0 1 122472
box -48 -56 720 834
use sg13g2_decap_8  FILLER_62_749
timestamp 1679585382
transform 1 0 147552 0 1 122472
box -48 -56 720 834
use sg13g2_fill_1  FILLER_62_756
timestamp 1677583258
transform 1 0 148224 0 1 122472
box -48 -56 144 834
use sg13g2_decap_8  FILLER_63_0
timestamp 1679585382
transform 1 0 75648 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_7
timestamp 1679585382
transform 1 0 76320 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_14
timestamp 1679585382
transform 1 0 76992 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_21
timestamp 1679585382
transform 1 0 77664 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_28
timestamp 1679585382
transform 1 0 78336 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_35
timestamp 1679585382
transform 1 0 79008 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_42
timestamp 1679585382
transform 1 0 79680 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_49
timestamp 1679585382
transform 1 0 80352 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_56
timestamp 1679585382
transform 1 0 81024 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_63
timestamp 1679585382
transform 1 0 81696 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_70
timestamp 1679585382
transform 1 0 82368 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_77
timestamp 1679585382
transform 1 0 83040 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_84
timestamp 1679585382
transform 1 0 83712 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_91
timestamp 1679585382
transform 1 0 84384 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_98
timestamp 1679585382
transform 1 0 85056 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_105
timestamp 1679585382
transform 1 0 85728 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_112
timestamp 1679585382
transform 1 0 86400 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_119
timestamp 1679585382
transform 1 0 87072 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_126
timestamp 1679585382
transform 1 0 87744 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_133
timestamp 1679585382
transform 1 0 88416 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_140
timestamp 1679585382
transform 1 0 89088 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_147
timestamp 1679585382
transform 1 0 89760 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_154
timestamp 1679585382
transform 1 0 90432 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_161
timestamp 1679585382
transform 1 0 91104 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_168
timestamp 1679585382
transform 1 0 91776 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_175
timestamp 1679585382
transform 1 0 92448 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_182
timestamp 1679585382
transform 1 0 93120 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_189
timestamp 1679585382
transform 1 0 93792 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_196
timestamp 1679585382
transform 1 0 94464 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_203
timestamp 1679585382
transform 1 0 95136 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_210
timestamp 1679585382
transform 1 0 95808 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_217
timestamp 1679585382
transform 1 0 96480 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_224
timestamp 1679585382
transform 1 0 97152 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_231
timestamp 1679585382
transform 1 0 97824 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_238
timestamp 1679585382
transform 1 0 98496 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_245
timestamp 1679585382
transform 1 0 99168 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_252
timestamp 1679585382
transform 1 0 99840 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_259
timestamp 1679585382
transform 1 0 100512 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_266
timestamp 1679585382
transform 1 0 101184 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_273
timestamp 1679585382
transform 1 0 101856 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_280
timestamp 1679585382
transform 1 0 102528 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_287
timestamp 1679585382
transform 1 0 103200 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_294
timestamp 1679585382
transform 1 0 103872 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_301
timestamp 1679585382
transform 1 0 104544 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_308
timestamp 1679585382
transform 1 0 105216 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_315
timestamp 1679585382
transform 1 0 105888 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_322
timestamp 1679585382
transform 1 0 106560 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_329
timestamp 1679585382
transform 1 0 107232 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_336
timestamp 1679585382
transform 1 0 107904 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_343
timestamp 1679585382
transform 1 0 108576 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_350
timestamp 1679585382
transform 1 0 109248 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_357
timestamp 1679585382
transform 1 0 109920 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_364
timestamp 1679585382
transform 1 0 110592 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_371
timestamp 1679585382
transform 1 0 111264 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_378
timestamp 1679585382
transform 1 0 111936 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_385
timestamp 1679585382
transform 1 0 112608 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_392
timestamp 1679585382
transform 1 0 113280 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_399
timestamp 1679585382
transform 1 0 113952 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_406
timestamp 1679585382
transform 1 0 114624 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_413
timestamp 1679585382
transform 1 0 115296 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_420
timestamp 1679585382
transform 1 0 115968 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_427
timestamp 1679585382
transform 1 0 116640 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_434
timestamp 1679585382
transform 1 0 117312 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_441
timestamp 1679585382
transform 1 0 117984 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_4  FILLER_63_448
timestamp 1679581501
transform 1 0 118656 0 -1 123984
box -48 -56 432 834
use sg13g2_fill_1  FILLER_63_452
timestamp 1677583258
transform 1 0 119040 0 -1 123984
box -48 -56 144 834
use sg13g2_decap_8  FILLER_63_480
timestamp 1679585382
transform 1 0 121728 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_487
timestamp 1679585382
transform 1 0 122400 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_494
timestamp 1679585382
transform 1 0 123072 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_501
timestamp 1679585382
transform 1 0 123744 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_508
timestamp 1679585382
transform 1 0 124416 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_515
timestamp 1679585382
transform 1 0 125088 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_522
timestamp 1679585382
transform 1 0 125760 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_529
timestamp 1679585382
transform 1 0 126432 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_536
timestamp 1679585382
transform 1 0 127104 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_543
timestamp 1679585382
transform 1 0 127776 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_550
timestamp 1679585382
transform 1 0 128448 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_557
timestamp 1679585382
transform 1 0 129120 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_564
timestamp 1679585382
transform 1 0 129792 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_571
timestamp 1679585382
transform 1 0 130464 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_578
timestamp 1679585382
transform 1 0 131136 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_585
timestamp 1679585382
transform 1 0 131808 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_592
timestamp 1679585382
transform 1 0 132480 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_599
timestamp 1679585382
transform 1 0 133152 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_606
timestamp 1679585382
transform 1 0 133824 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_613
timestamp 1679585382
transform 1 0 134496 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_620
timestamp 1679585382
transform 1 0 135168 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_627
timestamp 1679585382
transform 1 0 135840 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_634
timestamp 1679585382
transform 1 0 136512 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_641
timestamp 1679585382
transform 1 0 137184 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_648
timestamp 1679585382
transform 1 0 137856 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_655
timestamp 1679585382
transform 1 0 138528 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_662
timestamp 1679585382
transform 1 0 139200 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_669
timestamp 1679585382
transform 1 0 139872 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_676
timestamp 1679585382
transform 1 0 140544 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_683
timestamp 1679585382
transform 1 0 141216 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_690
timestamp 1679585382
transform 1 0 141888 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_697
timestamp 1679585382
transform 1 0 142560 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_704
timestamp 1679585382
transform 1 0 143232 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_711
timestamp 1679585382
transform 1 0 143904 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_718
timestamp 1679585382
transform 1 0 144576 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_725
timestamp 1679585382
transform 1 0 145248 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_732
timestamp 1679585382
transform 1 0 145920 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_739
timestamp 1679585382
transform 1 0 146592 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_63_746
timestamp 1679585382
transform 1 0 147264 0 -1 123984
box -48 -56 720 834
use sg13g2_decap_4  FILLER_63_753
timestamp 1679581501
transform 1 0 147936 0 -1 123984
box -48 -56 432 834
use sg13g2_decap_8  FILLER_64_0
timestamp 1679585382
transform 1 0 75648 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_7
timestamp 1679585382
transform 1 0 76320 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_14
timestamp 1679585382
transform 1 0 76992 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_21
timestamp 1679585382
transform 1 0 77664 0 1 123984
box -48 -56 720 834
use sg13g2_decap_4  FILLER_64_28
timestamp 1679581501
transform 1 0 78336 0 1 123984
box -48 -56 432 834
use sg13g2_fill_1  FILLER_64_32
timestamp 1677583258
transform 1 0 78720 0 1 123984
box -48 -56 144 834
use sg13g2_decap_8  FILLER_64_42
timestamp 1679585382
transform 1 0 79680 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_49
timestamp 1679585382
transform 1 0 80352 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_56
timestamp 1679585382
transform 1 0 81024 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_63
timestamp 1679585382
transform 1 0 81696 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_70
timestamp 1679585382
transform 1 0 82368 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_77
timestamp 1679585382
transform 1 0 83040 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_84
timestamp 1679585382
transform 1 0 83712 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_91
timestamp 1679585382
transform 1 0 84384 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_98
timestamp 1679585382
transform 1 0 85056 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_105
timestamp 1679585382
transform 1 0 85728 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_112
timestamp 1679585382
transform 1 0 86400 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_119
timestamp 1679585382
transform 1 0 87072 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_126
timestamp 1679585382
transform 1 0 87744 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_133
timestamp 1679585382
transform 1 0 88416 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_140
timestamp 1679585382
transform 1 0 89088 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_147
timestamp 1679585382
transform 1 0 89760 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_154
timestamp 1679585382
transform 1 0 90432 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_161
timestamp 1679585382
transform 1 0 91104 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_168
timestamp 1679585382
transform 1 0 91776 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_175
timestamp 1679585382
transform 1 0 92448 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_182
timestamp 1679585382
transform 1 0 93120 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_189
timestamp 1679585382
transform 1 0 93792 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_196
timestamp 1679585382
transform 1 0 94464 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_203
timestamp 1679585382
transform 1 0 95136 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_210
timestamp 1679585382
transform 1 0 95808 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_217
timestamp 1679585382
transform 1 0 96480 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_224
timestamp 1679585382
transform 1 0 97152 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_231
timestamp 1679585382
transform 1 0 97824 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_238
timestamp 1679585382
transform 1 0 98496 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_245
timestamp 1679585382
transform 1 0 99168 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_252
timestamp 1679585382
transform 1 0 99840 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_259
timestamp 1679585382
transform 1 0 100512 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_266
timestamp 1679585382
transform 1 0 101184 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_273
timestamp 1679585382
transform 1 0 101856 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_280
timestamp 1679585382
transform 1 0 102528 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_287
timestamp 1679585382
transform 1 0 103200 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_294
timestamp 1679585382
transform 1 0 103872 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_301
timestamp 1679585382
transform 1 0 104544 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_308
timestamp 1679585382
transform 1 0 105216 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_315
timestamp 1679585382
transform 1 0 105888 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_322
timestamp 1679585382
transform 1 0 106560 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_329
timestamp 1679585382
transform 1 0 107232 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_336
timestamp 1679585382
transform 1 0 107904 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_343
timestamp 1679585382
transform 1 0 108576 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_350
timestamp 1679585382
transform 1 0 109248 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_357
timestamp 1679585382
transform 1 0 109920 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_364
timestamp 1679585382
transform 1 0 110592 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_371
timestamp 1679585382
transform 1 0 111264 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_378
timestamp 1679585382
transform 1 0 111936 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_385
timestamp 1679585382
transform 1 0 112608 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_392
timestamp 1679585382
transform 1 0 113280 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_399
timestamp 1679585382
transform 1 0 113952 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_406
timestamp 1679585382
transform 1 0 114624 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_413
timestamp 1679585382
transform 1 0 115296 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_420
timestamp 1679585382
transform 1 0 115968 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_427
timestamp 1679585382
transform 1 0 116640 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_434
timestamp 1679585382
transform 1 0 117312 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_441
timestamp 1679585382
transform 1 0 117984 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_448
timestamp 1679585382
transform 1 0 118656 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_455
timestamp 1679585382
transform 1 0 119328 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_462
timestamp 1679585382
transform 1 0 120000 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_469
timestamp 1679585382
transform 1 0 120672 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_476
timestamp 1679585382
transform 1 0 121344 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_483
timestamp 1679585382
transform 1 0 122016 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_490
timestamp 1679585382
transform 1 0 122688 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_497
timestamp 1679585382
transform 1 0 123360 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_504
timestamp 1679585382
transform 1 0 124032 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_511
timestamp 1679585382
transform 1 0 124704 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_518
timestamp 1679585382
transform 1 0 125376 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_525
timestamp 1679585382
transform 1 0 126048 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_532
timestamp 1679585382
transform 1 0 126720 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_539
timestamp 1679585382
transform 1 0 127392 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_546
timestamp 1679585382
transform 1 0 128064 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_553
timestamp 1679585382
transform 1 0 128736 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_560
timestamp 1679585382
transform 1 0 129408 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_567
timestamp 1679585382
transform 1 0 130080 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_574
timestamp 1679585382
transform 1 0 130752 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_581
timestamp 1679585382
transform 1 0 131424 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_588
timestamp 1679585382
transform 1 0 132096 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_595
timestamp 1679585382
transform 1 0 132768 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_602
timestamp 1679585382
transform 1 0 133440 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_609
timestamp 1679585382
transform 1 0 134112 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_616
timestamp 1679585382
transform 1 0 134784 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_623
timestamp 1679585382
transform 1 0 135456 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_630
timestamp 1679585382
transform 1 0 136128 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_637
timestamp 1679585382
transform 1 0 136800 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_644
timestamp 1679585382
transform 1 0 137472 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_651
timestamp 1679585382
transform 1 0 138144 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_658
timestamp 1679585382
transform 1 0 138816 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_665
timestamp 1679585382
transform 1 0 139488 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_672
timestamp 1679585382
transform 1 0 140160 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_679
timestamp 1679585382
transform 1 0 140832 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_686
timestamp 1679585382
transform 1 0 141504 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_693
timestamp 1679585382
transform 1 0 142176 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_700
timestamp 1679585382
transform 1 0 142848 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_707
timestamp 1679585382
transform 1 0 143520 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_714
timestamp 1679585382
transform 1 0 144192 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_721
timestamp 1679585382
transform 1 0 144864 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_728
timestamp 1679585382
transform 1 0 145536 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_735
timestamp 1679585382
transform 1 0 146208 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_742
timestamp 1679585382
transform 1 0 146880 0 1 123984
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_749
timestamp 1679585382
transform 1 0 147552 0 1 123984
box -48 -56 720 834
use sg13g2_fill_1  FILLER_64_756
timestamp 1677583258
transform 1 0 148224 0 1 123984
box -48 -56 144 834
use sg13g2_decap_8  FILLER_65_0
timestamp 1679585382
transform 1 0 75648 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_7
timestamp 1679585382
transform 1 0 76320 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_14
timestamp 1679585382
transform 1 0 76992 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_21
timestamp 1679585382
transform 1 0 77664 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_28
timestamp 1679585382
transform 1 0 78336 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_35
timestamp 1679585382
transform 1 0 79008 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_42
timestamp 1679585382
transform 1 0 79680 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_49
timestamp 1679585382
transform 1 0 80352 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_56
timestamp 1679585382
transform 1 0 81024 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_63
timestamp 1679585382
transform 1 0 81696 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_70
timestamp 1679585382
transform 1 0 82368 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_77
timestamp 1679585382
transform 1 0 83040 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_84
timestamp 1679585382
transform 1 0 83712 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_91
timestamp 1679585382
transform 1 0 84384 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_98
timestamp 1679585382
transform 1 0 85056 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_105
timestamp 1679585382
transform 1 0 85728 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_112
timestamp 1679585382
transform 1 0 86400 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_119
timestamp 1679585382
transform 1 0 87072 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_126
timestamp 1679585382
transform 1 0 87744 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_133
timestamp 1679585382
transform 1 0 88416 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_140
timestamp 1679585382
transform 1 0 89088 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_147
timestamp 1679585382
transform 1 0 89760 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_154
timestamp 1679585382
transform 1 0 90432 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_161
timestamp 1679585382
transform 1 0 91104 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_168
timestamp 1679585382
transform 1 0 91776 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_175
timestamp 1679585382
transform 1 0 92448 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_182
timestamp 1679585382
transform 1 0 93120 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_189
timestamp 1679585382
transform 1 0 93792 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_196
timestamp 1679585382
transform 1 0 94464 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_203
timestamp 1679585382
transform 1 0 95136 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_210
timestamp 1679585382
transform 1 0 95808 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_217
timestamp 1679585382
transform 1 0 96480 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_224
timestamp 1679585382
transform 1 0 97152 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_231
timestamp 1679585382
transform 1 0 97824 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_238
timestamp 1679585382
transform 1 0 98496 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_245
timestamp 1679585382
transform 1 0 99168 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_252
timestamp 1679585382
transform 1 0 99840 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_259
timestamp 1679585382
transform 1 0 100512 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_266
timestamp 1679585382
transform 1 0 101184 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_273
timestamp 1679585382
transform 1 0 101856 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_280
timestamp 1679585382
transform 1 0 102528 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_287
timestamp 1679585382
transform 1 0 103200 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_294
timestamp 1679585382
transform 1 0 103872 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_301
timestamp 1679585382
transform 1 0 104544 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_308
timestamp 1679585382
transform 1 0 105216 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_315
timestamp 1679585382
transform 1 0 105888 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_322
timestamp 1679585382
transform 1 0 106560 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_329
timestamp 1679585382
transform 1 0 107232 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_336
timestamp 1679585382
transform 1 0 107904 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_343
timestamp 1679585382
transform 1 0 108576 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_350
timestamp 1679585382
transform 1 0 109248 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_357
timestamp 1679585382
transform 1 0 109920 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_364
timestamp 1679585382
transform 1 0 110592 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_371
timestamp 1679585382
transform 1 0 111264 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_378
timestamp 1679585382
transform 1 0 111936 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_385
timestamp 1679585382
transform 1 0 112608 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_392
timestamp 1679585382
transform 1 0 113280 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_399
timestamp 1679585382
transform 1 0 113952 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_406
timestamp 1679585382
transform 1 0 114624 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_413
timestamp 1679585382
transform 1 0 115296 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_420
timestamp 1679585382
transform 1 0 115968 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_427
timestamp 1679585382
transform 1 0 116640 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_434
timestamp 1679585382
transform 1 0 117312 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_441
timestamp 1679585382
transform 1 0 117984 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_448
timestamp 1679585382
transform 1 0 118656 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_455
timestamp 1679585382
transform 1 0 119328 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_462
timestamp 1679585382
transform 1 0 120000 0 -1 125496
box -48 -56 720 834
use sg13g2_fill_2  FILLER_65_469
timestamp 1677583704
transform 1 0 120672 0 -1 125496
box -48 -56 240 834
use sg13g2_fill_1  FILLER_65_471
timestamp 1677583258
transform 1 0 120864 0 -1 125496
box -48 -56 144 834
use sg13g2_fill_2  FILLER_65_475
timestamp 1677583704
transform 1 0 121248 0 -1 125496
box -48 -56 240 834
use sg13g2_decap_8  FILLER_65_486
timestamp 1679585382
transform 1 0 122304 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_493
timestamp 1679585382
transform 1 0 122976 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_500
timestamp 1679585382
transform 1 0 123648 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_507
timestamp 1679585382
transform 1 0 124320 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_514
timestamp 1679585382
transform 1 0 124992 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_521
timestamp 1679585382
transform 1 0 125664 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_528
timestamp 1679585382
transform 1 0 126336 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_535
timestamp 1679585382
transform 1 0 127008 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_542
timestamp 1679585382
transform 1 0 127680 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_549
timestamp 1679585382
transform 1 0 128352 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_556
timestamp 1679585382
transform 1 0 129024 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_563
timestamp 1679585382
transform 1 0 129696 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_570
timestamp 1679585382
transform 1 0 130368 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_577
timestamp 1679585382
transform 1 0 131040 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_584
timestamp 1679585382
transform 1 0 131712 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_591
timestamp 1679585382
transform 1 0 132384 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_598
timestamp 1679585382
transform 1 0 133056 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_605
timestamp 1679585382
transform 1 0 133728 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_612
timestamp 1679585382
transform 1 0 134400 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_619
timestamp 1679585382
transform 1 0 135072 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_626
timestamp 1679585382
transform 1 0 135744 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_633
timestamp 1679585382
transform 1 0 136416 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_640
timestamp 1679585382
transform 1 0 137088 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_647
timestamp 1679585382
transform 1 0 137760 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_654
timestamp 1679585382
transform 1 0 138432 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_661
timestamp 1679585382
transform 1 0 139104 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_668
timestamp 1679585382
transform 1 0 139776 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_675
timestamp 1679585382
transform 1 0 140448 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_682
timestamp 1679585382
transform 1 0 141120 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_689
timestamp 1679585382
transform 1 0 141792 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_696
timestamp 1679585382
transform 1 0 142464 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_703
timestamp 1679585382
transform 1 0 143136 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_710
timestamp 1679585382
transform 1 0 143808 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_717
timestamp 1679585382
transform 1 0 144480 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_724
timestamp 1679585382
transform 1 0 145152 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_731
timestamp 1679585382
transform 1 0 145824 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_738
timestamp 1679585382
transform 1 0 146496 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_65_745
timestamp 1679585382
transform 1 0 147168 0 -1 125496
box -48 -56 720 834
use sg13g2_decap_4  FILLER_65_752
timestamp 1679581501
transform 1 0 147840 0 -1 125496
box -48 -56 432 834
use sg13g2_fill_1  FILLER_65_756
timestamp 1677583258
transform 1 0 148224 0 -1 125496
box -48 -56 144 834
use sg13g2_decap_8  FILLER_66_0
timestamp 1679585382
transform 1 0 75648 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_7
timestamp 1679585382
transform 1 0 76320 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_14
timestamp 1679585382
transform 1 0 76992 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_21
timestamp 1679585382
transform 1 0 77664 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_28
timestamp 1679585382
transform 1 0 78336 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_35
timestamp 1679585382
transform 1 0 79008 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_42
timestamp 1679585382
transform 1 0 79680 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_49
timestamp 1679585382
transform 1 0 80352 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_56
timestamp 1679585382
transform 1 0 81024 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_63
timestamp 1679585382
transform 1 0 81696 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_70
timestamp 1679585382
transform 1 0 82368 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_77
timestamp 1679585382
transform 1 0 83040 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_84
timestamp 1679585382
transform 1 0 83712 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_91
timestamp 1679585382
transform 1 0 84384 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_98
timestamp 1679585382
transform 1 0 85056 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_105
timestamp 1679585382
transform 1 0 85728 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_112
timestamp 1679585382
transform 1 0 86400 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_119
timestamp 1679585382
transform 1 0 87072 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_126
timestamp 1679585382
transform 1 0 87744 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_133
timestamp 1679585382
transform 1 0 88416 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_140
timestamp 1679585382
transform 1 0 89088 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_147
timestamp 1679585382
transform 1 0 89760 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_154
timestamp 1679585382
transform 1 0 90432 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_161
timestamp 1679585382
transform 1 0 91104 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_168
timestamp 1679585382
transform 1 0 91776 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_175
timestamp 1679585382
transform 1 0 92448 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_182
timestamp 1679585382
transform 1 0 93120 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_189
timestamp 1679585382
transform 1 0 93792 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_196
timestamp 1679585382
transform 1 0 94464 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_203
timestamp 1679585382
transform 1 0 95136 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_210
timestamp 1679585382
transform 1 0 95808 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_217
timestamp 1679585382
transform 1 0 96480 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_224
timestamp 1679585382
transform 1 0 97152 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_231
timestamp 1679585382
transform 1 0 97824 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_238
timestamp 1679585382
transform 1 0 98496 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_245
timestamp 1679585382
transform 1 0 99168 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_252
timestamp 1679585382
transform 1 0 99840 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_259
timestamp 1679585382
transform 1 0 100512 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_266
timestamp 1679585382
transform 1 0 101184 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_273
timestamp 1679585382
transform 1 0 101856 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_280
timestamp 1679585382
transform 1 0 102528 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_287
timestamp 1679585382
transform 1 0 103200 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_294
timestamp 1679585382
transform 1 0 103872 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_301
timestamp 1679585382
transform 1 0 104544 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_308
timestamp 1679585382
transform 1 0 105216 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_315
timestamp 1679585382
transform 1 0 105888 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_322
timestamp 1679585382
transform 1 0 106560 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_329
timestamp 1679585382
transform 1 0 107232 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_336
timestamp 1679585382
transform 1 0 107904 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_343
timestamp 1679585382
transform 1 0 108576 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_350
timestamp 1679585382
transform 1 0 109248 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_357
timestamp 1679585382
transform 1 0 109920 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_364
timestamp 1679585382
transform 1 0 110592 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_371
timestamp 1679585382
transform 1 0 111264 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_378
timestamp 1679585382
transform 1 0 111936 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_385
timestamp 1679585382
transform 1 0 112608 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_392
timestamp 1679585382
transform 1 0 113280 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_399
timestamp 1679585382
transform 1 0 113952 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_406
timestamp 1679585382
transform 1 0 114624 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_413
timestamp 1679585382
transform 1 0 115296 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_420
timestamp 1679585382
transform 1 0 115968 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_427
timestamp 1679585382
transform 1 0 116640 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_434
timestamp 1679585382
transform 1 0 117312 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_441
timestamp 1679585382
transform 1 0 117984 0 1 125496
box -48 -56 720 834
use sg13g2_fill_2  FILLER_66_448
timestamp 1677583704
transform 1 0 118656 0 1 125496
box -48 -56 240 834
use sg13g2_decap_8  FILLER_66_457
timestamp 1679585382
transform 1 0 119520 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_464
timestamp 1679585382
transform 1 0 120192 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_471
timestamp 1679585382
transform 1 0 120864 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_478
timestamp 1679585382
transform 1 0 121536 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_485
timestamp 1679585382
transform 1 0 122208 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_492
timestamp 1679585382
transform 1 0 122880 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_499
timestamp 1679585382
transform 1 0 123552 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_506
timestamp 1679585382
transform 1 0 124224 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_513
timestamp 1679585382
transform 1 0 124896 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_520
timestamp 1679585382
transform 1 0 125568 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_527
timestamp 1679585382
transform 1 0 126240 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_534
timestamp 1679585382
transform 1 0 126912 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_541
timestamp 1679585382
transform 1 0 127584 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_548
timestamp 1679585382
transform 1 0 128256 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_555
timestamp 1679585382
transform 1 0 128928 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_562
timestamp 1679585382
transform 1 0 129600 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_569
timestamp 1679585382
transform 1 0 130272 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_576
timestamp 1679585382
transform 1 0 130944 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_583
timestamp 1679585382
transform 1 0 131616 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_590
timestamp 1679585382
transform 1 0 132288 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_597
timestamp 1679585382
transform 1 0 132960 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_604
timestamp 1679585382
transform 1 0 133632 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_611
timestamp 1679585382
transform 1 0 134304 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_618
timestamp 1679585382
transform 1 0 134976 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_625
timestamp 1679585382
transform 1 0 135648 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_632
timestamp 1679585382
transform 1 0 136320 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_639
timestamp 1679585382
transform 1 0 136992 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_646
timestamp 1679585382
transform 1 0 137664 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_653
timestamp 1679585382
transform 1 0 138336 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_660
timestamp 1679585382
transform 1 0 139008 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_667
timestamp 1679585382
transform 1 0 139680 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_674
timestamp 1679585382
transform 1 0 140352 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_681
timestamp 1679585382
transform 1 0 141024 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_688
timestamp 1679585382
transform 1 0 141696 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_695
timestamp 1679585382
transform 1 0 142368 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_702
timestamp 1679585382
transform 1 0 143040 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_709
timestamp 1679585382
transform 1 0 143712 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_716
timestamp 1679585382
transform 1 0 144384 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_723
timestamp 1679585382
transform 1 0 145056 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_730
timestamp 1679585382
transform 1 0 145728 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_737
timestamp 1679585382
transform 1 0 146400 0 1 125496
box -48 -56 720 834
use sg13g2_decap_8  FILLER_66_744
timestamp 1679585382
transform 1 0 147072 0 1 125496
box -48 -56 720 834
use sg13g2_decap_4  FILLER_66_751
timestamp 1679581501
transform 1 0 147744 0 1 125496
box -48 -56 432 834
use sg13g2_fill_2  FILLER_66_755
timestamp 1677583704
transform 1 0 148128 0 1 125496
box -48 -56 240 834
use sg13g2_decap_8  FILLER_67_0
timestamp 1679585382
transform 1 0 75648 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_7
timestamp 1679585382
transform 1 0 76320 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_14
timestamp 1679585382
transform 1 0 76992 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_21
timestamp 1679585382
transform 1 0 77664 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_28
timestamp 1679585382
transform 1 0 78336 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_35
timestamp 1679585382
transform 1 0 79008 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_42
timestamp 1679585382
transform 1 0 79680 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_49
timestamp 1679585382
transform 1 0 80352 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_56
timestamp 1679585382
transform 1 0 81024 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_63
timestamp 1679585382
transform 1 0 81696 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_70
timestamp 1679585382
transform 1 0 82368 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_77
timestamp 1679585382
transform 1 0 83040 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_84
timestamp 1679585382
transform 1 0 83712 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_91
timestamp 1679585382
transform 1 0 84384 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_98
timestamp 1679585382
transform 1 0 85056 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_105
timestamp 1679585382
transform 1 0 85728 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_112
timestamp 1679585382
transform 1 0 86400 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_119
timestamp 1679585382
transform 1 0 87072 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_126
timestamp 1679585382
transform 1 0 87744 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_133
timestamp 1679585382
transform 1 0 88416 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_140
timestamp 1679585382
transform 1 0 89088 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_147
timestamp 1679585382
transform 1 0 89760 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_154
timestamp 1679585382
transform 1 0 90432 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_161
timestamp 1679585382
transform 1 0 91104 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_168
timestamp 1679585382
transform 1 0 91776 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_175
timestamp 1679585382
transform 1 0 92448 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_182
timestamp 1679585382
transform 1 0 93120 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_189
timestamp 1679585382
transform 1 0 93792 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_4  FILLER_67_202
timestamp 1679581501
transform 1 0 95040 0 -1 127008
box -48 -56 432 834
use sg13g2_decap_8  FILLER_67_212
timestamp 1679585382
transform 1 0 96000 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_219
timestamp 1679585382
transform 1 0 96672 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_226
timestamp 1679585382
transform 1 0 97344 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_233
timestamp 1679585382
transform 1 0 98016 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_240
timestamp 1679585382
transform 1 0 98688 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_247
timestamp 1679585382
transform 1 0 99360 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_254
timestamp 1679585382
transform 1 0 100032 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_261
timestamp 1679585382
transform 1 0 100704 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_268
timestamp 1679585382
transform 1 0 101376 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_275
timestamp 1679585382
transform 1 0 102048 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_282
timestamp 1679585382
transform 1 0 102720 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_289
timestamp 1679585382
transform 1 0 103392 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_296
timestamp 1679585382
transform 1 0 104064 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_303
timestamp 1679585382
transform 1 0 104736 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_310
timestamp 1679585382
transform 1 0 105408 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_317
timestamp 1679585382
transform 1 0 106080 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_324
timestamp 1679585382
transform 1 0 106752 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_331
timestamp 1679585382
transform 1 0 107424 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_338
timestamp 1679585382
transform 1 0 108096 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_345
timestamp 1679585382
transform 1 0 108768 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_352
timestamp 1679585382
transform 1 0 109440 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_359
timestamp 1679585382
transform 1 0 110112 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_366
timestamp 1679585382
transform 1 0 110784 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_373
timestamp 1679585382
transform 1 0 111456 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_380
timestamp 1679585382
transform 1 0 112128 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_387
timestamp 1679585382
transform 1 0 112800 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_394
timestamp 1679585382
transform 1 0 113472 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_401
timestamp 1679585382
transform 1 0 114144 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_408
timestamp 1679585382
transform 1 0 114816 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_415
timestamp 1679585382
transform 1 0 115488 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_422
timestamp 1679585382
transform 1 0 116160 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_429
timestamp 1679585382
transform 1 0 116832 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_436
timestamp 1679585382
transform 1 0 117504 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_443
timestamp 1679585382
transform 1 0 118176 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_450
timestamp 1679585382
transform 1 0 118848 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_457
timestamp 1679585382
transform 1 0 119520 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_464
timestamp 1679585382
transform 1 0 120192 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_471
timestamp 1679585382
transform 1 0 120864 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_478
timestamp 1679585382
transform 1 0 121536 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_485
timestamp 1679585382
transform 1 0 122208 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_492
timestamp 1679585382
transform 1 0 122880 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_499
timestamp 1679585382
transform 1 0 123552 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_506
timestamp 1679585382
transform 1 0 124224 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_513
timestamp 1679585382
transform 1 0 124896 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_520
timestamp 1679585382
transform 1 0 125568 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_527
timestamp 1679585382
transform 1 0 126240 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_534
timestamp 1679585382
transform 1 0 126912 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_541
timestamp 1679585382
transform 1 0 127584 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_548
timestamp 1679585382
transform 1 0 128256 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_555
timestamp 1679585382
transform 1 0 128928 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_562
timestamp 1679585382
transform 1 0 129600 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_569
timestamp 1679585382
transform 1 0 130272 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_576
timestamp 1679585382
transform 1 0 130944 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_583
timestamp 1679585382
transform 1 0 131616 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_590
timestamp 1679585382
transform 1 0 132288 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_597
timestamp 1679585382
transform 1 0 132960 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_604
timestamp 1679585382
transform 1 0 133632 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_611
timestamp 1679585382
transform 1 0 134304 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_618
timestamp 1679585382
transform 1 0 134976 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_625
timestamp 1679585382
transform 1 0 135648 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_632
timestamp 1679585382
transform 1 0 136320 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_639
timestamp 1679585382
transform 1 0 136992 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_646
timestamp 1679585382
transform 1 0 137664 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_653
timestamp 1679585382
transform 1 0 138336 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_660
timestamp 1679585382
transform 1 0 139008 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_667
timestamp 1679585382
transform 1 0 139680 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_674
timestamp 1679585382
transform 1 0 140352 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_681
timestamp 1679585382
transform 1 0 141024 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_688
timestamp 1679585382
transform 1 0 141696 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_695
timestamp 1679585382
transform 1 0 142368 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_702
timestamp 1679585382
transform 1 0 143040 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_709
timestamp 1679585382
transform 1 0 143712 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_716
timestamp 1679585382
transform 1 0 144384 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_723
timestamp 1679585382
transform 1 0 145056 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_730
timestamp 1679585382
transform 1 0 145728 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_737
timestamp 1679585382
transform 1 0 146400 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_67_744
timestamp 1679585382
transform 1 0 147072 0 -1 127008
box -48 -56 720 834
use sg13g2_decap_4  FILLER_67_751
timestamp 1679581501
transform 1 0 147744 0 -1 127008
box -48 -56 432 834
use sg13g2_fill_2  FILLER_67_755
timestamp 1677583704
transform 1 0 148128 0 -1 127008
box -48 -56 240 834
use sg13g2_decap_8  FILLER_68_0
timestamp 1679585382
transform 1 0 75648 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_7
timestamp 1679585382
transform 1 0 76320 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_14
timestamp 1679585382
transform 1 0 76992 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_21
timestamp 1679585382
transform 1 0 77664 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_28
timestamp 1679585382
transform 1 0 78336 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_35
timestamp 1679585382
transform 1 0 79008 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_42
timestamp 1679585382
transform 1 0 79680 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_49
timestamp 1679585382
transform 1 0 80352 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_56
timestamp 1679585382
transform 1 0 81024 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_63
timestamp 1679585382
transform 1 0 81696 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_70
timestamp 1679585382
transform 1 0 82368 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_77
timestamp 1679585382
transform 1 0 83040 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_84
timestamp 1679585382
transform 1 0 83712 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_91
timestamp 1679585382
transform 1 0 84384 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_98
timestamp 1679585382
transform 1 0 85056 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_105
timestamp 1679585382
transform 1 0 85728 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_112
timestamp 1679585382
transform 1 0 86400 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_119
timestamp 1679585382
transform 1 0 87072 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_126
timestamp 1679585382
transform 1 0 87744 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_133
timestamp 1679585382
transform 1 0 88416 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_140
timestamp 1679585382
transform 1 0 89088 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_147
timestamp 1679585382
transform 1 0 89760 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_154
timestamp 1679585382
transform 1 0 90432 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_161
timestamp 1679585382
transform 1 0 91104 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_168
timestamp 1679585382
transform 1 0 91776 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_175
timestamp 1679585382
transform 1 0 92448 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_182
timestamp 1679585382
transform 1 0 93120 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_189
timestamp 1679585382
transform 1 0 93792 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_202
timestamp 1679585382
transform 1 0 95040 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_209
timestamp 1679585382
transform 1 0 95712 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_216
timestamp 1679585382
transform 1 0 96384 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_223
timestamp 1679585382
transform 1 0 97056 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_230
timestamp 1679585382
transform 1 0 97728 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_237
timestamp 1679585382
transform 1 0 98400 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_244
timestamp 1679585382
transform 1 0 99072 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_251
timestamp 1679585382
transform 1 0 99744 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_258
timestamp 1679585382
transform 1 0 100416 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_265
timestamp 1679585382
transform 1 0 101088 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_272
timestamp 1679585382
transform 1 0 101760 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_279
timestamp 1679585382
transform 1 0 102432 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_286
timestamp 1679585382
transform 1 0 103104 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_293
timestamp 1679585382
transform 1 0 103776 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_300
timestamp 1679585382
transform 1 0 104448 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_307
timestamp 1679585382
transform 1 0 105120 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_314
timestamp 1679585382
transform 1 0 105792 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_321
timestamp 1679585382
transform 1 0 106464 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_328
timestamp 1679585382
transform 1 0 107136 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_335
timestamp 1679585382
transform 1 0 107808 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_342
timestamp 1679585382
transform 1 0 108480 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_349
timestamp 1679585382
transform 1 0 109152 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_356
timestamp 1679585382
transform 1 0 109824 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_363
timestamp 1679585382
transform 1 0 110496 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_370
timestamp 1679585382
transform 1 0 111168 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_377
timestamp 1679585382
transform 1 0 111840 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_384
timestamp 1679585382
transform 1 0 112512 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_391
timestamp 1679585382
transform 1 0 113184 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_398
timestamp 1679585382
transform 1 0 113856 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_405
timestamp 1679585382
transform 1 0 114528 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_412
timestamp 1679585382
transform 1 0 115200 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_419
timestamp 1679585382
transform 1 0 115872 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_426
timestamp 1679585382
transform 1 0 116544 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_433
timestamp 1679585382
transform 1 0 117216 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_440
timestamp 1679585382
transform 1 0 117888 0 1 127008
box -48 -56 720 834
use sg13g2_fill_2  FILLER_68_447
timestamp 1677583704
transform 1 0 118560 0 1 127008
box -48 -56 240 834
use sg13g2_decap_8  FILLER_68_454
timestamp 1679585382
transform 1 0 119232 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_461
timestamp 1679585382
transform 1 0 119904 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_468
timestamp 1679585382
transform 1 0 120576 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_475
timestamp 1679585382
transform 1 0 121248 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_482
timestamp 1679585382
transform 1 0 121920 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_489
timestamp 1679585382
transform 1 0 122592 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_496
timestamp 1679585382
transform 1 0 123264 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_503
timestamp 1679585382
transform 1 0 123936 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_510
timestamp 1679585382
transform 1 0 124608 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_517
timestamp 1679585382
transform 1 0 125280 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_524
timestamp 1679585382
transform 1 0 125952 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_531
timestamp 1679585382
transform 1 0 126624 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_538
timestamp 1679585382
transform 1 0 127296 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_545
timestamp 1679585382
transform 1 0 127968 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_552
timestamp 1679585382
transform 1 0 128640 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_559
timestamp 1679585382
transform 1 0 129312 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_566
timestamp 1679585382
transform 1 0 129984 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_573
timestamp 1679585382
transform 1 0 130656 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_580
timestamp 1679585382
transform 1 0 131328 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_587
timestamp 1679585382
transform 1 0 132000 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_594
timestamp 1679585382
transform 1 0 132672 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_601
timestamp 1679585382
transform 1 0 133344 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_608
timestamp 1679585382
transform 1 0 134016 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_615
timestamp 1679585382
transform 1 0 134688 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_622
timestamp 1679585382
transform 1 0 135360 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_629
timestamp 1679585382
transform 1 0 136032 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_636
timestamp 1679585382
transform 1 0 136704 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_643
timestamp 1679585382
transform 1 0 137376 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_650
timestamp 1679585382
transform 1 0 138048 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_657
timestamp 1679585382
transform 1 0 138720 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_664
timestamp 1679585382
transform 1 0 139392 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_671
timestamp 1679585382
transform 1 0 140064 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_678
timestamp 1679585382
transform 1 0 140736 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_685
timestamp 1679585382
transform 1 0 141408 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_692
timestamp 1679585382
transform 1 0 142080 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_699
timestamp 1679585382
transform 1 0 142752 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_706
timestamp 1679585382
transform 1 0 143424 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_713
timestamp 1679585382
transform 1 0 144096 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_720
timestamp 1679585382
transform 1 0 144768 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_727
timestamp 1679585382
transform 1 0 145440 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_734
timestamp 1679585382
transform 1 0 146112 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_741
timestamp 1679585382
transform 1 0 146784 0 1 127008
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_748
timestamp 1679585382
transform 1 0 147456 0 1 127008
box -48 -56 720 834
use sg13g2_fill_2  FILLER_68_755
timestamp 1677583704
transform 1 0 148128 0 1 127008
box -48 -56 240 834
use sg13g2_decap_8  FILLER_69_0
timestamp 1679585382
transform 1 0 75648 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_7
timestamp 1679585382
transform 1 0 76320 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_14
timestamp 1679585382
transform 1 0 76992 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_21
timestamp 1679585382
transform 1 0 77664 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_28
timestamp 1679585382
transform 1 0 78336 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_35
timestamp 1679585382
transform 1 0 79008 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_42
timestamp 1679585382
transform 1 0 79680 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_49
timestamp 1679585382
transform 1 0 80352 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_56
timestamp 1679585382
transform 1 0 81024 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_63
timestamp 1679585382
transform 1 0 81696 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_70
timestamp 1679585382
transform 1 0 82368 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_77
timestamp 1679585382
transform 1 0 83040 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_84
timestamp 1679585382
transform 1 0 83712 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_91
timestamp 1679585382
transform 1 0 84384 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_98
timestamp 1679585382
transform 1 0 85056 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_105
timestamp 1679585382
transform 1 0 85728 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_112
timestamp 1679585382
transform 1 0 86400 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_119
timestamp 1679585382
transform 1 0 87072 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_126
timestamp 1679585382
transform 1 0 87744 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_133
timestamp 1679585382
transform 1 0 88416 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_140
timestamp 1679585382
transform 1 0 89088 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_147
timestamp 1679585382
transform 1 0 89760 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_154
timestamp 1679585382
transform 1 0 90432 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_161
timestamp 1679585382
transform 1 0 91104 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_168
timestamp 1679585382
transform 1 0 91776 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_175
timestamp 1679585382
transform 1 0 92448 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_182
timestamp 1679585382
transform 1 0 93120 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_189
timestamp 1679585382
transform 1 0 93792 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_196
timestamp 1679585382
transform 1 0 94464 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_203
timestamp 1679585382
transform 1 0 95136 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_210
timestamp 1679585382
transform 1 0 95808 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_217
timestamp 1679585382
transform 1 0 96480 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_224
timestamp 1679585382
transform 1 0 97152 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_231
timestamp 1679585382
transform 1 0 97824 0 -1 128520
box -48 -56 720 834
use sg13g2_fill_2  FILLER_69_238
timestamp 1677583704
transform 1 0 98496 0 -1 128520
box -48 -56 240 834
use sg13g2_fill_1  FILLER_69_240
timestamp 1677583258
transform 1 0 98688 0 -1 128520
box -48 -56 144 834
use sg13g2_decap_8  FILLER_69_247
timestamp 1679585382
transform 1 0 99360 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_254
timestamp 1679585382
transform 1 0 100032 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_261
timestamp 1679585382
transform 1 0 100704 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_268
timestamp 1679585382
transform 1 0 101376 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_275
timestamp 1679585382
transform 1 0 102048 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_282
timestamp 1679585382
transform 1 0 102720 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_289
timestamp 1679585382
transform 1 0 103392 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_296
timestamp 1679585382
transform 1 0 104064 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_303
timestamp 1679585382
transform 1 0 104736 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_310
timestamp 1679585382
transform 1 0 105408 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_317
timestamp 1679585382
transform 1 0 106080 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_324
timestamp 1679585382
transform 1 0 106752 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_331
timestamp 1679585382
transform 1 0 107424 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_338
timestamp 1679585382
transform 1 0 108096 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_345
timestamp 1679585382
transform 1 0 108768 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_352
timestamp 1679585382
transform 1 0 109440 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_359
timestamp 1679585382
transform 1 0 110112 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_366
timestamp 1679585382
transform 1 0 110784 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_373
timestamp 1679585382
transform 1 0 111456 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_380
timestamp 1679585382
transform 1 0 112128 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_387
timestamp 1679585382
transform 1 0 112800 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_394
timestamp 1679585382
transform 1 0 113472 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_401
timestamp 1679585382
transform 1 0 114144 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_408
timestamp 1679585382
transform 1 0 114816 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_415
timestamp 1679585382
transform 1 0 115488 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_422
timestamp 1679585382
transform 1 0 116160 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_429
timestamp 1679585382
transform 1 0 116832 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_436
timestamp 1679585382
transform 1 0 117504 0 -1 128520
box -48 -56 720 834
use sg13g2_fill_1  FILLER_69_456
timestamp 1677583258
transform 1 0 119424 0 -1 128520
box -48 -56 144 834
use sg13g2_decap_8  FILLER_69_462
timestamp 1679585382
transform 1 0 120000 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_496
timestamp 1679585382
transform 1 0 123264 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_503
timestamp 1679585382
transform 1 0 123936 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_510
timestamp 1679585382
transform 1 0 124608 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_517
timestamp 1679585382
transform 1 0 125280 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_524
timestamp 1679585382
transform 1 0 125952 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_531
timestamp 1679585382
transform 1 0 126624 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_538
timestamp 1679585382
transform 1 0 127296 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_545
timestamp 1679585382
transform 1 0 127968 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_552
timestamp 1679585382
transform 1 0 128640 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_559
timestamp 1679585382
transform 1 0 129312 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_566
timestamp 1679585382
transform 1 0 129984 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_573
timestamp 1679585382
transform 1 0 130656 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_580
timestamp 1679585382
transform 1 0 131328 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_587
timestamp 1679585382
transform 1 0 132000 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_594
timestamp 1679585382
transform 1 0 132672 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_601
timestamp 1679585382
transform 1 0 133344 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_608
timestamp 1679585382
transform 1 0 134016 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_615
timestamp 1679585382
transform 1 0 134688 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_622
timestamp 1679585382
transform 1 0 135360 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_629
timestamp 1679585382
transform 1 0 136032 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_636
timestamp 1679585382
transform 1 0 136704 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_643
timestamp 1679585382
transform 1 0 137376 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_650
timestamp 1679585382
transform 1 0 138048 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_657
timestamp 1679585382
transform 1 0 138720 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_664
timestamp 1679585382
transform 1 0 139392 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_671
timestamp 1679585382
transform 1 0 140064 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_678
timestamp 1679585382
transform 1 0 140736 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_685
timestamp 1679585382
transform 1 0 141408 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_692
timestamp 1679585382
transform 1 0 142080 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_699
timestamp 1679585382
transform 1 0 142752 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_706
timestamp 1679585382
transform 1 0 143424 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_713
timestamp 1679585382
transform 1 0 144096 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_720
timestamp 1679585382
transform 1 0 144768 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_727
timestamp 1679585382
transform 1 0 145440 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_734
timestamp 1679585382
transform 1 0 146112 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_741
timestamp 1679585382
transform 1 0 146784 0 -1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_748
timestamp 1679585382
transform 1 0 147456 0 -1 128520
box -48 -56 720 834
use sg13g2_fill_2  FILLER_69_755
timestamp 1677583704
transform 1 0 148128 0 -1 128520
box -48 -56 240 834
use sg13g2_decap_8  FILLER_70_0
timestamp 1679585382
transform 1 0 75648 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_7
timestamp 1679585382
transform 1 0 76320 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_14
timestamp 1679585382
transform 1 0 76992 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_21
timestamp 1679585382
transform 1 0 77664 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_28
timestamp 1679585382
transform 1 0 78336 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_35
timestamp 1679585382
transform 1 0 79008 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_42
timestamp 1679585382
transform 1 0 79680 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_49
timestamp 1679585382
transform 1 0 80352 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_56
timestamp 1679585382
transform 1 0 81024 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_63
timestamp 1679585382
transform 1 0 81696 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_70
timestamp 1679585382
transform 1 0 82368 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_77
timestamp 1679585382
transform 1 0 83040 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_84
timestamp 1679585382
transform 1 0 83712 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_91
timestamp 1679585382
transform 1 0 84384 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_98
timestamp 1679585382
transform 1 0 85056 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_105
timestamp 1679585382
transform 1 0 85728 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_112
timestamp 1679585382
transform 1 0 86400 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_119
timestamp 1679585382
transform 1 0 87072 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_126
timestamp 1679585382
transform 1 0 87744 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_133
timestamp 1679585382
transform 1 0 88416 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_140
timestamp 1679585382
transform 1 0 89088 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_147
timestamp 1679585382
transform 1 0 89760 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_154
timestamp 1679585382
transform 1 0 90432 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_161
timestamp 1679585382
transform 1 0 91104 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_168
timestamp 1679585382
transform 1 0 91776 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_175
timestamp 1679585382
transform 1 0 92448 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_182
timestamp 1679585382
transform 1 0 93120 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_195
timestamp 1679585382
transform 1 0 94368 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_202
timestamp 1679585382
transform 1 0 95040 0 1 128520
box -48 -56 720 834
use sg13g2_fill_2  FILLER_70_209
timestamp 1677583704
transform 1 0 95712 0 1 128520
box -48 -56 240 834
use sg13g2_fill_1  FILLER_70_211
timestamp 1677583258
transform 1 0 95904 0 1 128520
box -48 -56 144 834
use sg13g2_decap_8  FILLER_70_221
timestamp 1679585382
transform 1 0 96864 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_228
timestamp 1679585382
transform 1 0 97536 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_235
timestamp 1679585382
transform 1 0 98208 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_242
timestamp 1679585382
transform 1 0 98880 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_249
timestamp 1679585382
transform 1 0 99552 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_256
timestamp 1679585382
transform 1 0 100224 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_263
timestamp 1679585382
transform 1 0 100896 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_270
timestamp 1679585382
transform 1 0 101568 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_277
timestamp 1679585382
transform 1 0 102240 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_284
timestamp 1679585382
transform 1 0 102912 0 1 128520
box -48 -56 720 834
use sg13g2_decap_4  FILLER_70_291
timestamp 1679581501
transform 1 0 103584 0 1 128520
box -48 -56 432 834
use sg13g2_decap_8  FILLER_70_299
timestamp 1679585382
transform 1 0 104352 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_306
timestamp 1679585382
transform 1 0 105024 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_313
timestamp 1679585382
transform 1 0 105696 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_320
timestamp 1679585382
transform 1 0 106368 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_327
timestamp 1679585382
transform 1 0 107040 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_334
timestamp 1679585382
transform 1 0 107712 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_341
timestamp 1679585382
transform 1 0 108384 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_348
timestamp 1679585382
transform 1 0 109056 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_355
timestamp 1679585382
transform 1 0 109728 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_362
timestamp 1679585382
transform 1 0 110400 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_369
timestamp 1679585382
transform 1 0 111072 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_376
timestamp 1679585382
transform 1 0 111744 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_383
timestamp 1679585382
transform 1 0 112416 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_390
timestamp 1679585382
transform 1 0 113088 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_397
timestamp 1679585382
transform 1 0 113760 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_404
timestamp 1679585382
transform 1 0 114432 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_411
timestamp 1679585382
transform 1 0 115104 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_418
timestamp 1679585382
transform 1 0 115776 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_425
timestamp 1679585382
transform 1 0 116448 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_432
timestamp 1679585382
transform 1 0 117120 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_439
timestamp 1679585382
transform 1 0 117792 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_446
timestamp 1679585382
transform 1 0 118464 0 1 128520
box -48 -56 720 834
use sg13g2_fill_2  FILLER_70_453
timestamp 1677583704
transform 1 0 119136 0 1 128520
box -48 -56 240 834
use sg13g2_fill_1  FILLER_70_455
timestamp 1677583258
transform 1 0 119328 0 1 128520
box -48 -56 144 834
use sg13g2_fill_2  FILLER_70_478
timestamp 1677583704
transform 1 0 121536 0 1 128520
box -48 -56 240 834
use sg13g2_fill_1  FILLER_70_480
timestamp 1677583258
transform 1 0 121728 0 1 128520
box -48 -56 144 834
use sg13g2_decap_8  FILLER_70_484
timestamp 1679585382
transform 1 0 122112 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_491
timestamp 1679585382
transform 1 0 122784 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_498
timestamp 1679585382
transform 1 0 123456 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_505
timestamp 1679585382
transform 1 0 124128 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_512
timestamp 1679585382
transform 1 0 124800 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_519
timestamp 1679585382
transform 1 0 125472 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_526
timestamp 1679585382
transform 1 0 126144 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_533
timestamp 1679585382
transform 1 0 126816 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_540
timestamp 1679585382
transform 1 0 127488 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_547
timestamp 1679585382
transform 1 0 128160 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_554
timestamp 1679585382
transform 1 0 128832 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_561
timestamp 1679585382
transform 1 0 129504 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_568
timestamp 1679585382
transform 1 0 130176 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_575
timestamp 1679585382
transform 1 0 130848 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_582
timestamp 1679585382
transform 1 0 131520 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_589
timestamp 1679585382
transform 1 0 132192 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_596
timestamp 1679585382
transform 1 0 132864 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_603
timestamp 1679585382
transform 1 0 133536 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_610
timestamp 1679585382
transform 1 0 134208 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_617
timestamp 1679585382
transform 1 0 134880 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_624
timestamp 1679585382
transform 1 0 135552 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_631
timestamp 1679585382
transform 1 0 136224 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_638
timestamp 1679585382
transform 1 0 136896 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_645
timestamp 1679585382
transform 1 0 137568 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_652
timestamp 1679585382
transform 1 0 138240 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_659
timestamp 1679585382
transform 1 0 138912 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_666
timestamp 1679585382
transform 1 0 139584 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_673
timestamp 1679585382
transform 1 0 140256 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_680
timestamp 1679585382
transform 1 0 140928 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_687
timestamp 1679585382
transform 1 0 141600 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_694
timestamp 1679585382
transform 1 0 142272 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_701
timestamp 1679585382
transform 1 0 142944 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_708
timestamp 1679585382
transform 1 0 143616 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_715
timestamp 1679585382
transform 1 0 144288 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_722
timestamp 1679585382
transform 1 0 144960 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_729
timestamp 1679585382
transform 1 0 145632 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_736
timestamp 1679585382
transform 1 0 146304 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_743
timestamp 1679585382
transform 1 0 146976 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_70_750
timestamp 1679585382
transform 1 0 147648 0 1 128520
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_0
timestamp 1679585382
transform 1 0 75648 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_7
timestamp 1679585382
transform 1 0 76320 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_14
timestamp 1679585382
transform 1 0 76992 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_21
timestamp 1679585382
transform 1 0 77664 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_28
timestamp 1679585382
transform 1 0 78336 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_35
timestamp 1679585382
transform 1 0 79008 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_42
timestamp 1679585382
transform 1 0 79680 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_49
timestamp 1679585382
transform 1 0 80352 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_56
timestamp 1679585382
transform 1 0 81024 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_63
timestamp 1679585382
transform 1 0 81696 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_70
timestamp 1679585382
transform 1 0 82368 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_77
timestamp 1679585382
transform 1 0 83040 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_84
timestamp 1679585382
transform 1 0 83712 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_91
timestamp 1679585382
transform 1 0 84384 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_98
timestamp 1679585382
transform 1 0 85056 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_105
timestamp 1679585382
transform 1 0 85728 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_112
timestamp 1679585382
transform 1 0 86400 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_119
timestamp 1679585382
transform 1 0 87072 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_126
timestamp 1679585382
transform 1 0 87744 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_133
timestamp 1679585382
transform 1 0 88416 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_140
timestamp 1679585382
transform 1 0 89088 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_147
timestamp 1679585382
transform 1 0 89760 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_154
timestamp 1679585382
transform 1 0 90432 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_161
timestamp 1679585382
transform 1 0 91104 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_168
timestamp 1679585382
transform 1 0 91776 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_175
timestamp 1679585382
transform 1 0 92448 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_182
timestamp 1679585382
transform 1 0 93120 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_189
timestamp 1679585382
transform 1 0 93792 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_196
timestamp 1679585382
transform 1 0 94464 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_203
timestamp 1679585382
transform 1 0 95136 0 -1 130032
box -48 -56 720 834
use sg13g2_fill_2  FILLER_71_210
timestamp 1677583704
transform 1 0 95808 0 -1 130032
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_212
timestamp 1677583258
transform 1 0 96000 0 -1 130032
box -48 -56 144 834
use sg13g2_fill_1  FILLER_71_222
timestamp 1677583258
transform 1 0 96960 0 -1 130032
box -48 -56 144 834
use sg13g2_decap_8  FILLER_71_228
timestamp 1679585382
transform 1 0 97536 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_235
timestamp 1679585382
transform 1 0 98208 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_242
timestamp 1679585382
transform 1 0 98880 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_249
timestamp 1679585382
transform 1 0 99552 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_256
timestamp 1679585382
transform 1 0 100224 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_263
timestamp 1679585382
transform 1 0 100896 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_270
timestamp 1679585382
transform 1 0 101568 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_277
timestamp 1679585382
transform 1 0 102240 0 -1 130032
box -48 -56 720 834
use sg13g2_fill_1  FILLER_71_284
timestamp 1677583258
transform 1 0 102912 0 -1 130032
box -48 -56 144 834
use sg13g2_fill_1  FILLER_71_289
timestamp 1677583258
transform 1 0 103392 0 -1 130032
box -48 -56 144 834
use sg13g2_decap_8  FILLER_71_317
timestamp 1679585382
transform 1 0 106080 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_324
timestamp 1679585382
transform 1 0 106752 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_331
timestamp 1679585382
transform 1 0 107424 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_338
timestamp 1679585382
transform 1 0 108096 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_345
timestamp 1679585382
transform 1 0 108768 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_352
timestamp 1679585382
transform 1 0 109440 0 -1 130032
box -48 -56 720 834
use sg13g2_fill_2  FILLER_71_359
timestamp 1677583704
transform 1 0 110112 0 -1 130032
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_361
timestamp 1677583258
transform 1 0 110304 0 -1 130032
box -48 -56 144 834
use sg13g2_decap_8  FILLER_71_387
timestamp 1679585382
transform 1 0 112800 0 -1 130032
box -48 -56 720 834
use sg13g2_fill_2  FILLER_71_394
timestamp 1677583704
transform 1 0 113472 0 -1 130032
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_396
timestamp 1677583258
transform 1 0 113664 0 -1 130032
box -48 -56 144 834
use sg13g2_decap_8  FILLER_71_422
timestamp 1679585382
transform 1 0 116160 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_429
timestamp 1679585382
transform 1 0 116832 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_436
timestamp 1679585382
transform 1 0 117504 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_443
timestamp 1679585382
transform 1 0 118176 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_450
timestamp 1679585382
transform 1 0 118848 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_457
timestamp 1679585382
transform 1 0 119520 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_464
timestamp 1679585382
transform 1 0 120192 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_471
timestamp 1679585382
transform 1 0 120864 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_478
timestamp 1679585382
transform 1 0 121536 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_485
timestamp 1679585382
transform 1 0 122208 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_492
timestamp 1679585382
transform 1 0 122880 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_499
timestamp 1679585382
transform 1 0 123552 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_506
timestamp 1679585382
transform 1 0 124224 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_513
timestamp 1679585382
transform 1 0 124896 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_520
timestamp 1679585382
transform 1 0 125568 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_527
timestamp 1679585382
transform 1 0 126240 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_534
timestamp 1679585382
transform 1 0 126912 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_541
timestamp 1679585382
transform 1 0 127584 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_548
timestamp 1679585382
transform 1 0 128256 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_555
timestamp 1679585382
transform 1 0 128928 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_562
timestamp 1679585382
transform 1 0 129600 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_569
timestamp 1679585382
transform 1 0 130272 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_576
timestamp 1679585382
transform 1 0 130944 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_583
timestamp 1679585382
transform 1 0 131616 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_590
timestamp 1679585382
transform 1 0 132288 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_597
timestamp 1679585382
transform 1 0 132960 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_604
timestamp 1679585382
transform 1 0 133632 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_611
timestamp 1679585382
transform 1 0 134304 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_618
timestamp 1679585382
transform 1 0 134976 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_625
timestamp 1679585382
transform 1 0 135648 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_632
timestamp 1679585382
transform 1 0 136320 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_639
timestamp 1679585382
transform 1 0 136992 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_646
timestamp 1679585382
transform 1 0 137664 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_653
timestamp 1679585382
transform 1 0 138336 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_660
timestamp 1679585382
transform 1 0 139008 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_667
timestamp 1679585382
transform 1 0 139680 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_674
timestamp 1679585382
transform 1 0 140352 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_681
timestamp 1679585382
transform 1 0 141024 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_688
timestamp 1679585382
transform 1 0 141696 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_695
timestamp 1679585382
transform 1 0 142368 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_702
timestamp 1679585382
transform 1 0 143040 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_709
timestamp 1679585382
transform 1 0 143712 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_716
timestamp 1679585382
transform 1 0 144384 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_723
timestamp 1679585382
transform 1 0 145056 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_730
timestamp 1679585382
transform 1 0 145728 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_737
timestamp 1679585382
transform 1 0 146400 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_744
timestamp 1679585382
transform 1 0 147072 0 -1 130032
box -48 -56 720 834
use sg13g2_decap_4  FILLER_71_751
timestamp 1679581501
transform 1 0 147744 0 -1 130032
box -48 -56 432 834
use sg13g2_fill_2  FILLER_71_755
timestamp 1677583704
transform 1 0 148128 0 -1 130032
box -48 -56 240 834
use sg13g2_decap_8  FILLER_72_0
timestamp 1679585382
transform 1 0 75648 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_7
timestamp 1679585382
transform 1 0 76320 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_14
timestamp 1679585382
transform 1 0 76992 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_21
timestamp 1679585382
transform 1 0 77664 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_28
timestamp 1679585382
transform 1 0 78336 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_35
timestamp 1679585382
transform 1 0 79008 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_42
timestamp 1679585382
transform 1 0 79680 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_49
timestamp 1679585382
transform 1 0 80352 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_56
timestamp 1679585382
transform 1 0 81024 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_63
timestamp 1679585382
transform 1 0 81696 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_70
timestamp 1679585382
transform 1 0 82368 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_77
timestamp 1679585382
transform 1 0 83040 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_84
timestamp 1679585382
transform 1 0 83712 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_91
timestamp 1679585382
transform 1 0 84384 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_98
timestamp 1679585382
transform 1 0 85056 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_105
timestamp 1679585382
transform 1 0 85728 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_112
timestamp 1679585382
transform 1 0 86400 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_119
timestamp 1679585382
transform 1 0 87072 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_126
timestamp 1679585382
transform 1 0 87744 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_133
timestamp 1679585382
transform 1 0 88416 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_140
timestamp 1679585382
transform 1 0 89088 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_147
timestamp 1679585382
transform 1 0 89760 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_154
timestamp 1679585382
transform 1 0 90432 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_161
timestamp 1679585382
transform 1 0 91104 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_168
timestamp 1679585382
transform 1 0 91776 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_175
timestamp 1679585382
transform 1 0 92448 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_182
timestamp 1679585382
transform 1 0 93120 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_189
timestamp 1679585382
transform 1 0 93792 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_196
timestamp 1679585382
transform 1 0 94464 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_203
timestamp 1679585382
transform 1 0 95136 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_210
timestamp 1679585382
transform 1 0 95808 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_217
timestamp 1679585382
transform 1 0 96480 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_224
timestamp 1679585382
transform 1 0 97152 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_235
timestamp 1679585382
transform 1 0 98208 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_242
timestamp 1679585382
transform 1 0 98880 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_249
timestamp 1679585382
transform 1 0 99552 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_256
timestamp 1679585382
transform 1 0 100224 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_263
timestamp 1679585382
transform 1 0 100896 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_270
timestamp 1679585382
transform 1 0 101568 0 1 130032
box -48 -56 720 834
use sg13g2_fill_2  FILLER_72_277
timestamp 1677583704
transform 1 0 102240 0 1 130032
box -48 -56 240 834
use sg13g2_decap_8  FILLER_72_287
timestamp 1679585382
transform 1 0 103200 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_294
timestamp 1679585382
transform 1 0 103872 0 1 130032
box -48 -56 720 834
use sg13g2_fill_1  FILLER_72_301
timestamp 1677583258
transform 1 0 104544 0 1 130032
box -48 -56 144 834
use sg13g2_decap_8  FILLER_72_311
timestamp 1679585382
transform 1 0 105504 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_318
timestamp 1679585382
transform 1 0 106176 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_325
timestamp 1679585382
transform 1 0 106848 0 1 130032
box -48 -56 720 834
use sg13g2_decap_4  FILLER_72_332
timestamp 1679581501
transform 1 0 107520 0 1 130032
box -48 -56 432 834
use sg13g2_fill_1  FILLER_72_336
timestamp 1677583258
transform 1 0 107904 0 1 130032
box -48 -56 144 834
use sg13g2_decap_8  FILLER_72_367
timestamp 1679585382
transform 1 0 110880 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_374
timestamp 1679585382
transform 1 0 111552 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_381
timestamp 1679585382
transform 1 0 112224 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_388
timestamp 1679585382
transform 1 0 112896 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_395
timestamp 1679585382
transform 1 0 113568 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_402
timestamp 1679585382
transform 1 0 114240 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_409
timestamp 1679585382
transform 1 0 114912 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_416
timestamp 1679585382
transform 1 0 115584 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_423
timestamp 1679585382
transform 1 0 116256 0 1 130032
box -48 -56 720 834
use sg13g2_decap_4  FILLER_72_430
timestamp 1679581501
transform 1 0 116928 0 1 130032
box -48 -56 432 834
use sg13g2_fill_1  FILLER_72_434
timestamp 1677583258
transform 1 0 117312 0 1 130032
box -48 -56 144 834
use sg13g2_decap_8  FILLER_72_439
timestamp 1679585382
transform 1 0 117792 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_446
timestamp 1679585382
transform 1 0 118464 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_453
timestamp 1679585382
transform 1 0 119136 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_460
timestamp 1679585382
transform 1 0 119808 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_467
timestamp 1679585382
transform 1 0 120480 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_474
timestamp 1679585382
transform 1 0 121152 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_481
timestamp 1679585382
transform 1 0 121824 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_488
timestamp 1679585382
transform 1 0 122496 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_495
timestamp 1679585382
transform 1 0 123168 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_502
timestamp 1679585382
transform 1 0 123840 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_509
timestamp 1679585382
transform 1 0 124512 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_516
timestamp 1679585382
transform 1 0 125184 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_523
timestamp 1679585382
transform 1 0 125856 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_530
timestamp 1679585382
transform 1 0 126528 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_537
timestamp 1679585382
transform 1 0 127200 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_544
timestamp 1679585382
transform 1 0 127872 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_551
timestamp 1679585382
transform 1 0 128544 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_558
timestamp 1679585382
transform 1 0 129216 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_565
timestamp 1679585382
transform 1 0 129888 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_572
timestamp 1679585382
transform 1 0 130560 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_579
timestamp 1679585382
transform 1 0 131232 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_586
timestamp 1679585382
transform 1 0 131904 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_593
timestamp 1679585382
transform 1 0 132576 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_600
timestamp 1679585382
transform 1 0 133248 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_607
timestamp 1679585382
transform 1 0 133920 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_614
timestamp 1679585382
transform 1 0 134592 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_621
timestamp 1679585382
transform 1 0 135264 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_628
timestamp 1679585382
transform 1 0 135936 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_635
timestamp 1679585382
transform 1 0 136608 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_642
timestamp 1679585382
transform 1 0 137280 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_649
timestamp 1679585382
transform 1 0 137952 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_656
timestamp 1679585382
transform 1 0 138624 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_663
timestamp 1679585382
transform 1 0 139296 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_670
timestamp 1679585382
transform 1 0 139968 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_677
timestamp 1679585382
transform 1 0 140640 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_684
timestamp 1679585382
transform 1 0 141312 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_691
timestamp 1679585382
transform 1 0 141984 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_698
timestamp 1679585382
transform 1 0 142656 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_705
timestamp 1679585382
transform 1 0 143328 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_712
timestamp 1679585382
transform 1 0 144000 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_719
timestamp 1679585382
transform 1 0 144672 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_726
timestamp 1679585382
transform 1 0 145344 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_733
timestamp 1679585382
transform 1 0 146016 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_740
timestamp 1679585382
transform 1 0 146688 0 1 130032
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_747
timestamp 1679585382
transform 1 0 147360 0 1 130032
box -48 -56 720 834
use sg13g2_fill_2  FILLER_72_754
timestamp 1677583704
transform 1 0 148032 0 1 130032
box -48 -56 240 834
use sg13g2_fill_1  FILLER_72_756
timestamp 1677583258
transform 1 0 148224 0 1 130032
box -48 -56 144 834
use sg13g2_decap_8  FILLER_73_0
timestamp 1679585382
transform 1 0 75648 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_7
timestamp 1679585382
transform 1 0 76320 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_14
timestamp 1679585382
transform 1 0 76992 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_21
timestamp 1679585382
transform 1 0 77664 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_28
timestamp 1679585382
transform 1 0 78336 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_35
timestamp 1679585382
transform 1 0 79008 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_42
timestamp 1679585382
transform 1 0 79680 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_49
timestamp 1679585382
transform 1 0 80352 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_56
timestamp 1679585382
transform 1 0 81024 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_63
timestamp 1679585382
transform 1 0 81696 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_70
timestamp 1679585382
transform 1 0 82368 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_77
timestamp 1679585382
transform 1 0 83040 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_84
timestamp 1679585382
transform 1 0 83712 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_91
timestamp 1679585382
transform 1 0 84384 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_98
timestamp 1679585382
transform 1 0 85056 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_105
timestamp 1679585382
transform 1 0 85728 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_112
timestamp 1679585382
transform 1 0 86400 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_119
timestamp 1679585382
transform 1 0 87072 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_126
timestamp 1679585382
transform 1 0 87744 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_133
timestamp 1679585382
transform 1 0 88416 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_140
timestamp 1679585382
transform 1 0 89088 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_147
timestamp 1679585382
transform 1 0 89760 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_154
timestamp 1679585382
transform 1 0 90432 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_161
timestamp 1679585382
transform 1 0 91104 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_168
timestamp 1679585382
transform 1 0 91776 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_175
timestamp 1679585382
transform 1 0 92448 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_182
timestamp 1679585382
transform 1 0 93120 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_189
timestamp 1679585382
transform 1 0 93792 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_196
timestamp 1679585382
transform 1 0 94464 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_203
timestamp 1679585382
transform 1 0 95136 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_210
timestamp 1679585382
transform 1 0 95808 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_217
timestamp 1679585382
transform 1 0 96480 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_224
timestamp 1679585382
transform 1 0 97152 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_231
timestamp 1679585382
transform 1 0 97824 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_238
timestamp 1679585382
transform 1 0 98496 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_245
timestamp 1679585382
transform 1 0 99168 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_261
timestamp 1679585382
transform 1 0 100704 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_4  FILLER_73_268
timestamp 1679581501
transform 1 0 101376 0 -1 131544
box -48 -56 432 834
use sg13g2_fill_2  FILLER_73_272
timestamp 1677583704
transform 1 0 101760 0 -1 131544
box -48 -56 240 834
use sg13g2_decap_8  FILLER_73_297
timestamp 1679585382
transform 1 0 104160 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_304
timestamp 1679585382
transform 1 0 104832 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_311
timestamp 1679585382
transform 1 0 105504 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_318
timestamp 1679585382
transform 1 0 106176 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_325
timestamp 1679585382
transform 1 0 106848 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_332
timestamp 1679585382
transform 1 0 107520 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_4  FILLER_73_339
timestamp 1679581501
transform 1 0 108192 0 -1 131544
box -48 -56 432 834
use sg13g2_fill_2  FILLER_73_343
timestamp 1677583704
transform 1 0 108576 0 -1 131544
box -48 -56 240 834
use sg13g2_fill_1  FILLER_73_364
timestamp 1677583258
transform 1 0 110592 0 -1 131544
box -48 -56 144 834
use sg13g2_decap_8  FILLER_73_374
timestamp 1679585382
transform 1 0 111552 0 -1 131544
box -48 -56 720 834
use sg13g2_fill_1  FILLER_73_386
timestamp 1677583258
transform 1 0 112704 0 -1 131544
box -48 -56 144 834
use sg13g2_decap_8  FILLER_73_394
timestamp 1679585382
transform 1 0 113472 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_401
timestamp 1679585382
transform 1 0 114144 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_414
timestamp 1679585382
transform 1 0 115392 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_421
timestamp 1679585382
transform 1 0 116064 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_428
timestamp 1679585382
transform 1 0 116736 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_435
timestamp 1679585382
transform 1 0 117408 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_442
timestamp 1679585382
transform 1 0 118080 0 -1 131544
box -48 -56 720 834
use sg13g2_fill_2  FILLER_73_449
timestamp 1677583704
transform 1 0 118752 0 -1 131544
box -48 -56 240 834
use sg13g2_fill_1  FILLER_73_451
timestamp 1677583258
transform 1 0 118944 0 -1 131544
box -48 -56 144 834
use sg13g2_decap_8  FILLER_73_457
timestamp 1679585382
transform 1 0 119520 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_464
timestamp 1679585382
transform 1 0 120192 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_471
timestamp 1679585382
transform 1 0 120864 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_478
timestamp 1679585382
transform 1 0 121536 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_485
timestamp 1679585382
transform 1 0 122208 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_492
timestamp 1679585382
transform 1 0 122880 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_499
timestamp 1679585382
transform 1 0 123552 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_506
timestamp 1679585382
transform 1 0 124224 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_513
timestamp 1679585382
transform 1 0 124896 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_520
timestamp 1679585382
transform 1 0 125568 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_527
timestamp 1679585382
transform 1 0 126240 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_534
timestamp 1679585382
transform 1 0 126912 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_541
timestamp 1679585382
transform 1 0 127584 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_548
timestamp 1679585382
transform 1 0 128256 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_555
timestamp 1679585382
transform 1 0 128928 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_562
timestamp 1679585382
transform 1 0 129600 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_569
timestamp 1679585382
transform 1 0 130272 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_576
timestamp 1679585382
transform 1 0 130944 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_583
timestamp 1679585382
transform 1 0 131616 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_590
timestamp 1679585382
transform 1 0 132288 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_597
timestamp 1679585382
transform 1 0 132960 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_604
timestamp 1679585382
transform 1 0 133632 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_611
timestamp 1679585382
transform 1 0 134304 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_618
timestamp 1679585382
transform 1 0 134976 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_625
timestamp 1679585382
transform 1 0 135648 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_632
timestamp 1679585382
transform 1 0 136320 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_639
timestamp 1679585382
transform 1 0 136992 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_646
timestamp 1679585382
transform 1 0 137664 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_653
timestamp 1679585382
transform 1 0 138336 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_660
timestamp 1679585382
transform 1 0 139008 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_667
timestamp 1679585382
transform 1 0 139680 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_674
timestamp 1679585382
transform 1 0 140352 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_681
timestamp 1679585382
transform 1 0 141024 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_688
timestamp 1679585382
transform 1 0 141696 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_695
timestamp 1679585382
transform 1 0 142368 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_702
timestamp 1679585382
transform 1 0 143040 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_709
timestamp 1679585382
transform 1 0 143712 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_716
timestamp 1679585382
transform 1 0 144384 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_723
timestamp 1679585382
transform 1 0 145056 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_730
timestamp 1679585382
transform 1 0 145728 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_737
timestamp 1679585382
transform 1 0 146400 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_73_744
timestamp 1679585382
transform 1 0 147072 0 -1 131544
box -48 -56 720 834
use sg13g2_decap_4  FILLER_73_751
timestamp 1679581501
transform 1 0 147744 0 -1 131544
box -48 -56 432 834
use sg13g2_fill_2  FILLER_73_755
timestamp 1677583704
transform 1 0 148128 0 -1 131544
box -48 -56 240 834
use sg13g2_decap_8  FILLER_74_0
timestamp 1679585382
transform 1 0 75648 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_7
timestamp 1679585382
transform 1 0 76320 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_14
timestamp 1679585382
transform 1 0 76992 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_21
timestamp 1679585382
transform 1 0 77664 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_28
timestamp 1679585382
transform 1 0 78336 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_35
timestamp 1679585382
transform 1 0 79008 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_42
timestamp 1679585382
transform 1 0 79680 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_49
timestamp 1679585382
transform 1 0 80352 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_56
timestamp 1679585382
transform 1 0 81024 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_63
timestamp 1679585382
transform 1 0 81696 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_70
timestamp 1679585382
transform 1 0 82368 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_77
timestamp 1679585382
transform 1 0 83040 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_84
timestamp 1679585382
transform 1 0 83712 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_91
timestamp 1679585382
transform 1 0 84384 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_98
timestamp 1679585382
transform 1 0 85056 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_105
timestamp 1679585382
transform 1 0 85728 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_112
timestamp 1679585382
transform 1 0 86400 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_119
timestamp 1679585382
transform 1 0 87072 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_126
timestamp 1679585382
transform 1 0 87744 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_133
timestamp 1679585382
transform 1 0 88416 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_140
timestamp 1679585382
transform 1 0 89088 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_147
timestamp 1679585382
transform 1 0 89760 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_154
timestamp 1679585382
transform 1 0 90432 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_161
timestamp 1679585382
transform 1 0 91104 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_168
timestamp 1679585382
transform 1 0 91776 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_175
timestamp 1679585382
transform 1 0 92448 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_182
timestamp 1679585382
transform 1 0 93120 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_189
timestamp 1679585382
transform 1 0 93792 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_196
timestamp 1679585382
transform 1 0 94464 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_203
timestamp 1679585382
transform 1 0 95136 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_210
timestamp 1679585382
transform 1 0 95808 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_217
timestamp 1679585382
transform 1 0 96480 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_224
timestamp 1679585382
transform 1 0 97152 0 1 131544
box -48 -56 720 834
use sg13g2_decap_4  FILLER_74_231
timestamp 1679581501
transform 1 0 97824 0 1 131544
box -48 -56 432 834
use sg13g2_fill_1  FILLER_74_235
timestamp 1677583258
transform 1 0 98208 0 1 131544
box -48 -56 144 834
use sg13g2_fill_2  FILLER_74_250
timestamp 1677583704
transform 1 0 99648 0 1 131544
box -48 -56 240 834
use sg13g2_fill_1  FILLER_74_252
timestamp 1677583258
transform 1 0 99840 0 1 131544
box -48 -56 144 834
use sg13g2_decap_8  FILLER_74_257
timestamp 1679585382
transform 1 0 100320 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_272
timestamp 1679585382
transform 1 0 101760 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_279
timestamp 1679585382
transform 1 0 102432 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_286
timestamp 1679585382
transform 1 0 103104 0 1 131544
box -48 -56 720 834
use sg13g2_decap_4  FILLER_74_293
timestamp 1679581501
transform 1 0 103776 0 1 131544
box -48 -56 432 834
use sg13g2_fill_1  FILLER_74_297
timestamp 1677583258
transform 1 0 104160 0 1 131544
box -48 -56 144 834
use sg13g2_decap_8  FILLER_74_302
timestamp 1679585382
transform 1 0 104640 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_309
timestamp 1679585382
transform 1 0 105312 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_316
timestamp 1679585382
transform 1 0 105984 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_323
timestamp 1679585382
transform 1 0 106656 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_330
timestamp 1679585382
transform 1 0 107328 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_337
timestamp 1679585382
transform 1 0 108000 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_344
timestamp 1679585382
transform 1 0 108672 0 1 131544
box -48 -56 720 834
use sg13g2_fill_2  FILLER_74_378
timestamp 1677583704
transform 1 0 111936 0 1 131544
box -48 -56 240 834
use sg13g2_decap_8  FILLER_74_395
timestamp 1679585382
transform 1 0 113568 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_402
timestamp 1679585382
transform 1 0 114240 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_409
timestamp 1679585382
transform 1 0 114912 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_416
timestamp 1679585382
transform 1 0 115584 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_423
timestamp 1679585382
transform 1 0 116256 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_430
timestamp 1679585382
transform 1 0 116928 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_437
timestamp 1679585382
transform 1 0 117600 0 1 131544
box -48 -56 720 834
use sg13g2_fill_1  FILLER_74_444
timestamp 1677583258
transform 1 0 118272 0 1 131544
box -48 -56 144 834
use sg13g2_decap_8  FILLER_74_448
timestamp 1679585382
transform 1 0 118656 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_455
timestamp 1679585382
transform 1 0 119328 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_462
timestamp 1679585382
transform 1 0 120000 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_469
timestamp 1679585382
transform 1 0 120672 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_476
timestamp 1679585382
transform 1 0 121344 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_483
timestamp 1679585382
transform 1 0 122016 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_490
timestamp 1679585382
transform 1 0 122688 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_497
timestamp 1679585382
transform 1 0 123360 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_504
timestamp 1679585382
transform 1 0 124032 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_511
timestamp 1679585382
transform 1 0 124704 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_518
timestamp 1679585382
transform 1 0 125376 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_525
timestamp 1679585382
transform 1 0 126048 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_532
timestamp 1679585382
transform 1 0 126720 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_539
timestamp 1679585382
transform 1 0 127392 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_546
timestamp 1679585382
transform 1 0 128064 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_553
timestamp 1679585382
transform 1 0 128736 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_560
timestamp 1679585382
transform 1 0 129408 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_567
timestamp 1679585382
transform 1 0 130080 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_574
timestamp 1679585382
transform 1 0 130752 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_581
timestamp 1679585382
transform 1 0 131424 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_588
timestamp 1679585382
transform 1 0 132096 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_595
timestamp 1679585382
transform 1 0 132768 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_602
timestamp 1679585382
transform 1 0 133440 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_609
timestamp 1679585382
transform 1 0 134112 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_616
timestamp 1679585382
transform 1 0 134784 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_623
timestamp 1679585382
transform 1 0 135456 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_630
timestamp 1679585382
transform 1 0 136128 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_637
timestamp 1679585382
transform 1 0 136800 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_644
timestamp 1679585382
transform 1 0 137472 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_651
timestamp 1679585382
transform 1 0 138144 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_658
timestamp 1679585382
transform 1 0 138816 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_665
timestamp 1679585382
transform 1 0 139488 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_672
timestamp 1679585382
transform 1 0 140160 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_679
timestamp 1679585382
transform 1 0 140832 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_686
timestamp 1679585382
transform 1 0 141504 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_693
timestamp 1679585382
transform 1 0 142176 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_700
timestamp 1679585382
transform 1 0 142848 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_707
timestamp 1679585382
transform 1 0 143520 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_714
timestamp 1679585382
transform 1 0 144192 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_721
timestamp 1679585382
transform 1 0 144864 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_728
timestamp 1679585382
transform 1 0 145536 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_735
timestamp 1679585382
transform 1 0 146208 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_742
timestamp 1679585382
transform 1 0 146880 0 1 131544
box -48 -56 720 834
use sg13g2_decap_8  FILLER_74_749
timestamp 1679585382
transform 1 0 147552 0 1 131544
box -48 -56 720 834
use sg13g2_fill_1  FILLER_74_756
timestamp 1677583258
transform 1 0 148224 0 1 131544
box -48 -56 144 834
use sg13g2_decap_8  FILLER_75_0
timestamp 1679585382
transform 1 0 75648 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_7
timestamp 1679585382
transform 1 0 76320 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_14
timestamp 1679585382
transform 1 0 76992 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_21
timestamp 1679585382
transform 1 0 77664 0 -1 133056
box -48 -56 720 834
use sg13g2_fill_2  FILLER_75_28
timestamp 1677583704
transform 1 0 78336 0 -1 133056
box -48 -56 240 834
use sg13g2_decap_8  FILLER_75_39
timestamp 1679585382
transform 1 0 79392 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_46
timestamp 1679585382
transform 1 0 80064 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_53
timestamp 1679585382
transform 1 0 80736 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_60
timestamp 1679585382
transform 1 0 81408 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_67
timestamp 1679585382
transform 1 0 82080 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_74
timestamp 1679585382
transform 1 0 82752 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_81
timestamp 1679585382
transform 1 0 83424 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_88
timestamp 1679585382
transform 1 0 84096 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_95
timestamp 1679585382
transform 1 0 84768 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_102
timestamp 1679585382
transform 1 0 85440 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_109
timestamp 1679585382
transform 1 0 86112 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_116
timestamp 1679585382
transform 1 0 86784 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_123
timestamp 1679585382
transform 1 0 87456 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_130
timestamp 1679585382
transform 1 0 88128 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_137
timestamp 1679585382
transform 1 0 88800 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_144
timestamp 1679585382
transform 1 0 89472 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_151
timestamp 1679585382
transform 1 0 90144 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_158
timestamp 1679585382
transform 1 0 90816 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_165
timestamp 1679585382
transform 1 0 91488 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_172
timestamp 1679585382
transform 1 0 92160 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_179
timestamp 1679585382
transform 1 0 92832 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_186
timestamp 1679585382
transform 1 0 93504 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_193
timestamp 1679585382
transform 1 0 94176 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_200
timestamp 1679585382
transform 1 0 94848 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_207
timestamp 1679585382
transform 1 0 95520 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_214
timestamp 1679585382
transform 1 0 96192 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_221
timestamp 1679585382
transform 1 0 96864 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_228
timestamp 1679585382
transform 1 0 97536 0 -1 133056
box -48 -56 720 834
use sg13g2_fill_2  FILLER_75_235
timestamp 1677583704
transform 1 0 98208 0 -1 133056
box -48 -56 240 834
use sg13g2_fill_1  FILLER_75_237
timestamp 1677583258
transform 1 0 98400 0 -1 133056
box -48 -56 144 834
use sg13g2_decap_8  FILLER_75_243
timestamp 1679585382
transform 1 0 98976 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_250
timestamp 1679585382
transform 1 0 99648 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_257
timestamp 1679585382
transform 1 0 100320 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_264
timestamp 1679585382
transform 1 0 100992 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_271
timestamp 1679585382
transform 1 0 101664 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_4  FILLER_75_278
timestamp 1679581501
transform 1 0 102336 0 -1 133056
box -48 -56 432 834
use sg13g2_fill_2  FILLER_75_282
timestamp 1677583704
transform 1 0 102720 0 -1 133056
box -48 -56 240 834
use sg13g2_decap_8  FILLER_75_320
timestamp 1679585382
transform 1 0 106368 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_327
timestamp 1679585382
transform 1 0 107040 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_334
timestamp 1679585382
transform 1 0 107712 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_341
timestamp 1679585382
transform 1 0 108384 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_348
timestamp 1679585382
transform 1 0 109056 0 -1 133056
box -48 -56 720 834
use sg13g2_fill_1  FILLER_75_355
timestamp 1677583258
transform 1 0 109728 0 -1 133056
box -48 -56 144 834
use sg13g2_decap_8  FILLER_75_360
timestamp 1679585382
transform 1 0 110208 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_367
timestamp 1679585382
transform 1 0 110880 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_374
timestamp 1679585382
transform 1 0 111552 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_381
timestamp 1679585382
transform 1 0 112224 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_388
timestamp 1679585382
transform 1 0 112896 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_395
timestamp 1679585382
transform 1 0 113568 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_402
timestamp 1679585382
transform 1 0 114240 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_409
timestamp 1679585382
transform 1 0 114912 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_416
timestamp 1679585382
transform 1 0 115584 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_423
timestamp 1679585382
transform 1 0 116256 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_430
timestamp 1679585382
transform 1 0 116928 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_437
timestamp 1679585382
transform 1 0 117600 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_444
timestamp 1679585382
transform 1 0 118272 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_4  FILLER_75_451
timestamp 1679581501
transform 1 0 118944 0 -1 133056
box -48 -56 432 834
use sg13g2_decap_8  FILLER_75_473
timestamp 1679585382
transform 1 0 121056 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_480
timestamp 1679585382
transform 1 0 121728 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_487
timestamp 1679585382
transform 1 0 122400 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_494
timestamp 1679585382
transform 1 0 123072 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_501
timestamp 1679585382
transform 1 0 123744 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_508
timestamp 1679585382
transform 1 0 124416 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_515
timestamp 1679585382
transform 1 0 125088 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_522
timestamp 1679585382
transform 1 0 125760 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_529
timestamp 1679585382
transform 1 0 126432 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_536
timestamp 1679585382
transform 1 0 127104 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_543
timestamp 1679585382
transform 1 0 127776 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_550
timestamp 1679585382
transform 1 0 128448 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_557
timestamp 1679585382
transform 1 0 129120 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_564
timestamp 1679585382
transform 1 0 129792 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_571
timestamp 1679585382
transform 1 0 130464 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_578
timestamp 1679585382
transform 1 0 131136 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_585
timestamp 1679585382
transform 1 0 131808 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_592
timestamp 1679585382
transform 1 0 132480 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_599
timestamp 1679585382
transform 1 0 133152 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_606
timestamp 1679585382
transform 1 0 133824 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_613
timestamp 1679585382
transform 1 0 134496 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_620
timestamp 1679585382
transform 1 0 135168 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_627
timestamp 1679585382
transform 1 0 135840 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_634
timestamp 1679585382
transform 1 0 136512 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_641
timestamp 1679585382
transform 1 0 137184 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_648
timestamp 1679585382
transform 1 0 137856 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_655
timestamp 1679585382
transform 1 0 138528 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_662
timestamp 1679585382
transform 1 0 139200 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_669
timestamp 1679585382
transform 1 0 139872 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_676
timestamp 1679585382
transform 1 0 140544 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_683
timestamp 1679585382
transform 1 0 141216 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_690
timestamp 1679585382
transform 1 0 141888 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_697
timestamp 1679585382
transform 1 0 142560 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_704
timestamp 1679585382
transform 1 0 143232 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_711
timestamp 1679585382
transform 1 0 143904 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_718
timestamp 1679585382
transform 1 0 144576 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_725
timestamp 1679585382
transform 1 0 145248 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_732
timestamp 1679585382
transform 1 0 145920 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_739
timestamp 1679585382
transform 1 0 146592 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_75_746
timestamp 1679585382
transform 1 0 147264 0 -1 133056
box -48 -56 720 834
use sg13g2_decap_4  FILLER_75_753
timestamp 1679581501
transform 1 0 147936 0 -1 133056
box -48 -56 432 834
use sg13g2_decap_8  FILLER_76_0
timestamp 1679585382
transform 1 0 75648 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_7
timestamp 1679585382
transform 1 0 76320 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_14
timestamp 1679585382
transform 1 0 76992 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_21
timestamp 1679585382
transform 1 0 77664 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_28
timestamp 1679585382
transform 1 0 78336 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_35
timestamp 1679585382
transform 1 0 79008 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_42
timestamp 1679585382
transform 1 0 79680 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_49
timestamp 1679585382
transform 1 0 80352 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_56
timestamp 1679585382
transform 1 0 81024 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_63
timestamp 1679585382
transform 1 0 81696 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_70
timestamp 1679585382
transform 1 0 82368 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_77
timestamp 1679585382
transform 1 0 83040 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_84
timestamp 1679585382
transform 1 0 83712 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_91
timestamp 1679585382
transform 1 0 84384 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_98
timestamp 1679585382
transform 1 0 85056 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_105
timestamp 1679585382
transform 1 0 85728 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_112
timestamp 1679585382
transform 1 0 86400 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_119
timestamp 1679585382
transform 1 0 87072 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_126
timestamp 1679585382
transform 1 0 87744 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_133
timestamp 1679585382
transform 1 0 88416 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_140
timestamp 1679585382
transform 1 0 89088 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_147
timestamp 1679585382
transform 1 0 89760 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_154
timestamp 1679585382
transform 1 0 90432 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_161
timestamp 1679585382
transform 1 0 91104 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_168
timestamp 1679585382
transform 1 0 91776 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_175
timestamp 1679585382
transform 1 0 92448 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_182
timestamp 1679585382
transform 1 0 93120 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_189
timestamp 1679585382
transform 1 0 93792 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_196
timestamp 1679585382
transform 1 0 94464 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_203
timestamp 1679585382
transform 1 0 95136 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_210
timestamp 1679585382
transform 1 0 95808 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_217
timestamp 1679585382
transform 1 0 96480 0 1 133056
box -48 -56 720 834
use sg13g2_decap_4  FILLER_76_224
timestamp 1679581501
transform 1 0 97152 0 1 133056
box -48 -56 432 834
use sg13g2_fill_2  FILLER_76_228
timestamp 1677583704
transform 1 0 97536 0 1 133056
box -48 -56 240 834
use sg13g2_decap_8  FILLER_76_243
timestamp 1679585382
transform 1 0 98976 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_250
timestamp 1679585382
transform 1 0 99648 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_257
timestamp 1679585382
transform 1 0 100320 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_264
timestamp 1679585382
transform 1 0 100992 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_271
timestamp 1679585382
transform 1 0 101664 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_278
timestamp 1679585382
transform 1 0 102336 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_285
timestamp 1679585382
transform 1 0 103008 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_292
timestamp 1679585382
transform 1 0 103680 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_299
timestamp 1679585382
transform 1 0 104352 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_306
timestamp 1679585382
transform 1 0 105024 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_313
timestamp 1679585382
transform 1 0 105696 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_320
timestamp 1679585382
transform 1 0 106368 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_327
timestamp 1679585382
transform 1 0 107040 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_334
timestamp 1679585382
transform 1 0 107712 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_341
timestamp 1679585382
transform 1 0 108384 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_348
timestamp 1679585382
transform 1 0 109056 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_355
timestamp 1679585382
transform 1 0 109728 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_362
timestamp 1679585382
transform 1 0 110400 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_369
timestamp 1679585382
transform 1 0 111072 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_376
timestamp 1679585382
transform 1 0 111744 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_383
timestamp 1679585382
transform 1 0 112416 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_390
timestamp 1679585382
transform 1 0 113088 0 1 133056
box -48 -56 720 834
use sg13g2_fill_2  FILLER_76_397
timestamp 1677583704
transform 1 0 113760 0 1 133056
box -48 -56 240 834
use sg13g2_decap_8  FILLER_76_412
timestamp 1679585382
transform 1 0 115200 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_419
timestamp 1679585382
transform 1 0 115872 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_426
timestamp 1679585382
transform 1 0 116544 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_433
timestamp 1679585382
transform 1 0 117216 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_440
timestamp 1679585382
transform 1 0 117888 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_447
timestamp 1679585382
transform 1 0 118560 0 1 133056
box -48 -56 720 834
use sg13g2_fill_1  FILLER_76_454
timestamp 1677583258
transform 1 0 119232 0 1 133056
box -48 -56 144 834
use sg13g2_decap_8  FILLER_76_482
timestamp 1679585382
transform 1 0 121920 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_489
timestamp 1679585382
transform 1 0 122592 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_496
timestamp 1679585382
transform 1 0 123264 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_503
timestamp 1679585382
transform 1 0 123936 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_510
timestamp 1679585382
transform 1 0 124608 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_517
timestamp 1679585382
transform 1 0 125280 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_524
timestamp 1679585382
transform 1 0 125952 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_531
timestamp 1679585382
transform 1 0 126624 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_538
timestamp 1679585382
transform 1 0 127296 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_545
timestamp 1679585382
transform 1 0 127968 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_552
timestamp 1679585382
transform 1 0 128640 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_559
timestamp 1679585382
transform 1 0 129312 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_566
timestamp 1679585382
transform 1 0 129984 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_573
timestamp 1679585382
transform 1 0 130656 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_580
timestamp 1679585382
transform 1 0 131328 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_587
timestamp 1679585382
transform 1 0 132000 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_594
timestamp 1679585382
transform 1 0 132672 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_601
timestamp 1679585382
transform 1 0 133344 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_608
timestamp 1679585382
transform 1 0 134016 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_615
timestamp 1679585382
transform 1 0 134688 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_622
timestamp 1679585382
transform 1 0 135360 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_629
timestamp 1679585382
transform 1 0 136032 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_636
timestamp 1679585382
transform 1 0 136704 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_643
timestamp 1679585382
transform 1 0 137376 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_650
timestamp 1679585382
transform 1 0 138048 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_657
timestamp 1679585382
transform 1 0 138720 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_664
timestamp 1679585382
transform 1 0 139392 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_671
timestamp 1679585382
transform 1 0 140064 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_678
timestamp 1679585382
transform 1 0 140736 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_685
timestamp 1679585382
transform 1 0 141408 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_692
timestamp 1679585382
transform 1 0 142080 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_699
timestamp 1679585382
transform 1 0 142752 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_706
timestamp 1679585382
transform 1 0 143424 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_713
timestamp 1679585382
transform 1 0 144096 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_720
timestamp 1679585382
transform 1 0 144768 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_727
timestamp 1679585382
transform 1 0 145440 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_734
timestamp 1679585382
transform 1 0 146112 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_741
timestamp 1679585382
transform 1 0 146784 0 1 133056
box -48 -56 720 834
use sg13g2_decap_8  FILLER_76_748
timestamp 1679585382
transform 1 0 147456 0 1 133056
box -48 -56 720 834
use sg13g2_fill_2  FILLER_76_755
timestamp 1677583704
transform 1 0 148128 0 1 133056
box -48 -56 240 834
use sg13g2_decap_8  FILLER_77_0
timestamp 1679585382
transform 1 0 75648 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_7
timestamp 1679585382
transform 1 0 76320 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_14
timestamp 1679585382
transform 1 0 76992 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_21
timestamp 1679585382
transform 1 0 77664 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_28
timestamp 1679585382
transform 1 0 78336 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_35
timestamp 1679585382
transform 1 0 79008 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_42
timestamp 1679585382
transform 1 0 79680 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_49
timestamp 1679585382
transform 1 0 80352 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_56
timestamp 1679585382
transform 1 0 81024 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_63
timestamp 1679585382
transform 1 0 81696 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_70
timestamp 1679585382
transform 1 0 82368 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_77
timestamp 1679585382
transform 1 0 83040 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_84
timestamp 1679585382
transform 1 0 83712 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_91
timestamp 1679585382
transform 1 0 84384 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_98
timestamp 1679585382
transform 1 0 85056 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_105
timestamp 1679585382
transform 1 0 85728 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_112
timestamp 1679585382
transform 1 0 86400 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_119
timestamp 1679585382
transform 1 0 87072 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_126
timestamp 1679585382
transform 1 0 87744 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_133
timestamp 1679585382
transform 1 0 88416 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_140
timestamp 1679585382
transform 1 0 89088 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_147
timestamp 1679585382
transform 1 0 89760 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_154
timestamp 1679585382
transform 1 0 90432 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_161
timestamp 1679585382
transform 1 0 91104 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_168
timestamp 1679585382
transform 1 0 91776 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_175
timestamp 1679585382
transform 1 0 92448 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_182
timestamp 1679585382
transform 1 0 93120 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_189
timestamp 1679585382
transform 1 0 93792 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_196
timestamp 1679585382
transform 1 0 94464 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_203
timestamp 1679585382
transform 1 0 95136 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_210
timestamp 1679585382
transform 1 0 95808 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_217
timestamp 1679585382
transform 1 0 96480 0 -1 134568
box -48 -56 720 834
use sg13g2_fill_2  FILLER_77_224
timestamp 1677583704
transform 1 0 97152 0 -1 134568
box -48 -56 240 834
use sg13g2_decap_8  FILLER_77_253
timestamp 1679585382
transform 1 0 99936 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_260
timestamp 1679585382
transform 1 0 100608 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_267
timestamp 1679585382
transform 1 0 101280 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_274
timestamp 1679585382
transform 1 0 101952 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_281
timestamp 1679585382
transform 1 0 102624 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_288
timestamp 1679585382
transform 1 0 103296 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_295
timestamp 1679585382
transform 1 0 103968 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_302
timestamp 1679585382
transform 1 0 104640 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_309
timestamp 1679585382
transform 1 0 105312 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_316
timestamp 1679585382
transform 1 0 105984 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_323
timestamp 1679585382
transform 1 0 106656 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_330
timestamp 1679585382
transform 1 0 107328 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_337
timestamp 1679585382
transform 1 0 108000 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_344
timestamp 1679585382
transform 1 0 108672 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_351
timestamp 1679585382
transform 1 0 109344 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_358
timestamp 1679585382
transform 1 0 110016 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_365
timestamp 1679585382
transform 1 0 110688 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_372
timestamp 1679585382
transform 1 0 111360 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_379
timestamp 1679585382
transform 1 0 112032 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_386
timestamp 1679585382
transform 1 0 112704 0 -1 134568
box -48 -56 720 834
use sg13g2_fill_1  FILLER_77_393
timestamp 1677583258
transform 1 0 113376 0 -1 134568
box -48 -56 144 834
use sg13g2_decap_8  FILLER_77_421
timestamp 1679585382
transform 1 0 116064 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_428
timestamp 1679585382
transform 1 0 116736 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_435
timestamp 1679585382
transform 1 0 117408 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_442
timestamp 1679585382
transform 1 0 118080 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_449
timestamp 1679585382
transform 1 0 118752 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_4  FILLER_77_456
timestamp 1679581501
transform 1 0 119424 0 -1 134568
box -48 -56 432 834
use sg13g2_decap_8  FILLER_77_464
timestamp 1679585382
transform 1 0 120192 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_471
timestamp 1679585382
transform 1 0 120864 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_478
timestamp 1679585382
transform 1 0 121536 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_485
timestamp 1679585382
transform 1 0 122208 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_492
timestamp 1679585382
transform 1 0 122880 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_499
timestamp 1679585382
transform 1 0 123552 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_506
timestamp 1679585382
transform 1 0 124224 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_513
timestamp 1679585382
transform 1 0 124896 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_520
timestamp 1679585382
transform 1 0 125568 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_527
timestamp 1679585382
transform 1 0 126240 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_534
timestamp 1679585382
transform 1 0 126912 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_541
timestamp 1679585382
transform 1 0 127584 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_548
timestamp 1679585382
transform 1 0 128256 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_555
timestamp 1679585382
transform 1 0 128928 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_562
timestamp 1679585382
transform 1 0 129600 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_569
timestamp 1679585382
transform 1 0 130272 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_576
timestamp 1679585382
transform 1 0 130944 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_583
timestamp 1679585382
transform 1 0 131616 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_590
timestamp 1679585382
transform 1 0 132288 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_597
timestamp 1679585382
transform 1 0 132960 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_604
timestamp 1679585382
transform 1 0 133632 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_611
timestamp 1679585382
transform 1 0 134304 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_618
timestamp 1679585382
transform 1 0 134976 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_625
timestamp 1679585382
transform 1 0 135648 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_632
timestamp 1679585382
transform 1 0 136320 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_639
timestamp 1679585382
transform 1 0 136992 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_646
timestamp 1679585382
transform 1 0 137664 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_653
timestamp 1679585382
transform 1 0 138336 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_660
timestamp 1679585382
transform 1 0 139008 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_667
timestamp 1679585382
transform 1 0 139680 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_674
timestamp 1679585382
transform 1 0 140352 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_681
timestamp 1679585382
transform 1 0 141024 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_688
timestamp 1679585382
transform 1 0 141696 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_695
timestamp 1679585382
transform 1 0 142368 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_702
timestamp 1679585382
transform 1 0 143040 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_709
timestamp 1679585382
transform 1 0 143712 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_716
timestamp 1679585382
transform 1 0 144384 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_723
timestamp 1679585382
transform 1 0 145056 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_730
timestamp 1679585382
transform 1 0 145728 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_737
timestamp 1679585382
transform 1 0 146400 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_77_744
timestamp 1679585382
transform 1 0 147072 0 -1 134568
box -48 -56 720 834
use sg13g2_decap_4  FILLER_77_751
timestamp 1679581501
transform 1 0 147744 0 -1 134568
box -48 -56 432 834
use sg13g2_fill_2  FILLER_77_755
timestamp 1677583704
transform 1 0 148128 0 -1 134568
box -48 -56 240 834
use sg13g2_decap_8  FILLER_78_0
timestamp 1679585382
transform 1 0 75648 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_7
timestamp 1679585382
transform 1 0 76320 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_14
timestamp 1679585382
transform 1 0 76992 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_21
timestamp 1679585382
transform 1 0 77664 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_28
timestamp 1679585382
transform 1 0 78336 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_35
timestamp 1679585382
transform 1 0 79008 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_42
timestamp 1679585382
transform 1 0 79680 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_49
timestamp 1679585382
transform 1 0 80352 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_56
timestamp 1679585382
transform 1 0 81024 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_63
timestamp 1679585382
transform 1 0 81696 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_70
timestamp 1679585382
transform 1 0 82368 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_77
timestamp 1679585382
transform 1 0 83040 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_84
timestamp 1679585382
transform 1 0 83712 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_91
timestamp 1679585382
transform 1 0 84384 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_98
timestamp 1679585382
transform 1 0 85056 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_105
timestamp 1679585382
transform 1 0 85728 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_112
timestamp 1679585382
transform 1 0 86400 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_119
timestamp 1679585382
transform 1 0 87072 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_126
timestamp 1679585382
transform 1 0 87744 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_133
timestamp 1679585382
transform 1 0 88416 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_140
timestamp 1679585382
transform 1 0 89088 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_147
timestamp 1679585382
transform 1 0 89760 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_154
timestamp 1679585382
transform 1 0 90432 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_161
timestamp 1679585382
transform 1 0 91104 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_168
timestamp 1679585382
transform 1 0 91776 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_175
timestamp 1679585382
transform 1 0 92448 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_182
timestamp 1679585382
transform 1 0 93120 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_189
timestamp 1679585382
transform 1 0 93792 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_196
timestamp 1679585382
transform 1 0 94464 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_203
timestamp 1679585382
transform 1 0 95136 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_210
timestamp 1679585382
transform 1 0 95808 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_217
timestamp 1679585382
transform 1 0 96480 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_224
timestamp 1679585382
transform 1 0 97152 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_231
timestamp 1679585382
transform 1 0 97824 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_238
timestamp 1679585382
transform 1 0 98496 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_245
timestamp 1679585382
transform 1 0 99168 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_252
timestamp 1679585382
transform 1 0 99840 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_259
timestamp 1679585382
transform 1 0 100512 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_266
timestamp 1679585382
transform 1 0 101184 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_273
timestamp 1679585382
transform 1 0 101856 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_280
timestamp 1679585382
transform 1 0 102528 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_287
timestamp 1679585382
transform 1 0 103200 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_294
timestamp 1679585382
transform 1 0 103872 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_301
timestamp 1679585382
transform 1 0 104544 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_308
timestamp 1679585382
transform 1 0 105216 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_315
timestamp 1679585382
transform 1 0 105888 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_322
timestamp 1679585382
transform 1 0 106560 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_329
timestamp 1679585382
transform 1 0 107232 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_336
timestamp 1679585382
transform 1 0 107904 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_343
timestamp 1679585382
transform 1 0 108576 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_350
timestamp 1679585382
transform 1 0 109248 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_357
timestamp 1679585382
transform 1 0 109920 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_364
timestamp 1679585382
transform 1 0 110592 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_371
timestamp 1679585382
transform 1 0 111264 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_378
timestamp 1679585382
transform 1 0 111936 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_385
timestamp 1679585382
transform 1 0 112608 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_392
timestamp 1679585382
transform 1 0 113280 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_399
timestamp 1679585382
transform 1 0 113952 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_406
timestamp 1679585382
transform 1 0 114624 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_413
timestamp 1679585382
transform 1 0 115296 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_420
timestamp 1679585382
transform 1 0 115968 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_427
timestamp 1679585382
transform 1 0 116640 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_434
timestamp 1679585382
transform 1 0 117312 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_441
timestamp 1679585382
transform 1 0 117984 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_448
timestamp 1679585382
transform 1 0 118656 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_455
timestamp 1679585382
transform 1 0 119328 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_462
timestamp 1679585382
transform 1 0 120000 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_469
timestamp 1679585382
transform 1 0 120672 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_476
timestamp 1679585382
transform 1 0 121344 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_483
timestamp 1679585382
transform 1 0 122016 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_490
timestamp 1679585382
transform 1 0 122688 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_497
timestamp 1679585382
transform 1 0 123360 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_504
timestamp 1679585382
transform 1 0 124032 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_511
timestamp 1679585382
transform 1 0 124704 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_518
timestamp 1679585382
transform 1 0 125376 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_525
timestamp 1679585382
transform 1 0 126048 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_532
timestamp 1679585382
transform 1 0 126720 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_539
timestamp 1679585382
transform 1 0 127392 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_546
timestamp 1679585382
transform 1 0 128064 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_553
timestamp 1679585382
transform 1 0 128736 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_560
timestamp 1679585382
transform 1 0 129408 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_567
timestamp 1679585382
transform 1 0 130080 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_574
timestamp 1679585382
transform 1 0 130752 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_581
timestamp 1679585382
transform 1 0 131424 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_588
timestamp 1679585382
transform 1 0 132096 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_595
timestamp 1679585382
transform 1 0 132768 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_602
timestamp 1679585382
transform 1 0 133440 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_609
timestamp 1679585382
transform 1 0 134112 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_616
timestamp 1679585382
transform 1 0 134784 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_623
timestamp 1679585382
transform 1 0 135456 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_630
timestamp 1679585382
transform 1 0 136128 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_637
timestamp 1679585382
transform 1 0 136800 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_644
timestamp 1679585382
transform 1 0 137472 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_651
timestamp 1679585382
transform 1 0 138144 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_658
timestamp 1679585382
transform 1 0 138816 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_665
timestamp 1679585382
transform 1 0 139488 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_672
timestamp 1679585382
transform 1 0 140160 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_679
timestamp 1679585382
transform 1 0 140832 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_686
timestamp 1679585382
transform 1 0 141504 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_693
timestamp 1679585382
transform 1 0 142176 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_700
timestamp 1679585382
transform 1 0 142848 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_707
timestamp 1679585382
transform 1 0 143520 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_714
timestamp 1679585382
transform 1 0 144192 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_721
timestamp 1679585382
transform 1 0 144864 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_728
timestamp 1679585382
transform 1 0 145536 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_735
timestamp 1679585382
transform 1 0 146208 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_742
timestamp 1679585382
transform 1 0 146880 0 1 134568
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_749
timestamp 1679585382
transform 1 0 147552 0 1 134568
box -48 -56 720 834
use sg13g2_fill_1  FILLER_78_756
timestamp 1677583258
transform 1 0 148224 0 1 134568
box -48 -56 144 834
use sg13g2_decap_8  FILLER_79_0
timestamp 1679585382
transform 1 0 75648 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_7
timestamp 1679585382
transform 1 0 76320 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_14
timestamp 1679585382
transform 1 0 76992 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_21
timestamp 1679585382
transform 1 0 77664 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_28
timestamp 1679585382
transform 1 0 78336 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_35
timestamp 1679585382
transform 1 0 79008 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_42
timestamp 1679585382
transform 1 0 79680 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_49
timestamp 1679585382
transform 1 0 80352 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_56
timestamp 1679585382
transform 1 0 81024 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_63
timestamp 1679585382
transform 1 0 81696 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_70
timestamp 1679585382
transform 1 0 82368 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_77
timestamp 1679585382
transform 1 0 83040 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_84
timestamp 1679585382
transform 1 0 83712 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_91
timestamp 1679585382
transform 1 0 84384 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_98
timestamp 1679585382
transform 1 0 85056 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_105
timestamp 1679585382
transform 1 0 85728 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_112
timestamp 1679585382
transform 1 0 86400 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_119
timestamp 1679585382
transform 1 0 87072 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_126
timestamp 1679585382
transform 1 0 87744 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_133
timestamp 1679585382
transform 1 0 88416 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_140
timestamp 1679585382
transform 1 0 89088 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_147
timestamp 1679585382
transform 1 0 89760 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_154
timestamp 1679585382
transform 1 0 90432 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_161
timestamp 1679585382
transform 1 0 91104 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_168
timestamp 1679585382
transform 1 0 91776 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_175
timestamp 1679585382
transform 1 0 92448 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_182
timestamp 1679585382
transform 1 0 93120 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_189
timestamp 1679585382
transform 1 0 93792 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_196
timestamp 1679585382
transform 1 0 94464 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_203
timestamp 1679585382
transform 1 0 95136 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_210
timestamp 1679585382
transform 1 0 95808 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_217
timestamp 1679585382
transform 1 0 96480 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_224
timestamp 1679585382
transform 1 0 97152 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_231
timestamp 1679585382
transform 1 0 97824 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_238
timestamp 1679585382
transform 1 0 98496 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_245
timestamp 1679585382
transform 1 0 99168 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_252
timestamp 1679585382
transform 1 0 99840 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_259
timestamp 1679585382
transform 1 0 100512 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_266
timestamp 1679585382
transform 1 0 101184 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_273
timestamp 1679585382
transform 1 0 101856 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_280
timestamp 1679585382
transform 1 0 102528 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_287
timestamp 1679585382
transform 1 0 103200 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_294
timestamp 1679585382
transform 1 0 103872 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_301
timestamp 1679585382
transform 1 0 104544 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_308
timestamp 1679585382
transform 1 0 105216 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_315
timestamp 1679585382
transform 1 0 105888 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_322
timestamp 1679585382
transform 1 0 106560 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_329
timestamp 1679585382
transform 1 0 107232 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_336
timestamp 1679585382
transform 1 0 107904 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_343
timestamp 1679585382
transform 1 0 108576 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_350
timestamp 1679585382
transform 1 0 109248 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_357
timestamp 1679585382
transform 1 0 109920 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_364
timestamp 1679585382
transform 1 0 110592 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_371
timestamp 1679585382
transform 1 0 111264 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_378
timestamp 1679585382
transform 1 0 111936 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_385
timestamp 1679585382
transform 1 0 112608 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_392
timestamp 1679585382
transform 1 0 113280 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_399
timestamp 1679585382
transform 1 0 113952 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_406
timestamp 1679585382
transform 1 0 114624 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_413
timestamp 1679585382
transform 1 0 115296 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_420
timestamp 1679585382
transform 1 0 115968 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_427
timestamp 1679585382
transform 1 0 116640 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_434
timestamp 1679585382
transform 1 0 117312 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_441
timestamp 1679585382
transform 1 0 117984 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_448
timestamp 1679585382
transform 1 0 118656 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_455
timestamp 1679585382
transform 1 0 119328 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_462
timestamp 1679585382
transform 1 0 120000 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_469
timestamp 1679585382
transform 1 0 120672 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_476
timestamp 1679585382
transform 1 0 121344 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_483
timestamp 1679585382
transform 1 0 122016 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_490
timestamp 1679585382
transform 1 0 122688 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_497
timestamp 1679585382
transform 1 0 123360 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_504
timestamp 1679585382
transform 1 0 124032 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_511
timestamp 1679585382
transform 1 0 124704 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_518
timestamp 1679585382
transform 1 0 125376 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_525
timestamp 1679585382
transform 1 0 126048 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_532
timestamp 1679585382
transform 1 0 126720 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_539
timestamp 1679585382
transform 1 0 127392 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_546
timestamp 1679585382
transform 1 0 128064 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_553
timestamp 1679585382
transform 1 0 128736 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_560
timestamp 1679585382
transform 1 0 129408 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_567
timestamp 1679585382
transform 1 0 130080 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_574
timestamp 1679585382
transform 1 0 130752 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_581
timestamp 1679585382
transform 1 0 131424 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_588
timestamp 1679585382
transform 1 0 132096 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_595
timestamp 1679585382
transform 1 0 132768 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_602
timestamp 1679585382
transform 1 0 133440 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_609
timestamp 1679585382
transform 1 0 134112 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_616
timestamp 1679585382
transform 1 0 134784 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_623
timestamp 1679585382
transform 1 0 135456 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_630
timestamp 1679585382
transform 1 0 136128 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_637
timestamp 1679585382
transform 1 0 136800 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_644
timestamp 1679585382
transform 1 0 137472 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_651
timestamp 1679585382
transform 1 0 138144 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_658
timestamp 1679585382
transform 1 0 138816 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_665
timestamp 1679585382
transform 1 0 139488 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_672
timestamp 1679585382
transform 1 0 140160 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_679
timestamp 1679585382
transform 1 0 140832 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_686
timestamp 1679585382
transform 1 0 141504 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_693
timestamp 1679585382
transform 1 0 142176 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_700
timestamp 1679585382
transform 1 0 142848 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_707
timestamp 1679585382
transform 1 0 143520 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_714
timestamp 1679585382
transform 1 0 144192 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_721
timestamp 1679585382
transform 1 0 144864 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_728
timestamp 1679585382
transform 1 0 145536 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_735
timestamp 1679585382
transform 1 0 146208 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_742
timestamp 1679585382
transform 1 0 146880 0 -1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_79_749
timestamp 1679585382
transform 1 0 147552 0 -1 136080
box -48 -56 720 834
use sg13g2_fill_1  FILLER_79_756
timestamp 1677583258
transform 1 0 148224 0 -1 136080
box -48 -56 144 834
use sg13g2_decap_8  FILLER_80_0
timestamp 1679585382
transform 1 0 75648 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_7
timestamp 1679585382
transform 1 0 76320 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_14
timestamp 1679585382
transform 1 0 76992 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_21
timestamp 1679585382
transform 1 0 77664 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_28
timestamp 1679585382
transform 1 0 78336 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_35
timestamp 1679585382
transform 1 0 79008 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_42
timestamp 1679585382
transform 1 0 79680 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_49
timestamp 1679585382
transform 1 0 80352 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_56
timestamp 1679585382
transform 1 0 81024 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_63
timestamp 1679585382
transform 1 0 81696 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_70
timestamp 1679585382
transform 1 0 82368 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_77
timestamp 1679585382
transform 1 0 83040 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_84
timestamp 1679585382
transform 1 0 83712 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_91
timestamp 1679585382
transform 1 0 84384 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_98
timestamp 1679585382
transform 1 0 85056 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_105
timestamp 1679585382
transform 1 0 85728 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_112
timestamp 1679585382
transform 1 0 86400 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_119
timestamp 1679585382
transform 1 0 87072 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_126
timestamp 1679585382
transform 1 0 87744 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_133
timestamp 1679585382
transform 1 0 88416 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_140
timestamp 1679585382
transform 1 0 89088 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_147
timestamp 1679585382
transform 1 0 89760 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_154
timestamp 1679585382
transform 1 0 90432 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_161
timestamp 1679585382
transform 1 0 91104 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_168
timestamp 1679585382
transform 1 0 91776 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_175
timestamp 1679585382
transform 1 0 92448 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_182
timestamp 1679585382
transform 1 0 93120 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_189
timestamp 1679585382
transform 1 0 93792 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_196
timestamp 1679585382
transform 1 0 94464 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_203
timestamp 1679585382
transform 1 0 95136 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_210
timestamp 1679585382
transform 1 0 95808 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_217
timestamp 1679585382
transform 1 0 96480 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_224
timestamp 1679585382
transform 1 0 97152 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_231
timestamp 1679585382
transform 1 0 97824 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_238
timestamp 1679585382
transform 1 0 98496 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_245
timestamp 1679585382
transform 1 0 99168 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_252
timestamp 1679585382
transform 1 0 99840 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_259
timestamp 1679585382
transform 1 0 100512 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_266
timestamp 1679585382
transform 1 0 101184 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_273
timestamp 1679585382
transform 1 0 101856 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_280
timestamp 1679585382
transform 1 0 102528 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_287
timestamp 1679585382
transform 1 0 103200 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_294
timestamp 1679585382
transform 1 0 103872 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_301
timestamp 1679585382
transform 1 0 104544 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_308
timestamp 1679585382
transform 1 0 105216 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_315
timestamp 1679585382
transform 1 0 105888 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_322
timestamp 1679585382
transform 1 0 106560 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_329
timestamp 1679585382
transform 1 0 107232 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_336
timestamp 1679585382
transform 1 0 107904 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_343
timestamp 1679585382
transform 1 0 108576 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_350
timestamp 1679585382
transform 1 0 109248 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_357
timestamp 1679585382
transform 1 0 109920 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_364
timestamp 1679585382
transform 1 0 110592 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_371
timestamp 1679585382
transform 1 0 111264 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_378
timestamp 1679585382
transform 1 0 111936 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_385
timestamp 1679585382
transform 1 0 112608 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_392
timestamp 1679585382
transform 1 0 113280 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_399
timestamp 1679585382
transform 1 0 113952 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_406
timestamp 1679585382
transform 1 0 114624 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_413
timestamp 1679585382
transform 1 0 115296 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_420
timestamp 1679585382
transform 1 0 115968 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_427
timestamp 1679585382
transform 1 0 116640 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_434
timestamp 1679585382
transform 1 0 117312 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_441
timestamp 1679585382
transform 1 0 117984 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_448
timestamp 1679585382
transform 1 0 118656 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_455
timestamp 1679585382
transform 1 0 119328 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_462
timestamp 1679585382
transform 1 0 120000 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_469
timestamp 1679585382
transform 1 0 120672 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_476
timestamp 1679585382
transform 1 0 121344 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_483
timestamp 1679585382
transform 1 0 122016 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_490
timestamp 1679585382
transform 1 0 122688 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_497
timestamp 1679585382
transform 1 0 123360 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_504
timestamp 1679585382
transform 1 0 124032 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_511
timestamp 1679585382
transform 1 0 124704 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_518
timestamp 1679585382
transform 1 0 125376 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_525
timestamp 1679585382
transform 1 0 126048 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_532
timestamp 1679585382
transform 1 0 126720 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_539
timestamp 1679585382
transform 1 0 127392 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_546
timestamp 1679585382
transform 1 0 128064 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_553
timestamp 1679585382
transform 1 0 128736 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_560
timestamp 1679585382
transform 1 0 129408 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_567
timestamp 1679585382
transform 1 0 130080 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_574
timestamp 1679585382
transform 1 0 130752 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_581
timestamp 1679585382
transform 1 0 131424 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_588
timestamp 1679585382
transform 1 0 132096 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_595
timestamp 1679585382
transform 1 0 132768 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_602
timestamp 1679585382
transform 1 0 133440 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_609
timestamp 1679585382
transform 1 0 134112 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_616
timestamp 1679585382
transform 1 0 134784 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_623
timestamp 1679585382
transform 1 0 135456 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_630
timestamp 1679585382
transform 1 0 136128 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_637
timestamp 1679585382
transform 1 0 136800 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_644
timestamp 1679585382
transform 1 0 137472 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_651
timestamp 1679585382
transform 1 0 138144 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_658
timestamp 1679585382
transform 1 0 138816 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_665
timestamp 1679585382
transform 1 0 139488 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_672
timestamp 1679585382
transform 1 0 140160 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_679
timestamp 1679585382
transform 1 0 140832 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_686
timestamp 1679585382
transform 1 0 141504 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_693
timestamp 1679585382
transform 1 0 142176 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_700
timestamp 1679585382
transform 1 0 142848 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_707
timestamp 1679585382
transform 1 0 143520 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_714
timestamp 1679585382
transform 1 0 144192 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_721
timestamp 1679585382
transform 1 0 144864 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_728
timestamp 1679585382
transform 1 0 145536 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_735
timestamp 1679585382
transform 1 0 146208 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_742
timestamp 1679585382
transform 1 0 146880 0 1 136080
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_749
timestamp 1679585382
transform 1 0 147552 0 1 136080
box -48 -56 720 834
use sg13g2_fill_1  FILLER_80_756
timestamp 1677583258
transform 1 0 148224 0 1 136080
box -48 -56 144 834
use sg13g2_decap_8  FILLER_81_0
timestamp 1679585382
transform 1 0 75648 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_7
timestamp 1679585382
transform 1 0 76320 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_14
timestamp 1679585382
transform 1 0 76992 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_21
timestamp 1679585382
transform 1 0 77664 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_28
timestamp 1679585382
transform 1 0 78336 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_35
timestamp 1679585382
transform 1 0 79008 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_42
timestamp 1679585382
transform 1 0 79680 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_49
timestamp 1679585382
transform 1 0 80352 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_56
timestamp 1679585382
transform 1 0 81024 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_63
timestamp 1679585382
transform 1 0 81696 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_70
timestamp 1679585382
transform 1 0 82368 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_77
timestamp 1679585382
transform 1 0 83040 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_84
timestamp 1679585382
transform 1 0 83712 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_91
timestamp 1679585382
transform 1 0 84384 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_98
timestamp 1679585382
transform 1 0 85056 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_105
timestamp 1679585382
transform 1 0 85728 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_112
timestamp 1679585382
transform 1 0 86400 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_119
timestamp 1679585382
transform 1 0 87072 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_126
timestamp 1679585382
transform 1 0 87744 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_133
timestamp 1679585382
transform 1 0 88416 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_140
timestamp 1679585382
transform 1 0 89088 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_147
timestamp 1679585382
transform 1 0 89760 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_154
timestamp 1679585382
transform 1 0 90432 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_161
timestamp 1679585382
transform 1 0 91104 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_168
timestamp 1679585382
transform 1 0 91776 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_175
timestamp 1679585382
transform 1 0 92448 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_182
timestamp 1679585382
transform 1 0 93120 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_189
timestamp 1679585382
transform 1 0 93792 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_196
timestamp 1679585382
transform 1 0 94464 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_203
timestamp 1679585382
transform 1 0 95136 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_210
timestamp 1679585382
transform 1 0 95808 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_217
timestamp 1679585382
transform 1 0 96480 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_224
timestamp 1679585382
transform 1 0 97152 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_231
timestamp 1679585382
transform 1 0 97824 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_238
timestamp 1679585382
transform 1 0 98496 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_245
timestamp 1679585382
transform 1 0 99168 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_252
timestamp 1679585382
transform 1 0 99840 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_259
timestamp 1679585382
transform 1 0 100512 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_266
timestamp 1679585382
transform 1 0 101184 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_273
timestamp 1679585382
transform 1 0 101856 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_280
timestamp 1679585382
transform 1 0 102528 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_287
timestamp 1679585382
transform 1 0 103200 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_294
timestamp 1679585382
transform 1 0 103872 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_301
timestamp 1679585382
transform 1 0 104544 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_308
timestamp 1679585382
transform 1 0 105216 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_315
timestamp 1679585382
transform 1 0 105888 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_322
timestamp 1679585382
transform 1 0 106560 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_329
timestamp 1679585382
transform 1 0 107232 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_336
timestamp 1679585382
transform 1 0 107904 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_343
timestamp 1679585382
transform 1 0 108576 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_350
timestamp 1679585382
transform 1 0 109248 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_357
timestamp 1679585382
transform 1 0 109920 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_364
timestamp 1679585382
transform 1 0 110592 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_371
timestamp 1679585382
transform 1 0 111264 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_378
timestamp 1679585382
transform 1 0 111936 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_385
timestamp 1679585382
transform 1 0 112608 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_392
timestamp 1679585382
transform 1 0 113280 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_399
timestamp 1679585382
transform 1 0 113952 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_406
timestamp 1679585382
transform 1 0 114624 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_413
timestamp 1679585382
transform 1 0 115296 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_420
timestamp 1679585382
transform 1 0 115968 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_427
timestamp 1679585382
transform 1 0 116640 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_434
timestamp 1679585382
transform 1 0 117312 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_441
timestamp 1679585382
transform 1 0 117984 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_448
timestamp 1679585382
transform 1 0 118656 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_455
timestamp 1679585382
transform 1 0 119328 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_462
timestamp 1679585382
transform 1 0 120000 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_469
timestamp 1679585382
transform 1 0 120672 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_476
timestamp 1679585382
transform 1 0 121344 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_483
timestamp 1679585382
transform 1 0 122016 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_490
timestamp 1679585382
transform 1 0 122688 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_497
timestamp 1679585382
transform 1 0 123360 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_504
timestamp 1679585382
transform 1 0 124032 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_511
timestamp 1679585382
transform 1 0 124704 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_518
timestamp 1679585382
transform 1 0 125376 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_525
timestamp 1679585382
transform 1 0 126048 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_532
timestamp 1679585382
transform 1 0 126720 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_539
timestamp 1679585382
transform 1 0 127392 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_546
timestamp 1679585382
transform 1 0 128064 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_553
timestamp 1679585382
transform 1 0 128736 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_560
timestamp 1679585382
transform 1 0 129408 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_567
timestamp 1679585382
transform 1 0 130080 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_574
timestamp 1679585382
transform 1 0 130752 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_581
timestamp 1679585382
transform 1 0 131424 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_588
timestamp 1679585382
transform 1 0 132096 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_595
timestamp 1679585382
transform 1 0 132768 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_602
timestamp 1679585382
transform 1 0 133440 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_609
timestamp 1679585382
transform 1 0 134112 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_616
timestamp 1679585382
transform 1 0 134784 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_623
timestamp 1679585382
transform 1 0 135456 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_630
timestamp 1679585382
transform 1 0 136128 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_637
timestamp 1679585382
transform 1 0 136800 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_644
timestamp 1679585382
transform 1 0 137472 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_651
timestamp 1679585382
transform 1 0 138144 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_658
timestamp 1679585382
transform 1 0 138816 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_665
timestamp 1679585382
transform 1 0 139488 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_672
timestamp 1679585382
transform 1 0 140160 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_679
timestamp 1679585382
transform 1 0 140832 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_686
timestamp 1679585382
transform 1 0 141504 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_693
timestamp 1679585382
transform 1 0 142176 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_700
timestamp 1679585382
transform 1 0 142848 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_707
timestamp 1679585382
transform 1 0 143520 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_714
timestamp 1679585382
transform 1 0 144192 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_721
timestamp 1679585382
transform 1 0 144864 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_728
timestamp 1679585382
transform 1 0 145536 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_735
timestamp 1679585382
transform 1 0 146208 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_742
timestamp 1679585382
transform 1 0 146880 0 -1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_81_749
timestamp 1679585382
transform 1 0 147552 0 -1 137592
box -48 -56 720 834
use sg13g2_fill_1  FILLER_81_756
timestamp 1677583258
transform 1 0 148224 0 -1 137592
box -48 -56 144 834
use sg13g2_decap_8  FILLER_82_0
timestamp 1679585382
transform 1 0 75648 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_7
timestamp 1679585382
transform 1 0 76320 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_14
timestamp 1679585382
transform 1 0 76992 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_21
timestamp 1679585382
transform 1 0 77664 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_28
timestamp 1679585382
transform 1 0 78336 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_35
timestamp 1679585382
transform 1 0 79008 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_42
timestamp 1679585382
transform 1 0 79680 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_49
timestamp 1679585382
transform 1 0 80352 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_56
timestamp 1679585382
transform 1 0 81024 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_63
timestamp 1679585382
transform 1 0 81696 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_70
timestamp 1679585382
transform 1 0 82368 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_77
timestamp 1679585382
transform 1 0 83040 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_84
timestamp 1679585382
transform 1 0 83712 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_91
timestamp 1679585382
transform 1 0 84384 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_98
timestamp 1679585382
transform 1 0 85056 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_105
timestamp 1679585382
transform 1 0 85728 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_112
timestamp 1679585382
transform 1 0 86400 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_119
timestamp 1679585382
transform 1 0 87072 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_126
timestamp 1679585382
transform 1 0 87744 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_133
timestamp 1679585382
transform 1 0 88416 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_140
timestamp 1679585382
transform 1 0 89088 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_147
timestamp 1679585382
transform 1 0 89760 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_154
timestamp 1679585382
transform 1 0 90432 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_161
timestamp 1679585382
transform 1 0 91104 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_168
timestamp 1679585382
transform 1 0 91776 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_175
timestamp 1679585382
transform 1 0 92448 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_182
timestamp 1679585382
transform 1 0 93120 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_189
timestamp 1679585382
transform 1 0 93792 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_196
timestamp 1679585382
transform 1 0 94464 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_203
timestamp 1679585382
transform 1 0 95136 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_210
timestamp 1679585382
transform 1 0 95808 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_217
timestamp 1679585382
transform 1 0 96480 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_224
timestamp 1679585382
transform 1 0 97152 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_231
timestamp 1679585382
transform 1 0 97824 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_238
timestamp 1679585382
transform 1 0 98496 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_245
timestamp 1679585382
transform 1 0 99168 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_252
timestamp 1679585382
transform 1 0 99840 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_259
timestamp 1679585382
transform 1 0 100512 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_266
timestamp 1679585382
transform 1 0 101184 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_273
timestamp 1679585382
transform 1 0 101856 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_280
timestamp 1679585382
transform 1 0 102528 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_287
timestamp 1679585382
transform 1 0 103200 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_294
timestamp 1679585382
transform 1 0 103872 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_301
timestamp 1679585382
transform 1 0 104544 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_308
timestamp 1679585382
transform 1 0 105216 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_315
timestamp 1679585382
transform 1 0 105888 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_322
timestamp 1679585382
transform 1 0 106560 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_329
timestamp 1679585382
transform 1 0 107232 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_336
timestamp 1679585382
transform 1 0 107904 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_343
timestamp 1679585382
transform 1 0 108576 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_350
timestamp 1679585382
transform 1 0 109248 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_357
timestamp 1679585382
transform 1 0 109920 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_364
timestamp 1679585382
transform 1 0 110592 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_371
timestamp 1679585382
transform 1 0 111264 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_378
timestamp 1679585382
transform 1 0 111936 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_385
timestamp 1679585382
transform 1 0 112608 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_392
timestamp 1679585382
transform 1 0 113280 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_399
timestamp 1679585382
transform 1 0 113952 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_406
timestamp 1679585382
transform 1 0 114624 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_413
timestamp 1679585382
transform 1 0 115296 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_420
timestamp 1679585382
transform 1 0 115968 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_427
timestamp 1679585382
transform 1 0 116640 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_434
timestamp 1679585382
transform 1 0 117312 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_441
timestamp 1679585382
transform 1 0 117984 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_448
timestamp 1679585382
transform 1 0 118656 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_455
timestamp 1679585382
transform 1 0 119328 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_462
timestamp 1679585382
transform 1 0 120000 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_469
timestamp 1679585382
transform 1 0 120672 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_476
timestamp 1679585382
transform 1 0 121344 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_483
timestamp 1679585382
transform 1 0 122016 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_490
timestamp 1679585382
transform 1 0 122688 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_497
timestamp 1679585382
transform 1 0 123360 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_504
timestamp 1679585382
transform 1 0 124032 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_511
timestamp 1679585382
transform 1 0 124704 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_518
timestamp 1679585382
transform 1 0 125376 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_525
timestamp 1679585382
transform 1 0 126048 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_532
timestamp 1679585382
transform 1 0 126720 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_539
timestamp 1679585382
transform 1 0 127392 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_546
timestamp 1679585382
transform 1 0 128064 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_553
timestamp 1679585382
transform 1 0 128736 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_560
timestamp 1679585382
transform 1 0 129408 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_567
timestamp 1679585382
transform 1 0 130080 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_574
timestamp 1679585382
transform 1 0 130752 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_581
timestamp 1679585382
transform 1 0 131424 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_588
timestamp 1679585382
transform 1 0 132096 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_595
timestamp 1679585382
transform 1 0 132768 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_602
timestamp 1679585382
transform 1 0 133440 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_609
timestamp 1679585382
transform 1 0 134112 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_616
timestamp 1679585382
transform 1 0 134784 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_623
timestamp 1679585382
transform 1 0 135456 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_630
timestamp 1679585382
transform 1 0 136128 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_637
timestamp 1679585382
transform 1 0 136800 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_644
timestamp 1679585382
transform 1 0 137472 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_651
timestamp 1679585382
transform 1 0 138144 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_658
timestamp 1679585382
transform 1 0 138816 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_665
timestamp 1679585382
transform 1 0 139488 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_672
timestamp 1679585382
transform 1 0 140160 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_679
timestamp 1679585382
transform 1 0 140832 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_686
timestamp 1679585382
transform 1 0 141504 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_693
timestamp 1679585382
transform 1 0 142176 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_700
timestamp 1679585382
transform 1 0 142848 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_707
timestamp 1679585382
transform 1 0 143520 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_714
timestamp 1679585382
transform 1 0 144192 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_721
timestamp 1679585382
transform 1 0 144864 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_728
timestamp 1679585382
transform 1 0 145536 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_735
timestamp 1679585382
transform 1 0 146208 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_742
timestamp 1679585382
transform 1 0 146880 0 1 137592
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_749
timestamp 1679585382
transform 1 0 147552 0 1 137592
box -48 -56 720 834
use sg13g2_fill_1  FILLER_82_756
timestamp 1677583258
transform 1 0 148224 0 1 137592
box -48 -56 144 834
use sg13g2_decap_8  FILLER_83_0
timestamp 1679585382
transform 1 0 75648 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_7
timestamp 1679585382
transform 1 0 76320 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_14
timestamp 1679585382
transform 1 0 76992 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_21
timestamp 1679585382
transform 1 0 77664 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_28
timestamp 1679585382
transform 1 0 78336 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_35
timestamp 1679585382
transform 1 0 79008 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_42
timestamp 1679585382
transform 1 0 79680 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_49
timestamp 1679585382
transform 1 0 80352 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_56
timestamp 1679585382
transform 1 0 81024 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_63
timestamp 1679585382
transform 1 0 81696 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_70
timestamp 1679585382
transform 1 0 82368 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_77
timestamp 1679585382
transform 1 0 83040 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_84
timestamp 1679585382
transform 1 0 83712 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_91
timestamp 1679585382
transform 1 0 84384 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_98
timestamp 1679585382
transform 1 0 85056 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_105
timestamp 1679585382
transform 1 0 85728 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_112
timestamp 1679585382
transform 1 0 86400 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_119
timestamp 1679585382
transform 1 0 87072 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_126
timestamp 1679585382
transform 1 0 87744 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_133
timestamp 1679585382
transform 1 0 88416 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_140
timestamp 1679585382
transform 1 0 89088 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_147
timestamp 1679585382
transform 1 0 89760 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_154
timestamp 1679585382
transform 1 0 90432 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_161
timestamp 1679585382
transform 1 0 91104 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_168
timestamp 1679585382
transform 1 0 91776 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_175
timestamp 1679585382
transform 1 0 92448 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_182
timestamp 1679585382
transform 1 0 93120 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_189
timestamp 1679585382
transform 1 0 93792 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_196
timestamp 1679585382
transform 1 0 94464 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_203
timestamp 1679585382
transform 1 0 95136 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_210
timestamp 1679585382
transform 1 0 95808 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_217
timestamp 1679585382
transform 1 0 96480 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_224
timestamp 1679585382
transform 1 0 97152 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_231
timestamp 1679585382
transform 1 0 97824 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_238
timestamp 1679585382
transform 1 0 98496 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_245
timestamp 1679585382
transform 1 0 99168 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_252
timestamp 1679585382
transform 1 0 99840 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_259
timestamp 1679585382
transform 1 0 100512 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_266
timestamp 1679585382
transform 1 0 101184 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_273
timestamp 1679585382
transform 1 0 101856 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_280
timestamp 1679585382
transform 1 0 102528 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_287
timestamp 1679585382
transform 1 0 103200 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_294
timestamp 1679585382
transform 1 0 103872 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_301
timestamp 1679585382
transform 1 0 104544 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_308
timestamp 1679585382
transform 1 0 105216 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_315
timestamp 1679585382
transform 1 0 105888 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_322
timestamp 1679585382
transform 1 0 106560 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_329
timestamp 1679585382
transform 1 0 107232 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_336
timestamp 1679585382
transform 1 0 107904 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_343
timestamp 1679585382
transform 1 0 108576 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_350
timestamp 1679585382
transform 1 0 109248 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_357
timestamp 1679585382
transform 1 0 109920 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_364
timestamp 1679585382
transform 1 0 110592 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_371
timestamp 1679585382
transform 1 0 111264 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_378
timestamp 1679585382
transform 1 0 111936 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_385
timestamp 1679585382
transform 1 0 112608 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_392
timestamp 1679585382
transform 1 0 113280 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_399
timestamp 1679585382
transform 1 0 113952 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_406
timestamp 1679585382
transform 1 0 114624 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_413
timestamp 1679585382
transform 1 0 115296 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_420
timestamp 1679585382
transform 1 0 115968 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_427
timestamp 1679585382
transform 1 0 116640 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_434
timestamp 1679585382
transform 1 0 117312 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_441
timestamp 1679585382
transform 1 0 117984 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_448
timestamp 1679585382
transform 1 0 118656 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_455
timestamp 1679585382
transform 1 0 119328 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_462
timestamp 1679585382
transform 1 0 120000 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_469
timestamp 1679585382
transform 1 0 120672 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_476
timestamp 1679585382
transform 1 0 121344 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_483
timestamp 1679585382
transform 1 0 122016 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_490
timestamp 1679585382
transform 1 0 122688 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_497
timestamp 1679585382
transform 1 0 123360 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_504
timestamp 1679585382
transform 1 0 124032 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_511
timestamp 1679585382
transform 1 0 124704 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_518
timestamp 1679585382
transform 1 0 125376 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_525
timestamp 1679585382
transform 1 0 126048 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_532
timestamp 1679585382
transform 1 0 126720 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_539
timestamp 1679585382
transform 1 0 127392 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_546
timestamp 1679585382
transform 1 0 128064 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_553
timestamp 1679585382
transform 1 0 128736 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_560
timestamp 1679585382
transform 1 0 129408 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_567
timestamp 1679585382
transform 1 0 130080 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_574
timestamp 1679585382
transform 1 0 130752 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_581
timestamp 1679585382
transform 1 0 131424 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_588
timestamp 1679585382
transform 1 0 132096 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_595
timestamp 1679585382
transform 1 0 132768 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_602
timestamp 1679585382
transform 1 0 133440 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_609
timestamp 1679585382
transform 1 0 134112 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_616
timestamp 1679585382
transform 1 0 134784 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_623
timestamp 1679585382
transform 1 0 135456 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_630
timestamp 1679585382
transform 1 0 136128 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_637
timestamp 1679585382
transform 1 0 136800 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_644
timestamp 1679585382
transform 1 0 137472 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_651
timestamp 1679585382
transform 1 0 138144 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_658
timestamp 1679585382
transform 1 0 138816 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_665
timestamp 1679585382
transform 1 0 139488 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_672
timestamp 1679585382
transform 1 0 140160 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_679
timestamp 1679585382
transform 1 0 140832 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_686
timestamp 1679585382
transform 1 0 141504 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_693
timestamp 1679585382
transform 1 0 142176 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_700
timestamp 1679585382
transform 1 0 142848 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_707
timestamp 1679585382
transform 1 0 143520 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_714
timestamp 1679585382
transform 1 0 144192 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_721
timestamp 1679585382
transform 1 0 144864 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_728
timestamp 1679585382
transform 1 0 145536 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_735
timestamp 1679585382
transform 1 0 146208 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_742
timestamp 1679585382
transform 1 0 146880 0 -1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_83_749
timestamp 1679585382
transform 1 0 147552 0 -1 139104
box -48 -56 720 834
use sg13g2_fill_1  FILLER_83_756
timestamp 1677583258
transform 1 0 148224 0 -1 139104
box -48 -56 144 834
use sg13g2_decap_8  FILLER_84_0
timestamp 1679585382
transform 1 0 75648 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_7
timestamp 1679585382
transform 1 0 76320 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_14
timestamp 1679585382
transform 1 0 76992 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_21
timestamp 1679585382
transform 1 0 77664 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_28
timestamp 1679585382
transform 1 0 78336 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_35
timestamp 1679585382
transform 1 0 79008 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_42
timestamp 1679585382
transform 1 0 79680 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_49
timestamp 1679585382
transform 1 0 80352 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_56
timestamp 1679585382
transform 1 0 81024 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_63
timestamp 1679585382
transform 1 0 81696 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_70
timestamp 1679585382
transform 1 0 82368 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_77
timestamp 1679585382
transform 1 0 83040 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_84
timestamp 1679585382
transform 1 0 83712 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_91
timestamp 1679585382
transform 1 0 84384 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_98
timestamp 1679585382
transform 1 0 85056 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_105
timestamp 1679585382
transform 1 0 85728 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_112
timestamp 1679585382
transform 1 0 86400 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_119
timestamp 1679585382
transform 1 0 87072 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_126
timestamp 1679585382
transform 1 0 87744 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_133
timestamp 1679585382
transform 1 0 88416 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_140
timestamp 1679585382
transform 1 0 89088 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_147
timestamp 1679585382
transform 1 0 89760 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_154
timestamp 1679585382
transform 1 0 90432 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_161
timestamp 1679585382
transform 1 0 91104 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_168
timestamp 1679585382
transform 1 0 91776 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_175
timestamp 1679585382
transform 1 0 92448 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_182
timestamp 1679585382
transform 1 0 93120 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_189
timestamp 1679585382
transform 1 0 93792 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_196
timestamp 1679585382
transform 1 0 94464 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_203
timestamp 1679585382
transform 1 0 95136 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_210
timestamp 1679585382
transform 1 0 95808 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_217
timestamp 1679585382
transform 1 0 96480 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_224
timestamp 1679585382
transform 1 0 97152 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_231
timestamp 1679585382
transform 1 0 97824 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_238
timestamp 1679585382
transform 1 0 98496 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_245
timestamp 1679585382
transform 1 0 99168 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_252
timestamp 1679585382
transform 1 0 99840 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_259
timestamp 1679585382
transform 1 0 100512 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_266
timestamp 1679585382
transform 1 0 101184 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_273
timestamp 1679585382
transform 1 0 101856 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_280
timestamp 1679585382
transform 1 0 102528 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_287
timestamp 1679585382
transform 1 0 103200 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_294
timestamp 1679585382
transform 1 0 103872 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_301
timestamp 1679585382
transform 1 0 104544 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_308
timestamp 1679585382
transform 1 0 105216 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_315
timestamp 1679585382
transform 1 0 105888 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_322
timestamp 1679585382
transform 1 0 106560 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_329
timestamp 1679585382
transform 1 0 107232 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_336
timestamp 1679585382
transform 1 0 107904 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_343
timestamp 1679585382
transform 1 0 108576 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_350
timestamp 1679585382
transform 1 0 109248 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_357
timestamp 1679585382
transform 1 0 109920 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_364
timestamp 1679585382
transform 1 0 110592 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_371
timestamp 1679585382
transform 1 0 111264 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_378
timestamp 1679585382
transform 1 0 111936 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_385
timestamp 1679585382
transform 1 0 112608 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_392
timestamp 1679585382
transform 1 0 113280 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_399
timestamp 1679585382
transform 1 0 113952 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_406
timestamp 1679585382
transform 1 0 114624 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_413
timestamp 1679585382
transform 1 0 115296 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_420
timestamp 1679585382
transform 1 0 115968 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_427
timestamp 1679585382
transform 1 0 116640 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_434
timestamp 1679585382
transform 1 0 117312 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_441
timestamp 1679585382
transform 1 0 117984 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_448
timestamp 1679585382
transform 1 0 118656 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_455
timestamp 1679585382
transform 1 0 119328 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_462
timestamp 1679585382
transform 1 0 120000 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_469
timestamp 1679585382
transform 1 0 120672 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_476
timestamp 1679585382
transform 1 0 121344 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_483
timestamp 1679585382
transform 1 0 122016 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_490
timestamp 1679585382
transform 1 0 122688 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_497
timestamp 1679585382
transform 1 0 123360 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_504
timestamp 1679585382
transform 1 0 124032 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_511
timestamp 1679585382
transform 1 0 124704 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_518
timestamp 1679585382
transform 1 0 125376 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_525
timestamp 1679585382
transform 1 0 126048 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_532
timestamp 1679585382
transform 1 0 126720 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_539
timestamp 1679585382
transform 1 0 127392 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_546
timestamp 1679585382
transform 1 0 128064 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_553
timestamp 1679585382
transform 1 0 128736 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_560
timestamp 1679585382
transform 1 0 129408 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_567
timestamp 1679585382
transform 1 0 130080 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_574
timestamp 1679585382
transform 1 0 130752 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_581
timestamp 1679585382
transform 1 0 131424 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_588
timestamp 1679585382
transform 1 0 132096 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_595
timestamp 1679585382
transform 1 0 132768 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_602
timestamp 1679585382
transform 1 0 133440 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_609
timestamp 1679585382
transform 1 0 134112 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_616
timestamp 1679585382
transform 1 0 134784 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_623
timestamp 1679585382
transform 1 0 135456 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_630
timestamp 1679585382
transform 1 0 136128 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_637
timestamp 1679585382
transform 1 0 136800 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_644
timestamp 1679585382
transform 1 0 137472 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_651
timestamp 1679585382
transform 1 0 138144 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_658
timestamp 1679585382
transform 1 0 138816 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_665
timestamp 1679585382
transform 1 0 139488 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_672
timestamp 1679585382
transform 1 0 140160 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_679
timestamp 1679585382
transform 1 0 140832 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_686
timestamp 1679585382
transform 1 0 141504 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_693
timestamp 1679585382
transform 1 0 142176 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_700
timestamp 1679585382
transform 1 0 142848 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_707
timestamp 1679585382
transform 1 0 143520 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_714
timestamp 1679585382
transform 1 0 144192 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_721
timestamp 1679585382
transform 1 0 144864 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_728
timestamp 1679585382
transform 1 0 145536 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_735
timestamp 1679585382
transform 1 0 146208 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_742
timestamp 1679585382
transform 1 0 146880 0 1 139104
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_749
timestamp 1679585382
transform 1 0 147552 0 1 139104
box -48 -56 720 834
use sg13g2_fill_1  FILLER_84_756
timestamp 1677583258
transform 1 0 148224 0 1 139104
box -48 -56 144 834
use sg13g2_decap_8  FILLER_85_0
timestamp 1679585382
transform 1 0 75648 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_7
timestamp 1679585382
transform 1 0 76320 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_14
timestamp 1679585382
transform 1 0 76992 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_21
timestamp 1679585382
transform 1 0 77664 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_28
timestamp 1679585382
transform 1 0 78336 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_35
timestamp 1679585382
transform 1 0 79008 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_42
timestamp 1679585382
transform 1 0 79680 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_49
timestamp 1679585382
transform 1 0 80352 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_56
timestamp 1679585382
transform 1 0 81024 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_63
timestamp 1679585382
transform 1 0 81696 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_70
timestamp 1679585382
transform 1 0 82368 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_77
timestamp 1679585382
transform 1 0 83040 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_84
timestamp 1679585382
transform 1 0 83712 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_91
timestamp 1679585382
transform 1 0 84384 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_98
timestamp 1679585382
transform 1 0 85056 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_105
timestamp 1679585382
transform 1 0 85728 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_112
timestamp 1679585382
transform 1 0 86400 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_119
timestamp 1679585382
transform 1 0 87072 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_126
timestamp 1679585382
transform 1 0 87744 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_133
timestamp 1679585382
transform 1 0 88416 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_140
timestamp 1679585382
transform 1 0 89088 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_147
timestamp 1679585382
transform 1 0 89760 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_154
timestamp 1679585382
transform 1 0 90432 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_161
timestamp 1679585382
transform 1 0 91104 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_168
timestamp 1679585382
transform 1 0 91776 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_175
timestamp 1679585382
transform 1 0 92448 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_182
timestamp 1679585382
transform 1 0 93120 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_189
timestamp 1679585382
transform 1 0 93792 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_196
timestamp 1679585382
transform 1 0 94464 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_203
timestamp 1679585382
transform 1 0 95136 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_210
timestamp 1679585382
transform 1 0 95808 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_217
timestamp 1679585382
transform 1 0 96480 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_224
timestamp 1679585382
transform 1 0 97152 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_231
timestamp 1679585382
transform 1 0 97824 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_238
timestamp 1679585382
transform 1 0 98496 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_245
timestamp 1679585382
transform 1 0 99168 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_252
timestamp 1679585382
transform 1 0 99840 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_259
timestamp 1679585382
transform 1 0 100512 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_266
timestamp 1679585382
transform 1 0 101184 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_273
timestamp 1679585382
transform 1 0 101856 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_280
timestamp 1679585382
transform 1 0 102528 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_287
timestamp 1679585382
transform 1 0 103200 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_294
timestamp 1679585382
transform 1 0 103872 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_301
timestamp 1679585382
transform 1 0 104544 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_308
timestamp 1679585382
transform 1 0 105216 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_315
timestamp 1679585382
transform 1 0 105888 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_322
timestamp 1679585382
transform 1 0 106560 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_329
timestamp 1679585382
transform 1 0 107232 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_336
timestamp 1679585382
transform 1 0 107904 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_343
timestamp 1679585382
transform 1 0 108576 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_350
timestamp 1679585382
transform 1 0 109248 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_357
timestamp 1679585382
transform 1 0 109920 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_364
timestamp 1679585382
transform 1 0 110592 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_371
timestamp 1679585382
transform 1 0 111264 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_378
timestamp 1679585382
transform 1 0 111936 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_385
timestamp 1679585382
transform 1 0 112608 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_392
timestamp 1679585382
transform 1 0 113280 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_399
timestamp 1679585382
transform 1 0 113952 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_406
timestamp 1679585382
transform 1 0 114624 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_413
timestamp 1679585382
transform 1 0 115296 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_420
timestamp 1679585382
transform 1 0 115968 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_427
timestamp 1679585382
transform 1 0 116640 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_434
timestamp 1679585382
transform 1 0 117312 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_441
timestamp 1679585382
transform 1 0 117984 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_448
timestamp 1679585382
transform 1 0 118656 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_455
timestamp 1679585382
transform 1 0 119328 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_462
timestamp 1679585382
transform 1 0 120000 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_469
timestamp 1679585382
transform 1 0 120672 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_476
timestamp 1679585382
transform 1 0 121344 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_483
timestamp 1679585382
transform 1 0 122016 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_490
timestamp 1679585382
transform 1 0 122688 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_497
timestamp 1679585382
transform 1 0 123360 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_504
timestamp 1679585382
transform 1 0 124032 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_511
timestamp 1679585382
transform 1 0 124704 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_518
timestamp 1679585382
transform 1 0 125376 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_525
timestamp 1679585382
transform 1 0 126048 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_532
timestamp 1679585382
transform 1 0 126720 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_539
timestamp 1679585382
transform 1 0 127392 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_546
timestamp 1679585382
transform 1 0 128064 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_553
timestamp 1679585382
transform 1 0 128736 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_560
timestamp 1679585382
transform 1 0 129408 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_567
timestamp 1679585382
transform 1 0 130080 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_574
timestamp 1679585382
transform 1 0 130752 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_581
timestamp 1679585382
transform 1 0 131424 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_588
timestamp 1679585382
transform 1 0 132096 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_595
timestamp 1679585382
transform 1 0 132768 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_602
timestamp 1679585382
transform 1 0 133440 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_609
timestamp 1679585382
transform 1 0 134112 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_616
timestamp 1679585382
transform 1 0 134784 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_623
timestamp 1679585382
transform 1 0 135456 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_630
timestamp 1679585382
transform 1 0 136128 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_637
timestamp 1679585382
transform 1 0 136800 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_644
timestamp 1679585382
transform 1 0 137472 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_651
timestamp 1679585382
transform 1 0 138144 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_658
timestamp 1679585382
transform 1 0 138816 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_665
timestamp 1679585382
transform 1 0 139488 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_672
timestamp 1679585382
transform 1 0 140160 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_679
timestamp 1679585382
transform 1 0 140832 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_686
timestamp 1679585382
transform 1 0 141504 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_693
timestamp 1679585382
transform 1 0 142176 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_700
timestamp 1679585382
transform 1 0 142848 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_707
timestamp 1679585382
transform 1 0 143520 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_714
timestamp 1679585382
transform 1 0 144192 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_721
timestamp 1679585382
transform 1 0 144864 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_728
timestamp 1679585382
transform 1 0 145536 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_735
timestamp 1679585382
transform 1 0 146208 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_742
timestamp 1679585382
transform 1 0 146880 0 -1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_749
timestamp 1679585382
transform 1 0 147552 0 -1 140616
box -48 -56 720 834
use sg13g2_fill_1  FILLER_85_756
timestamp 1677583258
transform 1 0 148224 0 -1 140616
box -48 -56 144 834
use sg13g2_decap_8  FILLER_86_0
timestamp 1679585382
transform 1 0 75648 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_7
timestamp 1679585382
transform 1 0 76320 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_14
timestamp 1679585382
transform 1 0 76992 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_21
timestamp 1679585382
transform 1 0 77664 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_28
timestamp 1679585382
transform 1 0 78336 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_35
timestamp 1679585382
transform 1 0 79008 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_42
timestamp 1679585382
transform 1 0 79680 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_49
timestamp 1679585382
transform 1 0 80352 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_56
timestamp 1679585382
transform 1 0 81024 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_63
timestamp 1679585382
transform 1 0 81696 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_70
timestamp 1679585382
transform 1 0 82368 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_77
timestamp 1679585382
transform 1 0 83040 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_84
timestamp 1679585382
transform 1 0 83712 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_91
timestamp 1679585382
transform 1 0 84384 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_98
timestamp 1679585382
transform 1 0 85056 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_105
timestamp 1679585382
transform 1 0 85728 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_112
timestamp 1679585382
transform 1 0 86400 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_119
timestamp 1679585382
transform 1 0 87072 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_126
timestamp 1679585382
transform 1 0 87744 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_133
timestamp 1679585382
transform 1 0 88416 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_140
timestamp 1679585382
transform 1 0 89088 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_147
timestamp 1679585382
transform 1 0 89760 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_154
timestamp 1679585382
transform 1 0 90432 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_161
timestamp 1679585382
transform 1 0 91104 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_168
timestamp 1679585382
transform 1 0 91776 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_175
timestamp 1679585382
transform 1 0 92448 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_182
timestamp 1679585382
transform 1 0 93120 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_189
timestamp 1679585382
transform 1 0 93792 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_196
timestamp 1679585382
transform 1 0 94464 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_203
timestamp 1679585382
transform 1 0 95136 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_210
timestamp 1679585382
transform 1 0 95808 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_217
timestamp 1679585382
transform 1 0 96480 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_224
timestamp 1679585382
transform 1 0 97152 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_231
timestamp 1679585382
transform 1 0 97824 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_238
timestamp 1679585382
transform 1 0 98496 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_245
timestamp 1679585382
transform 1 0 99168 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_252
timestamp 1679585382
transform 1 0 99840 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_259
timestamp 1679585382
transform 1 0 100512 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_266
timestamp 1679585382
transform 1 0 101184 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_273
timestamp 1679585382
transform 1 0 101856 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_280
timestamp 1679585382
transform 1 0 102528 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_287
timestamp 1679585382
transform 1 0 103200 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_294
timestamp 1679585382
transform 1 0 103872 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_301
timestamp 1679585382
transform 1 0 104544 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_308
timestamp 1679585382
transform 1 0 105216 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_315
timestamp 1679585382
transform 1 0 105888 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_322
timestamp 1679585382
transform 1 0 106560 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_329
timestamp 1679585382
transform 1 0 107232 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_336
timestamp 1679585382
transform 1 0 107904 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_343
timestamp 1679585382
transform 1 0 108576 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_350
timestamp 1679585382
transform 1 0 109248 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_357
timestamp 1679585382
transform 1 0 109920 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_364
timestamp 1679585382
transform 1 0 110592 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_371
timestamp 1679585382
transform 1 0 111264 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_378
timestamp 1679585382
transform 1 0 111936 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_385
timestamp 1679585382
transform 1 0 112608 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_392
timestamp 1679585382
transform 1 0 113280 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_399
timestamp 1679585382
transform 1 0 113952 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_406
timestamp 1679585382
transform 1 0 114624 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_413
timestamp 1679585382
transform 1 0 115296 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_420
timestamp 1679585382
transform 1 0 115968 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_427
timestamp 1679585382
transform 1 0 116640 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_434
timestamp 1679585382
transform 1 0 117312 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_441
timestamp 1679585382
transform 1 0 117984 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_448
timestamp 1679585382
transform 1 0 118656 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_455
timestamp 1679585382
transform 1 0 119328 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_462
timestamp 1679585382
transform 1 0 120000 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_469
timestamp 1679585382
transform 1 0 120672 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_476
timestamp 1679585382
transform 1 0 121344 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_483
timestamp 1679585382
transform 1 0 122016 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_490
timestamp 1679585382
transform 1 0 122688 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_497
timestamp 1679585382
transform 1 0 123360 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_504
timestamp 1679585382
transform 1 0 124032 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_511
timestamp 1679585382
transform 1 0 124704 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_518
timestamp 1679585382
transform 1 0 125376 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_525
timestamp 1679585382
transform 1 0 126048 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_532
timestamp 1679585382
transform 1 0 126720 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_539
timestamp 1679585382
transform 1 0 127392 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_546
timestamp 1679585382
transform 1 0 128064 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_553
timestamp 1679585382
transform 1 0 128736 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_560
timestamp 1679585382
transform 1 0 129408 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_567
timestamp 1679585382
transform 1 0 130080 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_574
timestamp 1679585382
transform 1 0 130752 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_581
timestamp 1679585382
transform 1 0 131424 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_588
timestamp 1679585382
transform 1 0 132096 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_595
timestamp 1679585382
transform 1 0 132768 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_602
timestamp 1679585382
transform 1 0 133440 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_609
timestamp 1679585382
transform 1 0 134112 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_616
timestamp 1679585382
transform 1 0 134784 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_623
timestamp 1679585382
transform 1 0 135456 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_630
timestamp 1679585382
transform 1 0 136128 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_637
timestamp 1679585382
transform 1 0 136800 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_644
timestamp 1679585382
transform 1 0 137472 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_651
timestamp 1679585382
transform 1 0 138144 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_658
timestamp 1679585382
transform 1 0 138816 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_665
timestamp 1679585382
transform 1 0 139488 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_672
timestamp 1679585382
transform 1 0 140160 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_679
timestamp 1679585382
transform 1 0 140832 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_686
timestamp 1679585382
transform 1 0 141504 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_693
timestamp 1679585382
transform 1 0 142176 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_700
timestamp 1679585382
transform 1 0 142848 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_707
timestamp 1679585382
transform 1 0 143520 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_714
timestamp 1679585382
transform 1 0 144192 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_721
timestamp 1679585382
transform 1 0 144864 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_728
timestamp 1679585382
transform 1 0 145536 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_735
timestamp 1679585382
transform 1 0 146208 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_742
timestamp 1679585382
transform 1 0 146880 0 1 140616
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_749
timestamp 1679585382
transform 1 0 147552 0 1 140616
box -48 -56 720 834
use sg13g2_fill_1  FILLER_86_756
timestamp 1677583258
transform 1 0 148224 0 1 140616
box -48 -56 144 834
use sg13g2_decap_8  FILLER_87_0
timestamp 1679585382
transform 1 0 75648 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_7
timestamp 1679585382
transform 1 0 76320 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_14
timestamp 1679585382
transform 1 0 76992 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_21
timestamp 1679585382
transform 1 0 77664 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_28
timestamp 1679585382
transform 1 0 78336 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_35
timestamp 1679585382
transform 1 0 79008 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_42
timestamp 1679585382
transform 1 0 79680 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_49
timestamp 1679585382
transform 1 0 80352 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_56
timestamp 1679585382
transform 1 0 81024 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_63
timestamp 1679585382
transform 1 0 81696 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_70
timestamp 1679585382
transform 1 0 82368 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_77
timestamp 1679585382
transform 1 0 83040 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_84
timestamp 1679585382
transform 1 0 83712 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_91
timestamp 1679585382
transform 1 0 84384 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_98
timestamp 1679585382
transform 1 0 85056 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_105
timestamp 1679585382
transform 1 0 85728 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_112
timestamp 1679585382
transform 1 0 86400 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_119
timestamp 1679585382
transform 1 0 87072 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_126
timestamp 1679585382
transform 1 0 87744 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_133
timestamp 1679585382
transform 1 0 88416 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_140
timestamp 1679585382
transform 1 0 89088 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_147
timestamp 1679585382
transform 1 0 89760 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_154
timestamp 1679585382
transform 1 0 90432 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_161
timestamp 1679585382
transform 1 0 91104 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_168
timestamp 1679585382
transform 1 0 91776 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_175
timestamp 1679585382
transform 1 0 92448 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_182
timestamp 1679585382
transform 1 0 93120 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_189
timestamp 1679585382
transform 1 0 93792 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_196
timestamp 1679585382
transform 1 0 94464 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_203
timestamp 1679585382
transform 1 0 95136 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_210
timestamp 1679585382
transform 1 0 95808 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_217
timestamp 1679585382
transform 1 0 96480 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_224
timestamp 1679585382
transform 1 0 97152 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_231
timestamp 1679585382
transform 1 0 97824 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_238
timestamp 1679585382
transform 1 0 98496 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_245
timestamp 1679585382
transform 1 0 99168 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_252
timestamp 1679585382
transform 1 0 99840 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_259
timestamp 1679585382
transform 1 0 100512 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_266
timestamp 1679585382
transform 1 0 101184 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_273
timestamp 1679585382
transform 1 0 101856 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_280
timestamp 1679585382
transform 1 0 102528 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_287
timestamp 1679585382
transform 1 0 103200 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_294
timestamp 1679585382
transform 1 0 103872 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_301
timestamp 1679585382
transform 1 0 104544 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_308
timestamp 1679585382
transform 1 0 105216 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_315
timestamp 1679585382
transform 1 0 105888 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_322
timestamp 1679585382
transform 1 0 106560 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_329
timestamp 1679585382
transform 1 0 107232 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_336
timestamp 1679585382
transform 1 0 107904 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_343
timestamp 1679585382
transform 1 0 108576 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_350
timestamp 1679585382
transform 1 0 109248 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_357
timestamp 1679585382
transform 1 0 109920 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_364
timestamp 1679585382
transform 1 0 110592 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_371
timestamp 1679585382
transform 1 0 111264 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_378
timestamp 1679585382
transform 1 0 111936 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_385
timestamp 1679585382
transform 1 0 112608 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_392
timestamp 1679585382
transform 1 0 113280 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_399
timestamp 1679585382
transform 1 0 113952 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_406
timestamp 1679585382
transform 1 0 114624 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_413
timestamp 1679585382
transform 1 0 115296 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_420
timestamp 1679585382
transform 1 0 115968 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_427
timestamp 1679585382
transform 1 0 116640 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_434
timestamp 1679585382
transform 1 0 117312 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_441
timestamp 1679585382
transform 1 0 117984 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_448
timestamp 1679585382
transform 1 0 118656 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_455
timestamp 1679585382
transform 1 0 119328 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_462
timestamp 1679585382
transform 1 0 120000 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_469
timestamp 1679585382
transform 1 0 120672 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_476
timestamp 1679585382
transform 1 0 121344 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_483
timestamp 1679585382
transform 1 0 122016 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_490
timestamp 1679585382
transform 1 0 122688 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_497
timestamp 1679585382
transform 1 0 123360 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_504
timestamp 1679585382
transform 1 0 124032 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_511
timestamp 1679585382
transform 1 0 124704 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_518
timestamp 1679585382
transform 1 0 125376 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_525
timestamp 1679585382
transform 1 0 126048 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_532
timestamp 1679585382
transform 1 0 126720 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_539
timestamp 1679585382
transform 1 0 127392 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_546
timestamp 1679585382
transform 1 0 128064 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_553
timestamp 1679585382
transform 1 0 128736 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_560
timestamp 1679585382
transform 1 0 129408 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_567
timestamp 1679585382
transform 1 0 130080 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_574
timestamp 1679585382
transform 1 0 130752 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_581
timestamp 1679585382
transform 1 0 131424 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_588
timestamp 1679585382
transform 1 0 132096 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_595
timestamp 1679585382
transform 1 0 132768 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_602
timestamp 1679585382
transform 1 0 133440 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_609
timestamp 1679585382
transform 1 0 134112 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_616
timestamp 1679585382
transform 1 0 134784 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_623
timestamp 1679585382
transform 1 0 135456 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_630
timestamp 1679585382
transform 1 0 136128 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_637
timestamp 1679585382
transform 1 0 136800 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_644
timestamp 1679585382
transform 1 0 137472 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_651
timestamp 1679585382
transform 1 0 138144 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_658
timestamp 1679585382
transform 1 0 138816 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_665
timestamp 1679585382
transform 1 0 139488 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_672
timestamp 1679585382
transform 1 0 140160 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_679
timestamp 1679585382
transform 1 0 140832 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_686
timestamp 1679585382
transform 1 0 141504 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_693
timestamp 1679585382
transform 1 0 142176 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_700
timestamp 1679585382
transform 1 0 142848 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_707
timestamp 1679585382
transform 1 0 143520 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_714
timestamp 1679585382
transform 1 0 144192 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_721
timestamp 1679585382
transform 1 0 144864 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_728
timestamp 1679585382
transform 1 0 145536 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_735
timestamp 1679585382
transform 1 0 146208 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_742
timestamp 1679585382
transform 1 0 146880 0 -1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_87_749
timestamp 1679585382
transform 1 0 147552 0 -1 142128
box -48 -56 720 834
use sg13g2_fill_1  FILLER_87_756
timestamp 1677583258
transform 1 0 148224 0 -1 142128
box -48 -56 144 834
use sg13g2_decap_8  FILLER_88_0
timestamp 1679585382
transform 1 0 75648 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_7
timestamp 1679585382
transform 1 0 76320 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_14
timestamp 1679585382
transform 1 0 76992 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_21
timestamp 1679585382
transform 1 0 77664 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_28
timestamp 1679585382
transform 1 0 78336 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_35
timestamp 1679585382
transform 1 0 79008 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_42
timestamp 1679585382
transform 1 0 79680 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_49
timestamp 1679585382
transform 1 0 80352 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_56
timestamp 1679585382
transform 1 0 81024 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_63
timestamp 1679585382
transform 1 0 81696 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_70
timestamp 1679585382
transform 1 0 82368 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_77
timestamp 1679585382
transform 1 0 83040 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_84
timestamp 1679585382
transform 1 0 83712 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_91
timestamp 1679585382
transform 1 0 84384 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_98
timestamp 1679585382
transform 1 0 85056 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_105
timestamp 1679585382
transform 1 0 85728 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_112
timestamp 1679585382
transform 1 0 86400 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_119
timestamp 1679585382
transform 1 0 87072 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_126
timestamp 1679585382
transform 1 0 87744 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_133
timestamp 1679585382
transform 1 0 88416 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_140
timestamp 1679585382
transform 1 0 89088 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_147
timestamp 1679585382
transform 1 0 89760 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_154
timestamp 1679585382
transform 1 0 90432 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_161
timestamp 1679585382
transform 1 0 91104 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_168
timestamp 1679585382
transform 1 0 91776 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_175
timestamp 1679585382
transform 1 0 92448 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_182
timestamp 1679585382
transform 1 0 93120 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_189
timestamp 1679585382
transform 1 0 93792 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_196
timestamp 1679585382
transform 1 0 94464 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_203
timestamp 1679585382
transform 1 0 95136 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_210
timestamp 1679585382
transform 1 0 95808 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_217
timestamp 1679585382
transform 1 0 96480 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_224
timestamp 1679585382
transform 1 0 97152 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_231
timestamp 1679585382
transform 1 0 97824 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_238
timestamp 1679585382
transform 1 0 98496 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_245
timestamp 1679585382
transform 1 0 99168 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_252
timestamp 1679585382
transform 1 0 99840 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_259
timestamp 1679585382
transform 1 0 100512 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_266
timestamp 1679585382
transform 1 0 101184 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_273
timestamp 1679585382
transform 1 0 101856 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_280
timestamp 1679585382
transform 1 0 102528 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_287
timestamp 1679585382
transform 1 0 103200 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_294
timestamp 1679585382
transform 1 0 103872 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_301
timestamp 1679585382
transform 1 0 104544 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_308
timestamp 1679585382
transform 1 0 105216 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_315
timestamp 1679585382
transform 1 0 105888 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_322
timestamp 1679585382
transform 1 0 106560 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_329
timestamp 1679585382
transform 1 0 107232 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_336
timestamp 1679585382
transform 1 0 107904 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_343
timestamp 1679585382
transform 1 0 108576 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_350
timestamp 1679585382
transform 1 0 109248 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_357
timestamp 1679585382
transform 1 0 109920 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_364
timestamp 1679585382
transform 1 0 110592 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_371
timestamp 1679585382
transform 1 0 111264 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_378
timestamp 1679585382
transform 1 0 111936 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_385
timestamp 1679585382
transform 1 0 112608 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_392
timestamp 1679585382
transform 1 0 113280 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_399
timestamp 1679585382
transform 1 0 113952 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_406
timestamp 1679585382
transform 1 0 114624 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_413
timestamp 1679585382
transform 1 0 115296 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_420
timestamp 1679585382
transform 1 0 115968 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_427
timestamp 1679585382
transform 1 0 116640 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_434
timestamp 1679585382
transform 1 0 117312 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_441
timestamp 1679585382
transform 1 0 117984 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_448
timestamp 1679585382
transform 1 0 118656 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_455
timestamp 1679585382
transform 1 0 119328 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_462
timestamp 1679585382
transform 1 0 120000 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_469
timestamp 1679585382
transform 1 0 120672 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_476
timestamp 1679585382
transform 1 0 121344 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_483
timestamp 1679585382
transform 1 0 122016 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_490
timestamp 1679585382
transform 1 0 122688 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_497
timestamp 1679585382
transform 1 0 123360 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_504
timestamp 1679585382
transform 1 0 124032 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_511
timestamp 1679585382
transform 1 0 124704 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_518
timestamp 1679585382
transform 1 0 125376 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_525
timestamp 1679585382
transform 1 0 126048 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_532
timestamp 1679585382
transform 1 0 126720 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_539
timestamp 1679585382
transform 1 0 127392 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_546
timestamp 1679585382
transform 1 0 128064 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_553
timestamp 1679585382
transform 1 0 128736 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_560
timestamp 1679585382
transform 1 0 129408 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_567
timestamp 1679585382
transform 1 0 130080 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_574
timestamp 1679585382
transform 1 0 130752 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_581
timestamp 1679585382
transform 1 0 131424 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_588
timestamp 1679585382
transform 1 0 132096 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_595
timestamp 1679585382
transform 1 0 132768 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_602
timestamp 1679585382
transform 1 0 133440 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_609
timestamp 1679585382
transform 1 0 134112 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_616
timestamp 1679585382
transform 1 0 134784 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_623
timestamp 1679585382
transform 1 0 135456 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_630
timestamp 1679585382
transform 1 0 136128 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_637
timestamp 1679585382
transform 1 0 136800 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_644
timestamp 1679585382
transform 1 0 137472 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_651
timestamp 1679585382
transform 1 0 138144 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_658
timestamp 1679585382
transform 1 0 138816 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_665
timestamp 1679585382
transform 1 0 139488 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_672
timestamp 1679585382
transform 1 0 140160 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_679
timestamp 1679585382
transform 1 0 140832 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_686
timestamp 1679585382
transform 1 0 141504 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_693
timestamp 1679585382
transform 1 0 142176 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_700
timestamp 1679585382
transform 1 0 142848 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_707
timestamp 1679585382
transform 1 0 143520 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_714
timestamp 1679585382
transform 1 0 144192 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_721
timestamp 1679585382
transform 1 0 144864 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_728
timestamp 1679585382
transform 1 0 145536 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_735
timestamp 1679585382
transform 1 0 146208 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_742
timestamp 1679585382
transform 1 0 146880 0 1 142128
box -48 -56 720 834
use sg13g2_decap_8  FILLER_88_749
timestamp 1679585382
transform 1 0 147552 0 1 142128
box -48 -56 720 834
use sg13g2_fill_1  FILLER_88_756
timestamp 1677583258
transform 1 0 148224 0 1 142128
box -48 -56 144 834
use sg13g2_decap_8  FILLER_89_0
timestamp 1679585382
transform 1 0 75648 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_7
timestamp 1679585382
transform 1 0 76320 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_14
timestamp 1679585382
transform 1 0 76992 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_21
timestamp 1679585382
transform 1 0 77664 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_28
timestamp 1679585382
transform 1 0 78336 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_35
timestamp 1679585382
transform 1 0 79008 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_42
timestamp 1679585382
transform 1 0 79680 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_49
timestamp 1679585382
transform 1 0 80352 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_56
timestamp 1679585382
transform 1 0 81024 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_63
timestamp 1679585382
transform 1 0 81696 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_70
timestamp 1679585382
transform 1 0 82368 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_77
timestamp 1679585382
transform 1 0 83040 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_84
timestamp 1679585382
transform 1 0 83712 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_91
timestamp 1679585382
transform 1 0 84384 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_98
timestamp 1679585382
transform 1 0 85056 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_105
timestamp 1679585382
transform 1 0 85728 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_112
timestamp 1679585382
transform 1 0 86400 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_119
timestamp 1679585382
transform 1 0 87072 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_126
timestamp 1679585382
transform 1 0 87744 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_133
timestamp 1679585382
transform 1 0 88416 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_140
timestamp 1679585382
transform 1 0 89088 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_147
timestamp 1679585382
transform 1 0 89760 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_154
timestamp 1679585382
transform 1 0 90432 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_161
timestamp 1679585382
transform 1 0 91104 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_168
timestamp 1679585382
transform 1 0 91776 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_175
timestamp 1679585382
transform 1 0 92448 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_182
timestamp 1679585382
transform 1 0 93120 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_189
timestamp 1679585382
transform 1 0 93792 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_196
timestamp 1679585382
transform 1 0 94464 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_203
timestamp 1679585382
transform 1 0 95136 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_210
timestamp 1679585382
transform 1 0 95808 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_217
timestamp 1679585382
transform 1 0 96480 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_224
timestamp 1679585382
transform 1 0 97152 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_231
timestamp 1679585382
transform 1 0 97824 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_238
timestamp 1679585382
transform 1 0 98496 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_245
timestamp 1679585382
transform 1 0 99168 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_252
timestamp 1679585382
transform 1 0 99840 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_259
timestamp 1679585382
transform 1 0 100512 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_266
timestamp 1679585382
transform 1 0 101184 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_273
timestamp 1679585382
transform 1 0 101856 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_280
timestamp 1679585382
transform 1 0 102528 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_287
timestamp 1679585382
transform 1 0 103200 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_294
timestamp 1679585382
transform 1 0 103872 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_301
timestamp 1679585382
transform 1 0 104544 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_308
timestamp 1679585382
transform 1 0 105216 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_315
timestamp 1679585382
transform 1 0 105888 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_322
timestamp 1679585382
transform 1 0 106560 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_329
timestamp 1679585382
transform 1 0 107232 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_336
timestamp 1679585382
transform 1 0 107904 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_343
timestamp 1679585382
transform 1 0 108576 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_350
timestamp 1679585382
transform 1 0 109248 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_357
timestamp 1679585382
transform 1 0 109920 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_364
timestamp 1679585382
transform 1 0 110592 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_371
timestamp 1679585382
transform 1 0 111264 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_378
timestamp 1679585382
transform 1 0 111936 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_385
timestamp 1679585382
transform 1 0 112608 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_392
timestamp 1679585382
transform 1 0 113280 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_399
timestamp 1679585382
transform 1 0 113952 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_406
timestamp 1679585382
transform 1 0 114624 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_413
timestamp 1679585382
transform 1 0 115296 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_420
timestamp 1679585382
transform 1 0 115968 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_427
timestamp 1679585382
transform 1 0 116640 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_434
timestamp 1679585382
transform 1 0 117312 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_441
timestamp 1679585382
transform 1 0 117984 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_448
timestamp 1679585382
transform 1 0 118656 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_455
timestamp 1679585382
transform 1 0 119328 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_462
timestamp 1679585382
transform 1 0 120000 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_469
timestamp 1679585382
transform 1 0 120672 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_476
timestamp 1679585382
transform 1 0 121344 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_483
timestamp 1679585382
transform 1 0 122016 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_490
timestamp 1679585382
transform 1 0 122688 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_497
timestamp 1679585382
transform 1 0 123360 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_504
timestamp 1679585382
transform 1 0 124032 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_511
timestamp 1679585382
transform 1 0 124704 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_518
timestamp 1679585382
transform 1 0 125376 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_525
timestamp 1679585382
transform 1 0 126048 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_532
timestamp 1679585382
transform 1 0 126720 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_539
timestamp 1679585382
transform 1 0 127392 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_546
timestamp 1679585382
transform 1 0 128064 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_553
timestamp 1679585382
transform 1 0 128736 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_560
timestamp 1679585382
transform 1 0 129408 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_567
timestamp 1679585382
transform 1 0 130080 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_574
timestamp 1679585382
transform 1 0 130752 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_581
timestamp 1679585382
transform 1 0 131424 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_588
timestamp 1679585382
transform 1 0 132096 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_595
timestamp 1679585382
transform 1 0 132768 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_602
timestamp 1679585382
transform 1 0 133440 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_609
timestamp 1679585382
transform 1 0 134112 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_616
timestamp 1679585382
transform 1 0 134784 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_623
timestamp 1679585382
transform 1 0 135456 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_630
timestamp 1679585382
transform 1 0 136128 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_637
timestamp 1679585382
transform 1 0 136800 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_644
timestamp 1679585382
transform 1 0 137472 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_651
timestamp 1679585382
transform 1 0 138144 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_658
timestamp 1679585382
transform 1 0 138816 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_665
timestamp 1679585382
transform 1 0 139488 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_672
timestamp 1679585382
transform 1 0 140160 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_679
timestamp 1679585382
transform 1 0 140832 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_686
timestamp 1679585382
transform 1 0 141504 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_693
timestamp 1679585382
transform 1 0 142176 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_700
timestamp 1679585382
transform 1 0 142848 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_707
timestamp 1679585382
transform 1 0 143520 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_714
timestamp 1679585382
transform 1 0 144192 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_721
timestamp 1679585382
transform 1 0 144864 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_728
timestamp 1679585382
transform 1 0 145536 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_735
timestamp 1679585382
transform 1 0 146208 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_742
timestamp 1679585382
transform 1 0 146880 0 -1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_89_749
timestamp 1679585382
transform 1 0 147552 0 -1 143640
box -48 -56 720 834
use sg13g2_fill_1  FILLER_89_756
timestamp 1677583258
transform 1 0 148224 0 -1 143640
box -48 -56 144 834
use sg13g2_decap_8  FILLER_90_0
timestamp 1679585382
transform 1 0 75648 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_7
timestamp 1679585382
transform 1 0 76320 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_14
timestamp 1679585382
transform 1 0 76992 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_21
timestamp 1679585382
transform 1 0 77664 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_28
timestamp 1679585382
transform 1 0 78336 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_35
timestamp 1679585382
transform 1 0 79008 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_42
timestamp 1679585382
transform 1 0 79680 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_49
timestamp 1679585382
transform 1 0 80352 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_56
timestamp 1679585382
transform 1 0 81024 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_63
timestamp 1679585382
transform 1 0 81696 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_70
timestamp 1679585382
transform 1 0 82368 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_77
timestamp 1679585382
transform 1 0 83040 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_84
timestamp 1679585382
transform 1 0 83712 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_91
timestamp 1679585382
transform 1 0 84384 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_98
timestamp 1679585382
transform 1 0 85056 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_105
timestamp 1679585382
transform 1 0 85728 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_112
timestamp 1679585382
transform 1 0 86400 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_119
timestamp 1679585382
transform 1 0 87072 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_126
timestamp 1679585382
transform 1 0 87744 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_133
timestamp 1679585382
transform 1 0 88416 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_140
timestamp 1679585382
transform 1 0 89088 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_147
timestamp 1679585382
transform 1 0 89760 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_154
timestamp 1679585382
transform 1 0 90432 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_161
timestamp 1679585382
transform 1 0 91104 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_168
timestamp 1679585382
transform 1 0 91776 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_175
timestamp 1679585382
transform 1 0 92448 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_182
timestamp 1679585382
transform 1 0 93120 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_189
timestamp 1679585382
transform 1 0 93792 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_196
timestamp 1679585382
transform 1 0 94464 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_203
timestamp 1679585382
transform 1 0 95136 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_210
timestamp 1679585382
transform 1 0 95808 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_217
timestamp 1679585382
transform 1 0 96480 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_224
timestamp 1679585382
transform 1 0 97152 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_231
timestamp 1679585382
transform 1 0 97824 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_238
timestamp 1679585382
transform 1 0 98496 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_245
timestamp 1679585382
transform 1 0 99168 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_252
timestamp 1679585382
transform 1 0 99840 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_259
timestamp 1679585382
transform 1 0 100512 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_266
timestamp 1679585382
transform 1 0 101184 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_273
timestamp 1679585382
transform 1 0 101856 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_280
timestamp 1679585382
transform 1 0 102528 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_287
timestamp 1679585382
transform 1 0 103200 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_294
timestamp 1679585382
transform 1 0 103872 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_301
timestamp 1679585382
transform 1 0 104544 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_308
timestamp 1679585382
transform 1 0 105216 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_315
timestamp 1679585382
transform 1 0 105888 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_322
timestamp 1679585382
transform 1 0 106560 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_329
timestamp 1679585382
transform 1 0 107232 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_336
timestamp 1679585382
transform 1 0 107904 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_343
timestamp 1679585382
transform 1 0 108576 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_350
timestamp 1679585382
transform 1 0 109248 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_357
timestamp 1679585382
transform 1 0 109920 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_364
timestamp 1679585382
transform 1 0 110592 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_371
timestamp 1679585382
transform 1 0 111264 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_378
timestamp 1679585382
transform 1 0 111936 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_385
timestamp 1679585382
transform 1 0 112608 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_392
timestamp 1679585382
transform 1 0 113280 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_399
timestamp 1679585382
transform 1 0 113952 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_406
timestamp 1679585382
transform 1 0 114624 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_413
timestamp 1679585382
transform 1 0 115296 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_420
timestamp 1679585382
transform 1 0 115968 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_427
timestamp 1679585382
transform 1 0 116640 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_434
timestamp 1679585382
transform 1 0 117312 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_441
timestamp 1679585382
transform 1 0 117984 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_448
timestamp 1679585382
transform 1 0 118656 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_455
timestamp 1679585382
transform 1 0 119328 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_462
timestamp 1679585382
transform 1 0 120000 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_469
timestamp 1679585382
transform 1 0 120672 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_476
timestamp 1679585382
transform 1 0 121344 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_483
timestamp 1679585382
transform 1 0 122016 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_490
timestamp 1679585382
transform 1 0 122688 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_497
timestamp 1679585382
transform 1 0 123360 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_504
timestamp 1679585382
transform 1 0 124032 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_511
timestamp 1679585382
transform 1 0 124704 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_518
timestamp 1679585382
transform 1 0 125376 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_525
timestamp 1679585382
transform 1 0 126048 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_532
timestamp 1679585382
transform 1 0 126720 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_539
timestamp 1679585382
transform 1 0 127392 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_546
timestamp 1679585382
transform 1 0 128064 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_553
timestamp 1679585382
transform 1 0 128736 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_560
timestamp 1679585382
transform 1 0 129408 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_567
timestamp 1679585382
transform 1 0 130080 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_574
timestamp 1679585382
transform 1 0 130752 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_581
timestamp 1679585382
transform 1 0 131424 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_588
timestamp 1679585382
transform 1 0 132096 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_595
timestamp 1679585382
transform 1 0 132768 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_602
timestamp 1679585382
transform 1 0 133440 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_609
timestamp 1679585382
transform 1 0 134112 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_616
timestamp 1679585382
transform 1 0 134784 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_623
timestamp 1679585382
transform 1 0 135456 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_630
timestamp 1679585382
transform 1 0 136128 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_637
timestamp 1679585382
transform 1 0 136800 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_644
timestamp 1679585382
transform 1 0 137472 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_651
timestamp 1679585382
transform 1 0 138144 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_658
timestamp 1679585382
transform 1 0 138816 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_665
timestamp 1679585382
transform 1 0 139488 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_672
timestamp 1679585382
transform 1 0 140160 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_679
timestamp 1679585382
transform 1 0 140832 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_686
timestamp 1679585382
transform 1 0 141504 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_693
timestamp 1679585382
transform 1 0 142176 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_700
timestamp 1679585382
transform 1 0 142848 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_707
timestamp 1679585382
transform 1 0 143520 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_714
timestamp 1679585382
transform 1 0 144192 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_721
timestamp 1679585382
transform 1 0 144864 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_728
timestamp 1679585382
transform 1 0 145536 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_735
timestamp 1679585382
transform 1 0 146208 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_742
timestamp 1679585382
transform 1 0 146880 0 1 143640
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_749
timestamp 1679585382
transform 1 0 147552 0 1 143640
box -48 -56 720 834
use sg13g2_fill_1  FILLER_90_756
timestamp 1677583258
transform 1 0 148224 0 1 143640
box -48 -56 144 834
use sg13g2_decap_8  FILLER_91_0
timestamp 1679585382
transform 1 0 75648 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_7
timestamp 1679585382
transform 1 0 76320 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_14
timestamp 1679585382
transform 1 0 76992 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_21
timestamp 1679585382
transform 1 0 77664 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_28
timestamp 1679585382
transform 1 0 78336 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_35
timestamp 1679585382
transform 1 0 79008 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_42
timestamp 1679585382
transform 1 0 79680 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_49
timestamp 1679585382
transform 1 0 80352 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_56
timestamp 1679585382
transform 1 0 81024 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_63
timestamp 1679585382
transform 1 0 81696 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_70
timestamp 1679585382
transform 1 0 82368 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_77
timestamp 1679585382
transform 1 0 83040 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_84
timestamp 1679585382
transform 1 0 83712 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_91
timestamp 1679585382
transform 1 0 84384 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_98
timestamp 1679585382
transform 1 0 85056 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_105
timestamp 1679585382
transform 1 0 85728 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_112
timestamp 1679585382
transform 1 0 86400 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_119
timestamp 1679585382
transform 1 0 87072 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_126
timestamp 1679585382
transform 1 0 87744 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_133
timestamp 1679585382
transform 1 0 88416 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_140
timestamp 1679585382
transform 1 0 89088 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_147
timestamp 1679585382
transform 1 0 89760 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_154
timestamp 1679585382
transform 1 0 90432 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_161
timestamp 1679585382
transform 1 0 91104 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_168
timestamp 1679585382
transform 1 0 91776 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_175
timestamp 1679585382
transform 1 0 92448 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_182
timestamp 1679585382
transform 1 0 93120 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_189
timestamp 1679585382
transform 1 0 93792 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_196
timestamp 1679585382
transform 1 0 94464 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_203
timestamp 1679585382
transform 1 0 95136 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_210
timestamp 1679585382
transform 1 0 95808 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_217
timestamp 1679585382
transform 1 0 96480 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_224
timestamp 1679585382
transform 1 0 97152 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_231
timestamp 1679585382
transform 1 0 97824 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_238
timestamp 1679585382
transform 1 0 98496 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_245
timestamp 1679585382
transform 1 0 99168 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_252
timestamp 1679585382
transform 1 0 99840 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_259
timestamp 1679585382
transform 1 0 100512 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_266
timestamp 1679585382
transform 1 0 101184 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_273
timestamp 1679585382
transform 1 0 101856 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_280
timestamp 1679585382
transform 1 0 102528 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_287
timestamp 1679585382
transform 1 0 103200 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_294
timestamp 1679585382
transform 1 0 103872 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_301
timestamp 1679585382
transform 1 0 104544 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_308
timestamp 1679585382
transform 1 0 105216 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_315
timestamp 1679585382
transform 1 0 105888 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_322
timestamp 1679585382
transform 1 0 106560 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_329
timestamp 1679585382
transform 1 0 107232 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_336
timestamp 1679585382
transform 1 0 107904 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_343
timestamp 1679585382
transform 1 0 108576 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_350
timestamp 1679585382
transform 1 0 109248 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_357
timestamp 1679585382
transform 1 0 109920 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_364
timestamp 1679585382
transform 1 0 110592 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_371
timestamp 1679585382
transform 1 0 111264 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_378
timestamp 1679585382
transform 1 0 111936 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_385
timestamp 1679585382
transform 1 0 112608 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_392
timestamp 1679585382
transform 1 0 113280 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_399
timestamp 1679585382
transform 1 0 113952 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_406
timestamp 1679585382
transform 1 0 114624 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_413
timestamp 1679585382
transform 1 0 115296 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_420
timestamp 1679585382
transform 1 0 115968 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_427
timestamp 1679585382
transform 1 0 116640 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_434
timestamp 1679585382
transform 1 0 117312 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_441
timestamp 1679585382
transform 1 0 117984 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_448
timestamp 1679585382
transform 1 0 118656 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_455
timestamp 1679585382
transform 1 0 119328 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_462
timestamp 1679585382
transform 1 0 120000 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_469
timestamp 1679585382
transform 1 0 120672 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_476
timestamp 1679585382
transform 1 0 121344 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_483
timestamp 1679585382
transform 1 0 122016 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_490
timestamp 1679585382
transform 1 0 122688 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_497
timestamp 1679585382
transform 1 0 123360 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_504
timestamp 1679585382
transform 1 0 124032 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_511
timestamp 1679585382
transform 1 0 124704 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_518
timestamp 1679585382
transform 1 0 125376 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_525
timestamp 1679585382
transform 1 0 126048 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_532
timestamp 1679585382
transform 1 0 126720 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_539
timestamp 1679585382
transform 1 0 127392 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_546
timestamp 1679585382
transform 1 0 128064 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_553
timestamp 1679585382
transform 1 0 128736 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_560
timestamp 1679585382
transform 1 0 129408 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_567
timestamp 1679585382
transform 1 0 130080 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_574
timestamp 1679585382
transform 1 0 130752 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_581
timestamp 1679585382
transform 1 0 131424 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_588
timestamp 1679585382
transform 1 0 132096 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_595
timestamp 1679585382
transform 1 0 132768 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_602
timestamp 1679585382
transform 1 0 133440 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_609
timestamp 1679585382
transform 1 0 134112 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_616
timestamp 1679585382
transform 1 0 134784 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_623
timestamp 1679585382
transform 1 0 135456 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_630
timestamp 1679585382
transform 1 0 136128 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_637
timestamp 1679585382
transform 1 0 136800 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_644
timestamp 1679585382
transform 1 0 137472 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_651
timestamp 1679585382
transform 1 0 138144 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_658
timestamp 1679585382
transform 1 0 138816 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_665
timestamp 1679585382
transform 1 0 139488 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_672
timestamp 1679585382
transform 1 0 140160 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_679
timestamp 1679585382
transform 1 0 140832 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_686
timestamp 1679585382
transform 1 0 141504 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_693
timestamp 1679585382
transform 1 0 142176 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_700
timestamp 1679585382
transform 1 0 142848 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_707
timestamp 1679585382
transform 1 0 143520 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_714
timestamp 1679585382
transform 1 0 144192 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_721
timestamp 1679585382
transform 1 0 144864 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_728
timestamp 1679585382
transform 1 0 145536 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_735
timestamp 1679585382
transform 1 0 146208 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_742
timestamp 1679585382
transform 1 0 146880 0 -1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_91_749
timestamp 1679585382
transform 1 0 147552 0 -1 145152
box -48 -56 720 834
use sg13g2_fill_1  FILLER_91_756
timestamp 1677583258
transform 1 0 148224 0 -1 145152
box -48 -56 144 834
use sg13g2_decap_8  FILLER_92_0
timestamp 1679585382
transform 1 0 75648 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_7
timestamp 1679585382
transform 1 0 76320 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_14
timestamp 1679585382
transform 1 0 76992 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_21
timestamp 1679585382
transform 1 0 77664 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_28
timestamp 1679585382
transform 1 0 78336 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_35
timestamp 1679585382
transform 1 0 79008 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_42
timestamp 1679585382
transform 1 0 79680 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_49
timestamp 1679585382
transform 1 0 80352 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_56
timestamp 1679585382
transform 1 0 81024 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_63
timestamp 1679585382
transform 1 0 81696 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_70
timestamp 1679585382
transform 1 0 82368 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_77
timestamp 1679585382
transform 1 0 83040 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_84
timestamp 1679585382
transform 1 0 83712 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_91
timestamp 1679585382
transform 1 0 84384 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_98
timestamp 1679585382
transform 1 0 85056 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_105
timestamp 1679585382
transform 1 0 85728 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_112
timestamp 1679585382
transform 1 0 86400 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_119
timestamp 1679585382
transform 1 0 87072 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_126
timestamp 1679585382
transform 1 0 87744 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_133
timestamp 1679585382
transform 1 0 88416 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_140
timestamp 1679585382
transform 1 0 89088 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_147
timestamp 1679585382
transform 1 0 89760 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_154
timestamp 1679585382
transform 1 0 90432 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_161
timestamp 1679585382
transform 1 0 91104 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_168
timestamp 1679585382
transform 1 0 91776 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_175
timestamp 1679585382
transform 1 0 92448 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_182
timestamp 1679585382
transform 1 0 93120 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_189
timestamp 1679585382
transform 1 0 93792 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_196
timestamp 1679585382
transform 1 0 94464 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_203
timestamp 1679585382
transform 1 0 95136 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_210
timestamp 1679585382
transform 1 0 95808 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_217
timestamp 1679585382
transform 1 0 96480 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_224
timestamp 1679585382
transform 1 0 97152 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_231
timestamp 1679585382
transform 1 0 97824 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_238
timestamp 1679585382
transform 1 0 98496 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_245
timestamp 1679585382
transform 1 0 99168 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_252
timestamp 1679585382
transform 1 0 99840 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_259
timestamp 1679585382
transform 1 0 100512 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_266
timestamp 1679585382
transform 1 0 101184 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_273
timestamp 1679585382
transform 1 0 101856 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_280
timestamp 1679585382
transform 1 0 102528 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_287
timestamp 1679585382
transform 1 0 103200 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_294
timestamp 1679585382
transform 1 0 103872 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_301
timestamp 1679585382
transform 1 0 104544 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_308
timestamp 1679585382
transform 1 0 105216 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_315
timestamp 1679585382
transform 1 0 105888 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_322
timestamp 1679585382
transform 1 0 106560 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_329
timestamp 1679585382
transform 1 0 107232 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_336
timestamp 1679585382
transform 1 0 107904 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_343
timestamp 1679585382
transform 1 0 108576 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_350
timestamp 1679585382
transform 1 0 109248 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_357
timestamp 1679585382
transform 1 0 109920 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_364
timestamp 1679585382
transform 1 0 110592 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_371
timestamp 1679585382
transform 1 0 111264 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_378
timestamp 1679585382
transform 1 0 111936 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_385
timestamp 1679585382
transform 1 0 112608 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_392
timestamp 1679585382
transform 1 0 113280 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_399
timestamp 1679585382
transform 1 0 113952 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_406
timestamp 1679585382
transform 1 0 114624 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_413
timestamp 1679585382
transform 1 0 115296 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_420
timestamp 1679585382
transform 1 0 115968 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_427
timestamp 1679585382
transform 1 0 116640 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_434
timestamp 1679585382
transform 1 0 117312 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_441
timestamp 1679585382
transform 1 0 117984 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_448
timestamp 1679585382
transform 1 0 118656 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_455
timestamp 1679585382
transform 1 0 119328 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_462
timestamp 1679585382
transform 1 0 120000 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_469
timestamp 1679585382
transform 1 0 120672 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_476
timestamp 1679585382
transform 1 0 121344 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_483
timestamp 1679585382
transform 1 0 122016 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_490
timestamp 1679585382
transform 1 0 122688 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_497
timestamp 1679585382
transform 1 0 123360 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_504
timestamp 1679585382
transform 1 0 124032 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_511
timestamp 1679585382
transform 1 0 124704 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_518
timestamp 1679585382
transform 1 0 125376 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_525
timestamp 1679585382
transform 1 0 126048 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_532
timestamp 1679585382
transform 1 0 126720 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_539
timestamp 1679585382
transform 1 0 127392 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_546
timestamp 1679585382
transform 1 0 128064 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_553
timestamp 1679585382
transform 1 0 128736 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_560
timestamp 1679585382
transform 1 0 129408 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_567
timestamp 1679585382
transform 1 0 130080 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_574
timestamp 1679585382
transform 1 0 130752 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_581
timestamp 1679585382
transform 1 0 131424 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_588
timestamp 1679585382
transform 1 0 132096 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_595
timestamp 1679585382
transform 1 0 132768 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_602
timestamp 1679585382
transform 1 0 133440 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_609
timestamp 1679585382
transform 1 0 134112 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_616
timestamp 1679585382
transform 1 0 134784 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_623
timestamp 1679585382
transform 1 0 135456 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_630
timestamp 1679585382
transform 1 0 136128 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_637
timestamp 1679585382
transform 1 0 136800 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_644
timestamp 1679585382
transform 1 0 137472 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_651
timestamp 1679585382
transform 1 0 138144 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_658
timestamp 1679585382
transform 1 0 138816 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_665
timestamp 1679585382
transform 1 0 139488 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_672
timestamp 1679585382
transform 1 0 140160 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_679
timestamp 1679585382
transform 1 0 140832 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_686
timestamp 1679585382
transform 1 0 141504 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_693
timestamp 1679585382
transform 1 0 142176 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_700
timestamp 1679585382
transform 1 0 142848 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_707
timestamp 1679585382
transform 1 0 143520 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_714
timestamp 1679585382
transform 1 0 144192 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_721
timestamp 1679585382
transform 1 0 144864 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_728
timestamp 1679585382
transform 1 0 145536 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_735
timestamp 1679585382
transform 1 0 146208 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_742
timestamp 1679585382
transform 1 0 146880 0 1 145152
box -48 -56 720 834
use sg13g2_decap_8  FILLER_92_749
timestamp 1679585382
transform 1 0 147552 0 1 145152
box -48 -56 720 834
use sg13g2_fill_1  FILLER_92_756
timestamp 1677583258
transform 1 0 148224 0 1 145152
box -48 -56 144 834
use sg13g2_decap_8  FILLER_93_0
timestamp 1679585382
transform 1 0 75648 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_7
timestamp 1679585382
transform 1 0 76320 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_14
timestamp 1679585382
transform 1 0 76992 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_21
timestamp 1679585382
transform 1 0 77664 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_28
timestamp 1679585382
transform 1 0 78336 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_35
timestamp 1679585382
transform 1 0 79008 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_42
timestamp 1679585382
transform 1 0 79680 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_49
timestamp 1679585382
transform 1 0 80352 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_56
timestamp 1679585382
transform 1 0 81024 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_63
timestamp 1679585382
transform 1 0 81696 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_70
timestamp 1679585382
transform 1 0 82368 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_77
timestamp 1679585382
transform 1 0 83040 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_84
timestamp 1679585382
transform 1 0 83712 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_91
timestamp 1679585382
transform 1 0 84384 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_98
timestamp 1679585382
transform 1 0 85056 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_105
timestamp 1679585382
transform 1 0 85728 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_112
timestamp 1679585382
transform 1 0 86400 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_119
timestamp 1679585382
transform 1 0 87072 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_126
timestamp 1679585382
transform 1 0 87744 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_133
timestamp 1679585382
transform 1 0 88416 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_140
timestamp 1679585382
transform 1 0 89088 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_147
timestamp 1679585382
transform 1 0 89760 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_154
timestamp 1679585382
transform 1 0 90432 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_161
timestamp 1679585382
transform 1 0 91104 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_168
timestamp 1679585382
transform 1 0 91776 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_175
timestamp 1679585382
transform 1 0 92448 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_182
timestamp 1679585382
transform 1 0 93120 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_189
timestamp 1679585382
transform 1 0 93792 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_196
timestamp 1679585382
transform 1 0 94464 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_203
timestamp 1679585382
transform 1 0 95136 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_210
timestamp 1679585382
transform 1 0 95808 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_217
timestamp 1679585382
transform 1 0 96480 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_224
timestamp 1679585382
transform 1 0 97152 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_231
timestamp 1679585382
transform 1 0 97824 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_238
timestamp 1679585382
transform 1 0 98496 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_245
timestamp 1679585382
transform 1 0 99168 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_252
timestamp 1679585382
transform 1 0 99840 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_259
timestamp 1679585382
transform 1 0 100512 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_266
timestamp 1679585382
transform 1 0 101184 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_273
timestamp 1679585382
transform 1 0 101856 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_280
timestamp 1679585382
transform 1 0 102528 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_287
timestamp 1679585382
transform 1 0 103200 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_294
timestamp 1679585382
transform 1 0 103872 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_301
timestamp 1679585382
transform 1 0 104544 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_308
timestamp 1679585382
transform 1 0 105216 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_315
timestamp 1679585382
transform 1 0 105888 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_322
timestamp 1679585382
transform 1 0 106560 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_329
timestamp 1679585382
transform 1 0 107232 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_336
timestamp 1679585382
transform 1 0 107904 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_343
timestamp 1679585382
transform 1 0 108576 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_350
timestamp 1679585382
transform 1 0 109248 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_357
timestamp 1679585382
transform 1 0 109920 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_364
timestamp 1679585382
transform 1 0 110592 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_371
timestamp 1679585382
transform 1 0 111264 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_378
timestamp 1679585382
transform 1 0 111936 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_385
timestamp 1679585382
transform 1 0 112608 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_392
timestamp 1679585382
transform 1 0 113280 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_399
timestamp 1679585382
transform 1 0 113952 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_406
timestamp 1679585382
transform 1 0 114624 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_413
timestamp 1679585382
transform 1 0 115296 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_420
timestamp 1679585382
transform 1 0 115968 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_427
timestamp 1679585382
transform 1 0 116640 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_434
timestamp 1679585382
transform 1 0 117312 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_441
timestamp 1679585382
transform 1 0 117984 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_448
timestamp 1679585382
transform 1 0 118656 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_455
timestamp 1679585382
transform 1 0 119328 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_462
timestamp 1679585382
transform 1 0 120000 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_469
timestamp 1679585382
transform 1 0 120672 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_476
timestamp 1679585382
transform 1 0 121344 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_483
timestamp 1679585382
transform 1 0 122016 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_490
timestamp 1679585382
transform 1 0 122688 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_497
timestamp 1679585382
transform 1 0 123360 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_504
timestamp 1679585382
transform 1 0 124032 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_511
timestamp 1679585382
transform 1 0 124704 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_518
timestamp 1679585382
transform 1 0 125376 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_525
timestamp 1679585382
transform 1 0 126048 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_532
timestamp 1679585382
transform 1 0 126720 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_539
timestamp 1679585382
transform 1 0 127392 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_546
timestamp 1679585382
transform 1 0 128064 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_553
timestamp 1679585382
transform 1 0 128736 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_560
timestamp 1679585382
transform 1 0 129408 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_567
timestamp 1679585382
transform 1 0 130080 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_574
timestamp 1679585382
transform 1 0 130752 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_581
timestamp 1679585382
transform 1 0 131424 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_588
timestamp 1679585382
transform 1 0 132096 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_595
timestamp 1679585382
transform 1 0 132768 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_602
timestamp 1679585382
transform 1 0 133440 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_609
timestamp 1679585382
transform 1 0 134112 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_616
timestamp 1679585382
transform 1 0 134784 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_623
timestamp 1679585382
transform 1 0 135456 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_630
timestamp 1679585382
transform 1 0 136128 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_637
timestamp 1679585382
transform 1 0 136800 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_644
timestamp 1679585382
transform 1 0 137472 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_651
timestamp 1679585382
transform 1 0 138144 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_658
timestamp 1679585382
transform 1 0 138816 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_665
timestamp 1679585382
transform 1 0 139488 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_672
timestamp 1679585382
transform 1 0 140160 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_679
timestamp 1679585382
transform 1 0 140832 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_686
timestamp 1679585382
transform 1 0 141504 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_693
timestamp 1679585382
transform 1 0 142176 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_700
timestamp 1679585382
transform 1 0 142848 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_707
timestamp 1679585382
transform 1 0 143520 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_714
timestamp 1679585382
transform 1 0 144192 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_721
timestamp 1679585382
transform 1 0 144864 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_728
timestamp 1679585382
transform 1 0 145536 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_735
timestamp 1679585382
transform 1 0 146208 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_742
timestamp 1679585382
transform 1 0 146880 0 -1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_93_749
timestamp 1679585382
transform 1 0 147552 0 -1 146664
box -48 -56 720 834
use sg13g2_fill_1  FILLER_93_756
timestamp 1677583258
transform 1 0 148224 0 -1 146664
box -48 -56 144 834
use sg13g2_decap_8  FILLER_94_0
timestamp 1679585382
transform 1 0 75648 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_7
timestamp 1679585382
transform 1 0 76320 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_14
timestamp 1679585382
transform 1 0 76992 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_21
timestamp 1679585382
transform 1 0 77664 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_28
timestamp 1679585382
transform 1 0 78336 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_35
timestamp 1679585382
transform 1 0 79008 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_42
timestamp 1679585382
transform 1 0 79680 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_49
timestamp 1679585382
transform 1 0 80352 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_56
timestamp 1679585382
transform 1 0 81024 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_63
timestamp 1679585382
transform 1 0 81696 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_70
timestamp 1679585382
transform 1 0 82368 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_77
timestamp 1679585382
transform 1 0 83040 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_84
timestamp 1679585382
transform 1 0 83712 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_91
timestamp 1679585382
transform 1 0 84384 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_98
timestamp 1679585382
transform 1 0 85056 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_105
timestamp 1679585382
transform 1 0 85728 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_112
timestamp 1679585382
transform 1 0 86400 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_119
timestamp 1679585382
transform 1 0 87072 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_126
timestamp 1679585382
transform 1 0 87744 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_133
timestamp 1679585382
transform 1 0 88416 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_140
timestamp 1679585382
transform 1 0 89088 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_147
timestamp 1679585382
transform 1 0 89760 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_154
timestamp 1679585382
transform 1 0 90432 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_161
timestamp 1679585382
transform 1 0 91104 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_168
timestamp 1679585382
transform 1 0 91776 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_175
timestamp 1679585382
transform 1 0 92448 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_182
timestamp 1679585382
transform 1 0 93120 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_189
timestamp 1679585382
transform 1 0 93792 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_196
timestamp 1679585382
transform 1 0 94464 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_203
timestamp 1679585382
transform 1 0 95136 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_210
timestamp 1679585382
transform 1 0 95808 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_217
timestamp 1679585382
transform 1 0 96480 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_224
timestamp 1679585382
transform 1 0 97152 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_231
timestamp 1679585382
transform 1 0 97824 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_238
timestamp 1679585382
transform 1 0 98496 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_245
timestamp 1679585382
transform 1 0 99168 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_252
timestamp 1679585382
transform 1 0 99840 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_259
timestamp 1679585382
transform 1 0 100512 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_266
timestamp 1679585382
transform 1 0 101184 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_273
timestamp 1679585382
transform 1 0 101856 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_280
timestamp 1679585382
transform 1 0 102528 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_287
timestamp 1679585382
transform 1 0 103200 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_294
timestamp 1679585382
transform 1 0 103872 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_301
timestamp 1679585382
transform 1 0 104544 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_308
timestamp 1679585382
transform 1 0 105216 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_315
timestamp 1679585382
transform 1 0 105888 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_322
timestamp 1679585382
transform 1 0 106560 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_329
timestamp 1679585382
transform 1 0 107232 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_336
timestamp 1679585382
transform 1 0 107904 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_343
timestamp 1679585382
transform 1 0 108576 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_350
timestamp 1679585382
transform 1 0 109248 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_357
timestamp 1679585382
transform 1 0 109920 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_364
timestamp 1679585382
transform 1 0 110592 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_371
timestamp 1679585382
transform 1 0 111264 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_378
timestamp 1679585382
transform 1 0 111936 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_385
timestamp 1679585382
transform 1 0 112608 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_392
timestamp 1679585382
transform 1 0 113280 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_399
timestamp 1679585382
transform 1 0 113952 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_406
timestamp 1679585382
transform 1 0 114624 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_413
timestamp 1679585382
transform 1 0 115296 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_420
timestamp 1679585382
transform 1 0 115968 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_427
timestamp 1679585382
transform 1 0 116640 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_434
timestamp 1679585382
transform 1 0 117312 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_441
timestamp 1679585382
transform 1 0 117984 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_448
timestamp 1679585382
transform 1 0 118656 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_455
timestamp 1679585382
transform 1 0 119328 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_462
timestamp 1679585382
transform 1 0 120000 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_469
timestamp 1679585382
transform 1 0 120672 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_476
timestamp 1679585382
transform 1 0 121344 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_483
timestamp 1679585382
transform 1 0 122016 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_490
timestamp 1679585382
transform 1 0 122688 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_497
timestamp 1679585382
transform 1 0 123360 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_504
timestamp 1679585382
transform 1 0 124032 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_511
timestamp 1679585382
transform 1 0 124704 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_518
timestamp 1679585382
transform 1 0 125376 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_525
timestamp 1679585382
transform 1 0 126048 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_532
timestamp 1679585382
transform 1 0 126720 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_539
timestamp 1679585382
transform 1 0 127392 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_546
timestamp 1679585382
transform 1 0 128064 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_553
timestamp 1679585382
transform 1 0 128736 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_560
timestamp 1679585382
transform 1 0 129408 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_567
timestamp 1679585382
transform 1 0 130080 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_574
timestamp 1679585382
transform 1 0 130752 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_581
timestamp 1679585382
transform 1 0 131424 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_588
timestamp 1679585382
transform 1 0 132096 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_595
timestamp 1679585382
transform 1 0 132768 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_602
timestamp 1679585382
transform 1 0 133440 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_609
timestamp 1679585382
transform 1 0 134112 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_616
timestamp 1679585382
transform 1 0 134784 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_623
timestamp 1679585382
transform 1 0 135456 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_630
timestamp 1679585382
transform 1 0 136128 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_637
timestamp 1679585382
transform 1 0 136800 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_644
timestamp 1679585382
transform 1 0 137472 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_651
timestamp 1679585382
transform 1 0 138144 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_658
timestamp 1679585382
transform 1 0 138816 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_665
timestamp 1679585382
transform 1 0 139488 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_672
timestamp 1679585382
transform 1 0 140160 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_679
timestamp 1679585382
transform 1 0 140832 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_686
timestamp 1679585382
transform 1 0 141504 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_693
timestamp 1679585382
transform 1 0 142176 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_700
timestamp 1679585382
transform 1 0 142848 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_707
timestamp 1679585382
transform 1 0 143520 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_714
timestamp 1679585382
transform 1 0 144192 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_721
timestamp 1679585382
transform 1 0 144864 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_728
timestamp 1679585382
transform 1 0 145536 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_735
timestamp 1679585382
transform 1 0 146208 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_742
timestamp 1679585382
transform 1 0 146880 0 1 146664
box -48 -56 720 834
use sg13g2_decap_8  FILLER_94_749
timestamp 1679585382
transform 1 0 147552 0 1 146664
box -48 -56 720 834
use sg13g2_fill_1  FILLER_94_756
timestamp 1677583258
transform 1 0 148224 0 1 146664
box -48 -56 144 834
use sg13g2_decap_8  FILLER_95_0
timestamp 1679585382
transform 1 0 75648 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_7
timestamp 1679585382
transform 1 0 76320 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_14
timestamp 1679585382
transform 1 0 76992 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_21
timestamp 1679585382
transform 1 0 77664 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_28
timestamp 1679585382
transform 1 0 78336 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_35
timestamp 1679585382
transform 1 0 79008 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_42
timestamp 1679585382
transform 1 0 79680 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_49
timestamp 1679585382
transform 1 0 80352 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_56
timestamp 1679585382
transform 1 0 81024 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_63
timestamp 1679585382
transform 1 0 81696 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_70
timestamp 1679585382
transform 1 0 82368 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_77
timestamp 1679585382
transform 1 0 83040 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_84
timestamp 1679585382
transform 1 0 83712 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_91
timestamp 1679585382
transform 1 0 84384 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_98
timestamp 1679585382
transform 1 0 85056 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_105
timestamp 1679585382
transform 1 0 85728 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_112
timestamp 1679585382
transform 1 0 86400 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_119
timestamp 1679585382
transform 1 0 87072 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_126
timestamp 1679585382
transform 1 0 87744 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_133
timestamp 1679585382
transform 1 0 88416 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_140
timestamp 1679585382
transform 1 0 89088 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_147
timestamp 1679585382
transform 1 0 89760 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_154
timestamp 1679585382
transform 1 0 90432 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_161
timestamp 1679585382
transform 1 0 91104 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_168
timestamp 1679585382
transform 1 0 91776 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_175
timestamp 1679585382
transform 1 0 92448 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_182
timestamp 1679585382
transform 1 0 93120 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_189
timestamp 1679585382
transform 1 0 93792 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_196
timestamp 1679585382
transform 1 0 94464 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_203
timestamp 1679585382
transform 1 0 95136 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_210
timestamp 1679585382
transform 1 0 95808 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_217
timestamp 1679585382
transform 1 0 96480 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_224
timestamp 1679585382
transform 1 0 97152 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_231
timestamp 1679585382
transform 1 0 97824 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_238
timestamp 1679585382
transform 1 0 98496 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_245
timestamp 1679585382
transform 1 0 99168 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_252
timestamp 1679585382
transform 1 0 99840 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_259
timestamp 1679585382
transform 1 0 100512 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_266
timestamp 1679585382
transform 1 0 101184 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_273
timestamp 1679585382
transform 1 0 101856 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_280
timestamp 1679585382
transform 1 0 102528 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_287
timestamp 1679585382
transform 1 0 103200 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_294
timestamp 1679585382
transform 1 0 103872 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_301
timestamp 1679585382
transform 1 0 104544 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_308
timestamp 1679585382
transform 1 0 105216 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_315
timestamp 1679585382
transform 1 0 105888 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_322
timestamp 1679585382
transform 1 0 106560 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_329
timestamp 1679585382
transform 1 0 107232 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_336
timestamp 1679585382
transform 1 0 107904 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_343
timestamp 1679585382
transform 1 0 108576 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_350
timestamp 1679585382
transform 1 0 109248 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_357
timestamp 1679585382
transform 1 0 109920 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_364
timestamp 1679585382
transform 1 0 110592 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_371
timestamp 1679585382
transform 1 0 111264 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_378
timestamp 1679585382
transform 1 0 111936 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_385
timestamp 1679585382
transform 1 0 112608 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_392
timestamp 1679585382
transform 1 0 113280 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_399
timestamp 1679585382
transform 1 0 113952 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_406
timestamp 1679585382
transform 1 0 114624 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_413
timestamp 1679585382
transform 1 0 115296 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_420
timestamp 1679585382
transform 1 0 115968 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_427
timestamp 1679585382
transform 1 0 116640 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_434
timestamp 1679585382
transform 1 0 117312 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_441
timestamp 1679585382
transform 1 0 117984 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_448
timestamp 1679585382
transform 1 0 118656 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_455
timestamp 1679585382
transform 1 0 119328 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_462
timestamp 1679585382
transform 1 0 120000 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_469
timestamp 1679585382
transform 1 0 120672 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_476
timestamp 1679585382
transform 1 0 121344 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_483
timestamp 1679585382
transform 1 0 122016 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_490
timestamp 1679585382
transform 1 0 122688 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_497
timestamp 1679585382
transform 1 0 123360 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_504
timestamp 1679585382
transform 1 0 124032 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_511
timestamp 1679585382
transform 1 0 124704 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_518
timestamp 1679585382
transform 1 0 125376 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_525
timestamp 1679585382
transform 1 0 126048 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_532
timestamp 1679585382
transform 1 0 126720 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_539
timestamp 1679585382
transform 1 0 127392 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_546
timestamp 1679585382
transform 1 0 128064 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_553
timestamp 1679585382
transform 1 0 128736 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_560
timestamp 1679585382
transform 1 0 129408 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_567
timestamp 1679585382
transform 1 0 130080 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_574
timestamp 1679585382
transform 1 0 130752 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_581
timestamp 1679585382
transform 1 0 131424 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_588
timestamp 1679585382
transform 1 0 132096 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_595
timestamp 1679585382
transform 1 0 132768 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_602
timestamp 1679585382
transform 1 0 133440 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_609
timestamp 1679585382
transform 1 0 134112 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_616
timestamp 1679585382
transform 1 0 134784 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_623
timestamp 1679585382
transform 1 0 135456 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_630
timestamp 1679585382
transform 1 0 136128 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_637
timestamp 1679585382
transform 1 0 136800 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_644
timestamp 1679585382
transform 1 0 137472 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_651
timestamp 1679585382
transform 1 0 138144 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_658
timestamp 1679585382
transform 1 0 138816 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_665
timestamp 1679585382
transform 1 0 139488 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_672
timestamp 1679585382
transform 1 0 140160 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_679
timestamp 1679585382
transform 1 0 140832 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_686
timestamp 1679585382
transform 1 0 141504 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_693
timestamp 1679585382
transform 1 0 142176 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_700
timestamp 1679585382
transform 1 0 142848 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_707
timestamp 1679585382
transform 1 0 143520 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_714
timestamp 1679585382
transform 1 0 144192 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_721
timestamp 1679585382
transform 1 0 144864 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_728
timestamp 1679585382
transform 1 0 145536 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_735
timestamp 1679585382
transform 1 0 146208 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_742
timestamp 1679585382
transform 1 0 146880 0 -1 148176
box -48 -56 720 834
use sg13g2_decap_8  FILLER_95_749
timestamp 1679585382
transform 1 0 147552 0 -1 148176
box -48 -56 720 834
use sg13g2_fill_1  FILLER_95_756
timestamp 1677583258
transform 1 0 148224 0 -1 148176
box -48 -56 144 834
use sg13g2_dlygate4sd3_1  hold11
timestamp 1677675658
transform 1 0 103584 0 1 95256
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold12
timestamp 1677675658
transform 1 0 119424 0 1 128520
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold13
timestamp 1677675658
transform 1 0 120288 0 1 128520
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold14
timestamp 1677675658
transform 1 0 78528 0 -1 133056
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold15
timestamp 1677675658
transform 1 0 96096 0 -1 130032
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold16
timestamp 1677675658
transform 1 0 98304 0 1 131544
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold17
timestamp 1677675658
transform -1 0 98976 0 1 133056
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold18
timestamp 1677675658
transform -1 0 111552 0 -1 131544
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold19
timestamp 1677675658
transform -1 0 110592 0 -1 131544
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold20
timestamp 1677675658
transform -1 0 121056 0 -1 133056
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold21
timestamp 1677675658
transform -1 0 120192 0 -1 133056
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold22
timestamp 1677675658
transform -1 0 122304 0 -1 125496
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold23
timestamp 1677675658
transform -1 0 115200 0 1 133056
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold24
timestamp 1677675658
transform 1 0 112704 0 1 131544
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold25
timestamp 1677675658
transform -1 0 105504 0 1 130032
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold26
timestamp 1677675658
transform -1 0 103296 0 -1 131544
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold27
timestamp 1677675658
transform 1 0 103296 0 -1 131544
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold28
timestamp 1677675658
transform 1 0 78816 0 1 123984
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold29
timestamp 1677675658
transform 1 0 96000 0 1 128520
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold30
timestamp 1677675658
transform 1 0 99840 0 -1 131544
box -48 -56 912 834
use sg13g2_dlygate4sd3_1  hold31
timestamp 1677675658
transform 1 0 102912 0 -1 133056
box -48 -56 912 834
use sg13g2_IOPadIn  inputs\[0\].input_pad
timestamp 1716382777
transform 0 1 28000 1 0 144000
box -124 0 16124 36000
use sg13g2_IOPadIn  inputs\[1\].input_pad
timestamp 1716382777
transform 0 1 28000 1 0 128000
box -124 0 16124 36000
use sg13g2_IOPadIn  inputs\[2\].input_pad
timestamp 1716382777
transform 0 1 28000 1 0 112000
box -124 0 16124 36000
use sg13g2_IOPadIn  inputs\[3\].input_pad
timestamp 1716382777
transform 0 1 28000 1 0 96000
box -124 0 16124 36000
use sg13g2_IOPadIn  inputs\[4\].input_pad
timestamp 1716382777
transform 0 1 28000 1 0 80000
box -124 0 16124 36000
use sg13g2_IOPadIn  inputs\[5\].input_pad
timestamp 1716382777
transform 0 1 28000 1 0 64000
box -124 0 16124 36000
use sg13g2_IOPadIn  inputs\[6\].input_pad
timestamp 1716382777
transform 1 0 112000 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadIn  inputs\[7\].input_pad
timestamp 1716382777
transform 1 0 96000 0 1 28000
box -124 0 16124 36000
use bondpad_70x70_novias  IO_BOND_clk_pad
timestamp 1590364920
transform 1 0 65000 0 1 14000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_inputs\[0\].input_pad
timestamp 1590364920
transform 0 1 14000 1 0 145000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_inputs\[1\].input_pad
timestamp 1590364920
transform 0 1 14000 1 0 129000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_inputs\[2\].input_pad
timestamp 1590364920
transform 0 1 14000 1 0 113000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_inputs\[3\].input_pad
timestamp 1590364920
transform 0 1 14000 1 0 97000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_inputs\[4\].input_pad
timestamp 1590364920
transform 0 1 14000 1 0 81000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_inputs\[5\].input_pad
timestamp 1590364920
transform 0 1 14000 1 0 65000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_inputs\[6\].input_pad
timestamp 1590364920
transform 1 0 113000 0 1 14000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_inputs\[7\].input_pad
timestamp 1590364920
transform 1 0 97000 0 1 14000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_iovdd_pads\[0\].iovdd_pad
timestamp 1590364920
transform 1 0 81000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_iovss_pads\[0\].iovss_pad
timestamp 1590364920
transform 1 0 65000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_outputs\[0\].output_pad
timestamp 1590364920
transform 1 0 145000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_outputs\[1\].output_pad
timestamp 1590364920
transform 1 0 129000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_outputs\[2\].output_pad
timestamp 1590364920
transform 1 0 113000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_outputs\[3\].output_pad
timestamp 1590364920
transform 1 0 97000 0 -1 210000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_outputs\[4\].output_pad
timestamp 1590364920
transform 0 -1 210000 1 0 145000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_outputs\[5\].output_pad
timestamp 1590364920
transform 0 -1 210000 1 0 129000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_outputs\[6\].output_pad
timestamp 1590364920
transform 0 -1 210000 1 0 113000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_outputs\[7\].output_pad
timestamp 1590364920
transform 0 -1 210000 1 0 97000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_outputs\[8\].output_pad
timestamp 1590364920
transform 0 -1 210000 1 0 81000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_outputs\[9\].output_pad
timestamp 1590364920
transform 0 -1 210000 1 0 65000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_rst_n_pad
timestamp 1590364920
transform 1 0 81000 0 1 14000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_vdd_pads\[0\].vdd_pad
timestamp 1590364920
transform 1 0 129000 0 1 14000
box 0 0 14000 14000
use bondpad_70x70_novias  IO_BOND_vss_pads\[0\].vss_pad
timestamp 1590364920
transform 1 0 145000 0 1 14000
box 0 0 14000 14000
use sg13g2_Corner  IO_CORNER_NORTH_EAST_INST
timestamp 1716382778
transform -1 0 196000 0 -1 196000
box 1076 1076 36124 36124
use sg13g2_Corner  IO_CORNER_NORTH_WEST_INST
timestamp 1716382778
transform 1 0 28000 0 -1 196000
box 1076 1076 36124 36124
use sg13g2_Corner  IO_CORNER_SOUTH_EAST_INST
timestamp 1716382778
transform -1 0 196000 0 1 28000
box 1076 1076 36124 36124
use sg13g2_Corner  IO_CORNER_SOUTH_WEST_INST
timestamp 1716382778
transform 1 0 28000 0 1 28000
box 1076 1076 36124 36124
use sg13g2_IOPadIOVdd  iovdd_pads\[0\].iovdd_pad
timestamp 1716382778
transform 1 0 80000 0 -1 196000
box -124 0 16124 35600
use sg13g2_IOPadIOVss  iovss_pads\[0\].iovss_pad
timestamp 1716382777
transform 1 0 64000 0 -1 196000
box -124 0 16124 35600
use sg13g2_IOPadOut30mA  outputs\[0\].output_pad
timestamp 1716382777
transform 1 0 144000 0 -1 196000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  outputs\[1\].output_pad
timestamp 1716382777
transform 1 0 128000 0 -1 196000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  outputs\[2\].output_pad
timestamp 1716382777
transform 1 0 112000 0 -1 196000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  outputs\[3\].output_pad
timestamp 1716382777
transform 1 0 96000 0 -1 196000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  outputs\[4\].output_pad
timestamp 1716382777
transform 0 -1 196000 1 0 144000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  outputs\[5\].output_pad
timestamp 1716382777
transform 0 -1 196000 1 0 128000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  outputs\[6\].output_pad
timestamp 1716382777
transform 0 -1 196000 1 0 112000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  outputs\[7\].output_pad
timestamp 1716382777
transform 0 -1 196000 1 0 96000
box -124 0 16124 36000
use sg13g2_tielo  outputs\[8\].output_pad_1
timestamp 1680007837
transform 1 0 147936 0 1 87696
box -48 -56 432 834
use sg13g2_IOPadOut30mA  outputs\[8\].output_pad
timestamp 1716382777
transform 0 -1 196000 1 0 80000
box -124 0 16124 36000
use sg13g2_IOPadOut30mA  outputs\[9\].output_pad
timestamp 1716382777
transform 0 -1 196000 1 0 64000
box -124 0 16124 36000
use sg13g2_tielo  outputs\[9\].output_pad_2
timestamp 1680007837
transform 1 0 147936 0 1 75600
box -48 -56 432 834
use sg13g2_IOPadIn  rst_n_pad
timestamp 1716382777
transform 1 0 80000 0 1 28000
box -124 0 16124 36000
use sg13g2_IOPadVdd  vdd_pads\[0\].vdd_pad
timestamp 1716382777
transform 1 0 128000 0 1 28000
box -124 0 16124 35600
use sg13g2_IOPadVss  vss_pads\[0\].vss_pad
timestamp 1716382777
transform 1 0 144000 0 1 28000
box -124 0 16124 35600
<< labels >>
flabel metal7 s 81000 196000 95000 210000 0 FreeSans 102400 0 0 0 IOVDD
port 0 nsew power input
flabel metal7 s 65000 196000 79000 210000 0 FreeSans 102400 0 0 0 IOVSS
port 1 nsew ground input
flabel metal7 s 129000 14000 143000 28000 0 FreeSans 102400 0 0 0 VDD
port 2 nsew power input
flabel metal7 s 145000 14000 159000 28000 0 FreeSans 102400 0 0 0 VSS
port 3 nsew ground input
flabel metal7 s 65000 14000 79000 28000 0 FreeSans 102400 0 0 0 clk_PAD
port 4 nsew signal bidirectional
flabel metal7 s 14000 145000 28000 159000 0 FreeSans 102400 0 0 0 input_PAD[0]
port 5 nsew signal bidirectional
flabel metal7 s 14000 129000 28000 143000 0 FreeSans 102400 0 0 0 input_PAD[1]
port 6 nsew signal bidirectional
flabel metal7 s 14000 113000 28000 127000 0 FreeSans 102400 0 0 0 input_PAD[2]
port 7 nsew signal bidirectional
flabel metal7 s 14000 97000 28000 111000 0 FreeSans 102400 0 0 0 input_PAD[3]
port 8 nsew signal bidirectional
flabel metal7 s 14000 81000 28000 95000 0 FreeSans 102400 0 0 0 input_PAD[4]
port 9 nsew signal bidirectional
flabel metal7 s 14000 65000 28000 79000 0 FreeSans 102400 0 0 0 input_PAD[5]
port 10 nsew signal bidirectional
flabel metal7 s 113000 14000 127000 28000 0 FreeSans 102400 0 0 0 input_PAD[6]
port 11 nsew signal bidirectional
flabel metal7 s 97000 14000 111000 28000 0 FreeSans 102400 0 0 0 input_PAD[7]
port 12 nsew signal bidirectional
flabel metal7 s 145000 196000 159000 210000 0 FreeSans 102400 0 0 0 output_PAD[0]
port 13 nsew signal bidirectional
flabel metal7 s 129000 196000 143000 210000 0 FreeSans 102400 0 0 0 output_PAD[1]
port 14 nsew signal bidirectional
flabel metal7 s 113000 196000 127000 210000 0 FreeSans 102400 0 0 0 output_PAD[2]
port 15 nsew signal bidirectional
flabel metal7 s 97000 196000 111000 210000 0 FreeSans 102400 0 0 0 output_PAD[3]
port 16 nsew signal bidirectional
flabel metal7 s 196000 145000 210000 159000 0 FreeSans 102400 0 0 0 output_PAD[4]
port 17 nsew signal bidirectional
flabel metal7 s 196000 129000 210000 143000 0 FreeSans 102400 0 0 0 output_PAD[5]
port 18 nsew signal bidirectional
flabel metal7 s 196000 113000 210000 127000 0 FreeSans 102400 0 0 0 output_PAD[6]
port 19 nsew signal bidirectional
flabel metal7 s 196000 97000 210000 111000 0 FreeSans 102400 0 0 0 output_PAD[7]
port 20 nsew signal bidirectional
flabel metal7 s 196000 81000 210000 95000 0 FreeSans 102400 0 0 0 output_PAD[8]
port 21 nsew signal bidirectional
flabel metal7 s 196000 65000 210000 79000 0 FreeSans 102400 0 0 0 output_PAD[9]
port 22 nsew signal bidirectional
flabel metal7 s 81000 14000 95000 28000 0 FreeSans 102400 0 0 0 rst_n_PAD
port 23 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 224000 224000
<< end >>
