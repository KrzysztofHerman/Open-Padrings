module FMD_QNC_Padframe28 (\IO_CORNER_NORTH_WEST_INST.iovdd_RING ,
    \IO_CORNER_NORTH_WEST_INST.iovss_RING ,
    \IO_CORNER_NORTH_WEST_INST.vdd_RING ,
    \IO_CORNER_NORTH_WEST_INST.vss_RING ,
    VSS,
    VDD,
    ui_PAD,
    uo_PAD);
 inout \IO_CORNER_NORTH_WEST_INST.iovdd_RING ;
 inout \IO_CORNER_NORTH_WEST_INST.iovss_RING ;
 inout \IO_CORNER_NORTH_WEST_INST.vdd_RING ;
 inout \IO_CORNER_NORTH_WEST_INST.vss_RING ;
 inout VSS;
 inout VDD;
 inout [11:0] ui_PAD;
 inout [11:0] uo_PAD;

 wire \ui_PAD2CORE[0] ;
 wire \ui_PAD2CORE[10] ;
 wire \ui_PAD2CORE[11] ;
 wire \ui_PAD2CORE[1] ;
 wire \ui_PAD2CORE[2] ;
 wire \ui_PAD2CORE[3] ;
 wire \ui_PAD2CORE[4] ;
 wire \ui_PAD2CORE[5] ;
 wire \ui_PAD2CORE[6] ;
 wire \ui_PAD2CORE[7] ;
 wire \ui_PAD2CORE[8] ;
 wire \ui_PAD2CORE[9] ;
 wire IOVDD;
 wire IOVSS;

 sg13g2_IOPadIOVdd sg13g2_IOPadIOVdd_north (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIOVss sg13g2_IOPadIOVss_north (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[0].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[0] ),
    .pad(ui_PAD[0]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[10].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[10] ),
    .pad(ui_PAD[10]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[11].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[11] ),
    .pad(ui_PAD[11]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[1].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[1] ),
    .pad(ui_PAD[1]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[2].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[2] ),
    .pad(ui_PAD[2]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[3].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[3] ),
    .pad(ui_PAD[3]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[4].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[4] ),
    .pad(ui_PAD[4]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[5].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[5] ),
    .pad(ui_PAD[5]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[6].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[6] ),
    .pad(ui_PAD[6]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[7].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[7] ),
    .pad(ui_PAD[7]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[8].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[8] ),
    .pad(ui_PAD[8]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[9].ui  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\ui_PAD2CORE[9] ),
    .pad(ui_PAD[9]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[0].uo  (.c2p(\ui_PAD2CORE[0] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[0]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[10].uo  (.c2p(\ui_PAD2CORE[10] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[10]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[11].uo  (.c2p(\ui_PAD2CORE[11] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[11]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[1].uo  (.c2p(\ui_PAD2CORE[1] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[1]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[2].uo  (.c2p(\ui_PAD2CORE[2] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[2]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[3].uo  (.c2p(\ui_PAD2CORE[3] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[3]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[4].uo  (.c2p(\ui_PAD2CORE[4] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[4]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[5].uo  (.c2p(\ui_PAD2CORE[5] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[5]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[6].uo  (.c2p(\ui_PAD2CORE[6] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[6]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[7].uo  (.c2p(\ui_PAD2CORE[7] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[7]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[8].uo  (.c2p(\ui_PAD2CORE[8] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[8]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[9].uo  (.c2p(\ui_PAD2CORE[9] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(uo_PAD[9]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadVdd sg13g2_IOPadVdd_south (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadVss sg13g2_IOPadVss_south (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_Corner IO_CORNER_NORTH_WEST_INST (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_Corner IO_CORNER_NORTH_EAST_INST (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_Corner IO_CORNER_SOUTH_WEST_INST (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_Corner IO_CORNER_SOUTH_EAST_INST (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 bondpad_70x70 IO_BOND_sg13g2_IOPadIOVdd_north (.pad(\IO_CORNER_NORTH_WEST_INST.iovdd_RING ));
 bondpad_70x70 IO_BOND_sg13g2_IOPadIOVss_north (.pad(\IO_CORNER_NORTH_WEST_INST.iovss_RING ));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[0].ui  (.pad(ui_PAD[0]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[10].ui  (.pad(ui_PAD[10]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[11].ui  (.pad(ui_PAD[11]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[1].ui  (.pad(ui_PAD[1]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[2].ui  (.pad(ui_PAD[2]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[3].ui  (.pad(ui_PAD[3]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[4].ui  (.pad(ui_PAD[4]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[5].ui  (.pad(ui_PAD[5]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[6].ui  (.pad(ui_PAD[6]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[7].ui  (.pad(ui_PAD[7]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[8].ui  (.pad(ui_PAD[8]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[9].ui  (.pad(ui_PAD[9]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[0].uo  (.pad(uo_PAD[0]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[10].uo  (.pad(uo_PAD[10]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[11].uo  (.pad(uo_PAD[11]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[1].uo  (.pad(uo_PAD[1]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[2].uo  (.pad(uo_PAD[2]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[3].uo  (.pad(uo_PAD[3]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[4].uo  (.pad(uo_PAD[4]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[5].uo  (.pad(uo_PAD[5]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[6].uo  (.pad(uo_PAD[6]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[7].uo  (.pad(uo_PAD[7]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[8].uo  (.pad(uo_PAD[8]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[9].uo  (.pad(uo_PAD[9]));
 bondpad_70x70 IO_BOND_sg13g2_IOPadVdd_south (.pad(\IO_CORNER_NORTH_WEST_INST.vdd_RING ));
 bondpad_70x70 IO_BOND_sg13g2_IOPadVss_south (.pad(\IO_CORNER_NORTH_WEST_INST.vss_RING ));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_96_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_97_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_98_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_99_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_100_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_101_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_102_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_103_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_104_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_105_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_106_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_107_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_108_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_109_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_110_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_111_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_112_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_113_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_114_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_115_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_116_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_117_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_118_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_119_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_120_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_121_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_122_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_123_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_124_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_125_1001 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_763 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_770 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_777 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_784 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_791 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_798 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_805 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_812 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_819 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_826 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_833 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_840 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_847 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_854 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_861 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_868 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_875 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_882 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_889 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_896 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_903 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_910 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_917 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_924 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_931 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_938 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_945 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_952 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_959 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_966 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_973 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_980 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_987 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_994 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_126_1001 (.VDD(VDD),
    .VSS(VSS));
endmodule
