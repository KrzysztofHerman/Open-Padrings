module FMD_QNC_Padframe24 (ui_PAD,
    uo_PAD);
 inout [9:0] ui_PAD;
 inout [9:0] uo_PAD;

 wire \ui_PAD2CORE[0] ;
 wire \ui_PAD2CORE[1] ;
 wire \ui_PAD2CORE[2] ;
 wire \ui_PAD2CORE[3] ;
 wire \ui_PAD2CORE[4] ;
 wire \ui_PAD2CORE[5] ;
 wire \ui_PAD2CORE[6] ;
 wire \ui_PAD2CORE[7] ;
 wire \ui_PAD2CORE[8] ;
 wire \ui_PAD2CORE[9] ;

 sg13g2_IOPadIOVdd sg13g2_IOPadIOVdd_north ();
 sg13g2_IOPadIOVss sg13g2_IOPadIOVss_north ();
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[0].ui  (.p2c(\ui_PAD2CORE[0] ),
    .pad(ui_PAD[0]));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[1].ui  (.p2c(\ui_PAD2CORE[1] ),
    .pad(ui_PAD[1]));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[2].ui  (.p2c(\ui_PAD2CORE[2] ),
    .pad(ui_PAD[2]));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[3].ui  (.p2c(\ui_PAD2CORE[3] ),
    .pad(ui_PAD[3]));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[4].ui  (.p2c(\ui_PAD2CORE[4] ),
    .pad(ui_PAD[4]));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[5].ui  (.p2c(\ui_PAD2CORE[5] ),
    .pad(ui_PAD[5]));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[6].ui  (.p2c(\ui_PAD2CORE[6] ),
    .pad(ui_PAD[6]));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[7].ui  (.p2c(\ui_PAD2CORE[7] ),
    .pad(ui_PAD[7]));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[8].ui  (.p2c(\ui_PAD2CORE[8] ),
    .pad(ui_PAD[8]));
 sg13g2_IOPadIn \sg13g2_IOPadIn_ui[9].ui  (.p2c(\ui_PAD2CORE[9] ),
    .pad(ui_PAD[9]));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[0].uo  (.c2p(\ui_PAD2CORE[0] ),
    .pad(uo_PAD[0]));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[1].uo  (.c2p(\ui_PAD2CORE[1] ),
    .pad(uo_PAD[1]));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[2].uo  (.c2p(\ui_PAD2CORE[2] ),
    .pad(uo_PAD[2]));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[3].uo  (.c2p(\ui_PAD2CORE[3] ),
    .pad(uo_PAD[3]));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[4].uo  (.c2p(\ui_PAD2CORE[4] ),
    .pad(uo_PAD[4]));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[5].uo  (.c2p(\ui_PAD2CORE[5] ),
    .pad(uo_PAD[5]));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[6].uo  (.c2p(\ui_PAD2CORE[6] ),
    .pad(uo_PAD[6]));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[7].uo  (.c2p(\ui_PAD2CORE[7] ),
    .pad(uo_PAD[7]));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[8].uo  (.c2p(\ui_PAD2CORE[8] ),
    .pad(uo_PAD[8]));
 sg13g2_IOPadOut30mA \sg13g2_IOPadOut30mA_uo[9].uo  (.c2p(\ui_PAD2CORE[9] ),
    .pad(uo_PAD[9]));
 sg13g2_IOPadVdd sg13g2_IOPadVdd_south ();
 sg13g2_IOPadVss sg13g2_IOPadVss_south ();
 sg13g2_Corner IO_CORNER_NORTH_WEST_INST ();
 sg13g2_Corner IO_CORNER_NORTH_EAST_INST ();
 sg13g2_Corner IO_CORNER_SOUTH_WEST_INST ();
 sg13g2_Corner IO_CORNER_SOUTH_EAST_INST ();
 bondpad_70x70 IO_BOND_sg13g2_IOPadIOVdd_north (.pad(\IO_CORNER_NORTH_WEST_INST.iovdd_RING ));
 bondpad_70x70 IO_BOND_sg13g2_IOPadIOVss_north (.pad(\IO_CORNER_NORTH_WEST_INST.iovss_RING ));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[0].ui  (.pad(ui_PAD[0]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[1].ui  (.pad(ui_PAD[1]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[2].ui  (.pad(ui_PAD[2]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[3].ui  (.pad(ui_PAD[3]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[4].ui  (.pad(ui_PAD[4]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[5].ui  (.pad(ui_PAD[5]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[6].ui  (.pad(ui_PAD[6]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[7].ui  (.pad(ui_PAD[7]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[8].ui  (.pad(ui_PAD[8]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadIn_ui[9].ui  (.pad(ui_PAD[9]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[0].uo  (.pad(uo_PAD[0]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[1].uo  (.pad(uo_PAD[1]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[2].uo  (.pad(uo_PAD[2]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[3].uo  (.pad(uo_PAD[3]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[4].uo  (.pad(uo_PAD[4]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[5].uo  (.pad(uo_PAD[5]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[6].uo  (.pad(uo_PAD[6]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[7].uo  (.pad(uo_PAD[7]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[8].uo  (.pad(uo_PAD[8]));
 bondpad_70x70 \IO_BOND_sg13g2_IOPadOut30mA_uo[9].uo  (.pad(uo_PAD[9]));
 bondpad_70x70 IO_BOND_sg13g2_IOPadVdd_south (.pad(\IO_CORNER_NORTH_WEST_INST.vdd_RING ));
 bondpad_70x70 IO_BOND_sg13g2_IOPadVss_south (.pad(\IO_CORNER_NORTH_WEST_INST.vss_RING ));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_fill_1 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_fill_1 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_fill_1 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_fill_1 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_fill_1 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_fill_1 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_fill_1 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_fill_1 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_fill_1 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_fill_1 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_fill_1 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_fill_1 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_fill_1 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_fill_1 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_fill_1 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_fill_1 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_fill_1 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_fill_1 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_fill_1 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_fill_1 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_fill_1 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_fill_1 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_decap_8 FILLER_22_406 ();
 sg13g2_decap_8 FILLER_22_413 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_decap_8 FILLER_22_427 ();
 sg13g2_decap_8 FILLER_22_434 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_8 FILLER_22_483 ();
 sg13g2_decap_8 FILLER_22_490 ();
 sg13g2_decap_8 FILLER_22_497 ();
 sg13g2_decap_8 FILLER_22_504 ();
 sg13g2_decap_8 FILLER_22_511 ();
 sg13g2_decap_8 FILLER_22_518 ();
 sg13g2_decap_8 FILLER_22_525 ();
 sg13g2_decap_8 FILLER_22_532 ();
 sg13g2_decap_8 FILLER_22_539 ();
 sg13g2_decap_8 FILLER_22_546 ();
 sg13g2_decap_8 FILLER_22_553 ();
 sg13g2_decap_8 FILLER_22_560 ();
 sg13g2_decap_8 FILLER_22_567 ();
 sg13g2_decap_8 FILLER_22_574 ();
 sg13g2_decap_8 FILLER_22_581 ();
 sg13g2_decap_8 FILLER_22_588 ();
 sg13g2_decap_8 FILLER_22_595 ();
 sg13g2_decap_8 FILLER_22_602 ();
 sg13g2_decap_8 FILLER_22_609 ();
 sg13g2_decap_8 FILLER_22_616 ();
 sg13g2_decap_8 FILLER_22_623 ();
 sg13g2_decap_8 FILLER_22_630 ();
 sg13g2_decap_8 FILLER_22_637 ();
 sg13g2_decap_8 FILLER_22_644 ();
 sg13g2_decap_8 FILLER_22_651 ();
 sg13g2_decap_8 FILLER_22_658 ();
 sg13g2_decap_8 FILLER_22_665 ();
 sg13g2_decap_8 FILLER_22_672 ();
 sg13g2_decap_8 FILLER_22_679 ();
 sg13g2_decap_8 FILLER_22_686 ();
 sg13g2_decap_8 FILLER_22_693 ();
 sg13g2_decap_8 FILLER_22_700 ();
 sg13g2_decap_8 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_714 ();
 sg13g2_decap_8 FILLER_22_721 ();
 sg13g2_decap_8 FILLER_22_728 ();
 sg13g2_decap_8 FILLER_22_735 ();
 sg13g2_decap_8 FILLER_22_742 ();
 sg13g2_decap_8 FILLER_22_749 ();
 sg13g2_decap_8 FILLER_22_756 ();
 sg13g2_decap_8 FILLER_22_763 ();
 sg13g2_decap_8 FILLER_22_770 ();
 sg13g2_decap_8 FILLER_22_777 ();
 sg13g2_decap_8 FILLER_22_784 ();
 sg13g2_decap_8 FILLER_22_791 ();
 sg13g2_decap_8 FILLER_22_798 ();
 sg13g2_decap_8 FILLER_22_805 ();
 sg13g2_decap_8 FILLER_22_812 ();
 sg13g2_decap_8 FILLER_22_819 ();
 sg13g2_decap_8 FILLER_22_826 ();
 sg13g2_decap_8 FILLER_22_833 ();
 sg13g2_fill_1 FILLER_22_840 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_fill_1 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_301 ();
 sg13g2_decap_8 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_decap_8 FILLER_24_322 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_8 FILLER_24_357 ();
 sg13g2_decap_8 FILLER_24_364 ();
 sg13g2_decap_8 FILLER_24_371 ();
 sg13g2_decap_8 FILLER_24_378 ();
 sg13g2_decap_8 FILLER_24_385 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_decap_8 FILLER_24_406 ();
 sg13g2_decap_8 FILLER_24_413 ();
 sg13g2_decap_8 FILLER_24_420 ();
 sg13g2_decap_8 FILLER_24_427 ();
 sg13g2_decap_8 FILLER_24_434 ();
 sg13g2_decap_8 FILLER_24_441 ();
 sg13g2_decap_8 FILLER_24_448 ();
 sg13g2_decap_8 FILLER_24_455 ();
 sg13g2_decap_8 FILLER_24_462 ();
 sg13g2_decap_8 FILLER_24_469 ();
 sg13g2_decap_8 FILLER_24_476 ();
 sg13g2_decap_8 FILLER_24_483 ();
 sg13g2_decap_8 FILLER_24_490 ();
 sg13g2_decap_8 FILLER_24_497 ();
 sg13g2_decap_8 FILLER_24_504 ();
 sg13g2_decap_8 FILLER_24_511 ();
 sg13g2_decap_8 FILLER_24_518 ();
 sg13g2_decap_8 FILLER_24_525 ();
 sg13g2_decap_8 FILLER_24_532 ();
 sg13g2_decap_8 FILLER_24_539 ();
 sg13g2_decap_8 FILLER_24_546 ();
 sg13g2_decap_8 FILLER_24_553 ();
 sg13g2_decap_8 FILLER_24_560 ();
 sg13g2_decap_8 FILLER_24_567 ();
 sg13g2_decap_8 FILLER_24_574 ();
 sg13g2_decap_8 FILLER_24_581 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_8 FILLER_24_595 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_8 FILLER_24_609 ();
 sg13g2_decap_8 FILLER_24_616 ();
 sg13g2_decap_8 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_630 ();
 sg13g2_decap_8 FILLER_24_637 ();
 sg13g2_decap_8 FILLER_24_644 ();
 sg13g2_decap_8 FILLER_24_651 ();
 sg13g2_decap_8 FILLER_24_658 ();
 sg13g2_decap_8 FILLER_24_665 ();
 sg13g2_decap_8 FILLER_24_672 ();
 sg13g2_decap_8 FILLER_24_679 ();
 sg13g2_decap_8 FILLER_24_686 ();
 sg13g2_decap_8 FILLER_24_693 ();
 sg13g2_decap_8 FILLER_24_700 ();
 sg13g2_decap_8 FILLER_24_707 ();
 sg13g2_decap_8 FILLER_24_714 ();
 sg13g2_decap_8 FILLER_24_721 ();
 sg13g2_decap_8 FILLER_24_728 ();
 sg13g2_decap_8 FILLER_24_735 ();
 sg13g2_decap_8 FILLER_24_742 ();
 sg13g2_decap_8 FILLER_24_749 ();
 sg13g2_decap_8 FILLER_24_756 ();
 sg13g2_decap_8 FILLER_24_763 ();
 sg13g2_decap_8 FILLER_24_770 ();
 sg13g2_decap_8 FILLER_24_777 ();
 sg13g2_decap_8 FILLER_24_784 ();
 sg13g2_decap_8 FILLER_24_791 ();
 sg13g2_decap_8 FILLER_24_798 ();
 sg13g2_decap_8 FILLER_24_805 ();
 sg13g2_decap_8 FILLER_24_812 ();
 sg13g2_decap_8 FILLER_24_819 ();
 sg13g2_decap_8 FILLER_24_826 ();
 sg13g2_decap_8 FILLER_24_833 ();
 sg13g2_fill_1 FILLER_24_840 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_532 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_8 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_decap_8 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_581 ();
 sg13g2_decap_8 FILLER_25_588 ();
 sg13g2_decap_8 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_fill_1 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_decap_8 FILLER_26_462 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_8 FILLER_26_532 ();
 sg13g2_decap_8 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_651 ();
 sg13g2_decap_8 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_8 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_777 ();
 sg13g2_decap_8 FILLER_26_784 ();
 sg13g2_decap_8 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_fill_1 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_fill_1 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_decap_8 FILLER_28_427 ();
 sg13g2_decap_8 FILLER_28_434 ();
 sg13g2_decap_8 FILLER_28_441 ();
 sg13g2_decap_8 FILLER_28_448 ();
 sg13g2_decap_8 FILLER_28_455 ();
 sg13g2_decap_8 FILLER_28_462 ();
 sg13g2_decap_8 FILLER_28_469 ();
 sg13g2_decap_8 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_483 ();
 sg13g2_decap_8 FILLER_28_490 ();
 sg13g2_decap_8 FILLER_28_497 ();
 sg13g2_decap_8 FILLER_28_504 ();
 sg13g2_decap_8 FILLER_28_511 ();
 sg13g2_decap_8 FILLER_28_518 ();
 sg13g2_decap_8 FILLER_28_525 ();
 sg13g2_decap_8 FILLER_28_532 ();
 sg13g2_decap_8 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_546 ();
 sg13g2_decap_8 FILLER_28_553 ();
 sg13g2_decap_8 FILLER_28_560 ();
 sg13g2_decap_8 FILLER_28_567 ();
 sg13g2_decap_8 FILLER_28_574 ();
 sg13g2_decap_8 FILLER_28_581 ();
 sg13g2_decap_8 FILLER_28_588 ();
 sg13g2_decap_8 FILLER_28_595 ();
 sg13g2_decap_8 FILLER_28_602 ();
 sg13g2_decap_8 FILLER_28_609 ();
 sg13g2_decap_8 FILLER_28_616 ();
 sg13g2_decap_8 FILLER_28_623 ();
 sg13g2_decap_8 FILLER_28_630 ();
 sg13g2_decap_8 FILLER_28_637 ();
 sg13g2_decap_8 FILLER_28_644 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_decap_8 FILLER_28_665 ();
 sg13g2_decap_8 FILLER_28_672 ();
 sg13g2_decap_8 FILLER_28_679 ();
 sg13g2_decap_8 FILLER_28_686 ();
 sg13g2_decap_8 FILLER_28_693 ();
 sg13g2_decap_8 FILLER_28_700 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_fill_1 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_8 FILLER_29_189 ();
 sg13g2_decap_8 FILLER_29_196 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_210 ();
 sg13g2_decap_8 FILLER_29_217 ();
 sg13g2_decap_8 FILLER_29_224 ();
 sg13g2_decap_8 FILLER_29_231 ();
 sg13g2_decap_8 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_245 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_8 FILLER_29_273 ();
 sg13g2_decap_8 FILLER_29_280 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_decap_8 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_301 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_decap_8 FILLER_29_427 ();
 sg13g2_decap_8 FILLER_29_434 ();
 sg13g2_decap_8 FILLER_29_441 ();
 sg13g2_decap_8 FILLER_29_448 ();
 sg13g2_decap_8 FILLER_29_455 ();
 sg13g2_decap_8 FILLER_29_462 ();
 sg13g2_decap_8 FILLER_29_469 ();
 sg13g2_decap_8 FILLER_29_476 ();
 sg13g2_decap_8 FILLER_29_483 ();
 sg13g2_decap_8 FILLER_29_490 ();
 sg13g2_decap_8 FILLER_29_497 ();
 sg13g2_decap_8 FILLER_29_504 ();
 sg13g2_decap_8 FILLER_29_511 ();
 sg13g2_decap_8 FILLER_29_518 ();
 sg13g2_decap_8 FILLER_29_525 ();
 sg13g2_decap_8 FILLER_29_532 ();
 sg13g2_decap_8 FILLER_29_539 ();
 sg13g2_decap_8 FILLER_29_546 ();
 sg13g2_decap_8 FILLER_29_553 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_decap_8 FILLER_29_574 ();
 sg13g2_decap_8 FILLER_29_581 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_decap_8 FILLER_29_595 ();
 sg13g2_decap_8 FILLER_29_602 ();
 sg13g2_decap_8 FILLER_29_609 ();
 sg13g2_decap_8 FILLER_29_616 ();
 sg13g2_decap_8 FILLER_29_623 ();
 sg13g2_decap_8 FILLER_29_630 ();
 sg13g2_decap_8 FILLER_29_637 ();
 sg13g2_decap_8 FILLER_29_644 ();
 sg13g2_decap_8 FILLER_29_651 ();
 sg13g2_decap_8 FILLER_29_658 ();
 sg13g2_decap_8 FILLER_29_665 ();
 sg13g2_decap_8 FILLER_29_672 ();
 sg13g2_decap_8 FILLER_29_679 ();
 sg13g2_decap_8 FILLER_29_686 ();
 sg13g2_decap_8 FILLER_29_693 ();
 sg13g2_decap_8 FILLER_29_700 ();
 sg13g2_decap_8 FILLER_29_707 ();
 sg13g2_decap_8 FILLER_29_714 ();
 sg13g2_decap_8 FILLER_29_721 ();
 sg13g2_decap_8 FILLER_29_728 ();
 sg13g2_decap_8 FILLER_29_735 ();
 sg13g2_decap_8 FILLER_29_742 ();
 sg13g2_decap_8 FILLER_29_749 ();
 sg13g2_decap_8 FILLER_29_756 ();
 sg13g2_decap_8 FILLER_29_763 ();
 sg13g2_decap_8 FILLER_29_770 ();
 sg13g2_decap_8 FILLER_29_777 ();
 sg13g2_decap_8 FILLER_29_784 ();
 sg13g2_decap_8 FILLER_29_791 ();
 sg13g2_decap_8 FILLER_29_798 ();
 sg13g2_decap_8 FILLER_29_805 ();
 sg13g2_decap_8 FILLER_29_812 ();
 sg13g2_decap_8 FILLER_29_819 ();
 sg13g2_decap_8 FILLER_29_826 ();
 sg13g2_decap_8 FILLER_29_833 ();
 sg13g2_fill_1 FILLER_29_840 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_427 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_504 ();
 sg13g2_decap_8 FILLER_30_511 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_decap_8 FILLER_30_525 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_decap_8 FILLER_30_539 ();
 sg13g2_decap_8 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_decap_8 FILLER_30_581 ();
 sg13g2_decap_8 FILLER_30_588 ();
 sg13g2_decap_8 FILLER_30_595 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_decap_8 FILLER_30_623 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_fill_1 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_8 FILLER_31_511 ();
 sg13g2_decap_8 FILLER_31_518 ();
 sg13g2_decap_8 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_decap_8 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_567 ();
 sg13g2_decap_8 FILLER_31_574 ();
 sg13g2_decap_8 FILLER_31_581 ();
 sg13g2_decap_8 FILLER_31_588 ();
 sg13g2_decap_8 FILLER_31_595 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_decap_8 FILLER_31_609 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_decap_8 FILLER_31_623 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_8 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_decap_8 FILLER_31_679 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_8 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_763 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_fill_1 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_8 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_203 ();
 sg13g2_decap_8 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_217 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_8 FILLER_32_231 ();
 sg13g2_decap_8 FILLER_32_238 ();
 sg13g2_decap_8 FILLER_32_245 ();
 sg13g2_decap_8 FILLER_32_252 ();
 sg13g2_decap_8 FILLER_32_259 ();
 sg13g2_decap_8 FILLER_32_266 ();
 sg13g2_decap_8 FILLER_32_273 ();
 sg13g2_decap_8 FILLER_32_280 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_8 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_32_406 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_decap_8 FILLER_32_427 ();
 sg13g2_decap_8 FILLER_32_434 ();
 sg13g2_decap_8 FILLER_32_441 ();
 sg13g2_decap_8 FILLER_32_448 ();
 sg13g2_decap_8 FILLER_32_455 ();
 sg13g2_decap_8 FILLER_32_462 ();
 sg13g2_decap_8 FILLER_32_469 ();
 sg13g2_decap_8 FILLER_32_476 ();
 sg13g2_decap_8 FILLER_32_483 ();
 sg13g2_decap_8 FILLER_32_490 ();
 sg13g2_decap_8 FILLER_32_497 ();
 sg13g2_decap_8 FILLER_32_504 ();
 sg13g2_decap_8 FILLER_32_511 ();
 sg13g2_decap_8 FILLER_32_518 ();
 sg13g2_decap_8 FILLER_32_525 ();
 sg13g2_decap_8 FILLER_32_532 ();
 sg13g2_decap_8 FILLER_32_539 ();
 sg13g2_decap_8 FILLER_32_546 ();
 sg13g2_decap_8 FILLER_32_553 ();
 sg13g2_decap_8 FILLER_32_560 ();
 sg13g2_decap_8 FILLER_32_567 ();
 sg13g2_decap_8 FILLER_32_574 ();
 sg13g2_decap_8 FILLER_32_581 ();
 sg13g2_decap_8 FILLER_32_588 ();
 sg13g2_decap_8 FILLER_32_595 ();
 sg13g2_decap_8 FILLER_32_602 ();
 sg13g2_decap_8 FILLER_32_609 ();
 sg13g2_decap_8 FILLER_32_616 ();
 sg13g2_decap_8 FILLER_32_623 ();
 sg13g2_decap_8 FILLER_32_630 ();
 sg13g2_decap_8 FILLER_32_637 ();
 sg13g2_decap_8 FILLER_32_644 ();
 sg13g2_decap_8 FILLER_32_651 ();
 sg13g2_decap_8 FILLER_32_658 ();
 sg13g2_decap_8 FILLER_32_665 ();
 sg13g2_decap_8 FILLER_32_672 ();
 sg13g2_decap_8 FILLER_32_679 ();
 sg13g2_decap_8 FILLER_32_686 ();
 sg13g2_decap_8 FILLER_32_693 ();
 sg13g2_decap_8 FILLER_32_700 ();
 sg13g2_decap_8 FILLER_32_707 ();
 sg13g2_decap_8 FILLER_32_714 ();
 sg13g2_decap_8 FILLER_32_721 ();
 sg13g2_decap_8 FILLER_32_728 ();
 sg13g2_decap_8 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_742 ();
 sg13g2_decap_8 FILLER_32_749 ();
 sg13g2_decap_8 FILLER_32_756 ();
 sg13g2_decap_8 FILLER_32_763 ();
 sg13g2_decap_8 FILLER_32_770 ();
 sg13g2_decap_8 FILLER_32_777 ();
 sg13g2_decap_8 FILLER_32_784 ();
 sg13g2_decap_8 FILLER_32_791 ();
 sg13g2_decap_8 FILLER_32_798 ();
 sg13g2_decap_8 FILLER_32_805 ();
 sg13g2_decap_8 FILLER_32_812 ();
 sg13g2_decap_8 FILLER_32_819 ();
 sg13g2_decap_8 FILLER_32_826 ();
 sg13g2_decap_8 FILLER_32_833 ();
 sg13g2_fill_1 FILLER_32_840 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_441 ();
 sg13g2_decap_8 FILLER_33_448 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_decap_8 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_476 ();
 sg13g2_decap_8 FILLER_33_483 ();
 sg13g2_decap_8 FILLER_33_490 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_decap_8 FILLER_33_511 ();
 sg13g2_decap_8 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_decap_8 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_546 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_decap_8 FILLER_33_560 ();
 sg13g2_decap_8 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_decap_8 FILLER_33_581 ();
 sg13g2_decap_8 FILLER_33_588 ();
 sg13g2_decap_8 FILLER_33_595 ();
 sg13g2_decap_8 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_609 ();
 sg13g2_decap_8 FILLER_33_616 ();
 sg13g2_decap_8 FILLER_33_623 ();
 sg13g2_decap_8 FILLER_33_630 ();
 sg13g2_decap_8 FILLER_33_637 ();
 sg13g2_decap_8 FILLER_33_644 ();
 sg13g2_decap_8 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_decap_8 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_fill_1 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_203 ();
 sg13g2_decap_8 FILLER_34_210 ();
 sg13g2_decap_8 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_224 ();
 sg13g2_decap_8 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_238 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_decap_8 FILLER_34_252 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_decap_8 FILLER_34_280 ();
 sg13g2_decap_8 FILLER_34_287 ();
 sg13g2_decap_8 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_322 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_406 ();
 sg13g2_decap_8 FILLER_34_413 ();
 sg13g2_decap_8 FILLER_34_420 ();
 sg13g2_decap_8 FILLER_34_427 ();
 sg13g2_decap_8 FILLER_34_434 ();
 sg13g2_decap_8 FILLER_34_441 ();
 sg13g2_decap_8 FILLER_34_448 ();
 sg13g2_decap_8 FILLER_34_455 ();
 sg13g2_decap_8 FILLER_34_462 ();
 sg13g2_decap_8 FILLER_34_469 ();
 sg13g2_decap_8 FILLER_34_476 ();
 sg13g2_decap_8 FILLER_34_483 ();
 sg13g2_decap_8 FILLER_34_490 ();
 sg13g2_decap_8 FILLER_34_497 ();
 sg13g2_decap_8 FILLER_34_504 ();
 sg13g2_decap_8 FILLER_34_511 ();
 sg13g2_decap_8 FILLER_34_518 ();
 sg13g2_decap_8 FILLER_34_525 ();
 sg13g2_decap_8 FILLER_34_532 ();
 sg13g2_decap_8 FILLER_34_539 ();
 sg13g2_decap_8 FILLER_34_546 ();
 sg13g2_decap_8 FILLER_34_553 ();
 sg13g2_decap_8 FILLER_34_560 ();
 sg13g2_decap_8 FILLER_34_567 ();
 sg13g2_decap_8 FILLER_34_574 ();
 sg13g2_decap_8 FILLER_34_581 ();
 sg13g2_decap_8 FILLER_34_588 ();
 sg13g2_decap_8 FILLER_34_595 ();
 sg13g2_decap_8 FILLER_34_602 ();
 sg13g2_decap_8 FILLER_34_609 ();
 sg13g2_decap_8 FILLER_34_616 ();
 sg13g2_decap_8 FILLER_34_623 ();
 sg13g2_decap_8 FILLER_34_630 ();
 sg13g2_decap_8 FILLER_34_637 ();
 sg13g2_decap_8 FILLER_34_644 ();
 sg13g2_decap_8 FILLER_34_651 ();
 sg13g2_decap_8 FILLER_34_658 ();
 sg13g2_decap_8 FILLER_34_665 ();
 sg13g2_decap_8 FILLER_34_672 ();
 sg13g2_decap_8 FILLER_34_679 ();
 sg13g2_decap_8 FILLER_34_686 ();
 sg13g2_decap_8 FILLER_34_693 ();
 sg13g2_decap_8 FILLER_34_700 ();
 sg13g2_decap_8 FILLER_34_707 ();
 sg13g2_decap_8 FILLER_34_714 ();
 sg13g2_decap_8 FILLER_34_721 ();
 sg13g2_decap_8 FILLER_34_728 ();
 sg13g2_decap_8 FILLER_34_735 ();
 sg13g2_decap_8 FILLER_34_742 ();
 sg13g2_decap_8 FILLER_34_749 ();
 sg13g2_decap_8 FILLER_34_756 ();
 sg13g2_decap_8 FILLER_34_763 ();
 sg13g2_decap_8 FILLER_34_770 ();
 sg13g2_decap_8 FILLER_34_777 ();
 sg13g2_decap_8 FILLER_34_784 ();
 sg13g2_decap_8 FILLER_34_791 ();
 sg13g2_decap_8 FILLER_34_798 ();
 sg13g2_decap_8 FILLER_34_805 ();
 sg13g2_decap_8 FILLER_34_812 ();
 sg13g2_decap_8 FILLER_34_819 ();
 sg13g2_decap_8 FILLER_34_826 ();
 sg13g2_decap_8 FILLER_34_833 ();
 sg13g2_fill_1 FILLER_34_840 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_decap_8 FILLER_35_427 ();
 sg13g2_decap_8 FILLER_35_434 ();
 sg13g2_decap_8 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_448 ();
 sg13g2_decap_8 FILLER_35_455 ();
 sg13g2_decap_8 FILLER_35_462 ();
 sg13g2_decap_8 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_decap_8 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_490 ();
 sg13g2_decap_8 FILLER_35_497 ();
 sg13g2_decap_8 FILLER_35_504 ();
 sg13g2_decap_8 FILLER_35_511 ();
 sg13g2_decap_8 FILLER_35_518 ();
 sg13g2_decap_8 FILLER_35_525 ();
 sg13g2_decap_8 FILLER_35_532 ();
 sg13g2_decap_8 FILLER_35_539 ();
 sg13g2_decap_8 FILLER_35_546 ();
 sg13g2_decap_8 FILLER_35_553 ();
 sg13g2_decap_8 FILLER_35_560 ();
 sg13g2_decap_8 FILLER_35_567 ();
 sg13g2_decap_8 FILLER_35_574 ();
 sg13g2_decap_8 FILLER_35_581 ();
 sg13g2_decap_8 FILLER_35_588 ();
 sg13g2_decap_8 FILLER_35_595 ();
 sg13g2_decap_8 FILLER_35_602 ();
 sg13g2_decap_8 FILLER_35_609 ();
 sg13g2_decap_8 FILLER_35_616 ();
 sg13g2_decap_8 FILLER_35_623 ();
 sg13g2_decap_8 FILLER_35_630 ();
 sg13g2_decap_8 FILLER_35_637 ();
 sg13g2_decap_8 FILLER_35_644 ();
 sg13g2_decap_8 FILLER_35_651 ();
 sg13g2_decap_8 FILLER_35_658 ();
 sg13g2_decap_8 FILLER_35_665 ();
 sg13g2_decap_8 FILLER_35_672 ();
 sg13g2_decap_8 FILLER_35_679 ();
 sg13g2_decap_8 FILLER_35_686 ();
 sg13g2_decap_8 FILLER_35_693 ();
 sg13g2_decap_8 FILLER_35_700 ();
 sg13g2_decap_8 FILLER_35_707 ();
 sg13g2_decap_8 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_721 ();
 sg13g2_decap_8 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_749 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_777 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_fill_1 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_36_406 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_420 ();
 sg13g2_decap_8 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_434 ();
 sg13g2_decap_8 FILLER_36_441 ();
 sg13g2_decap_8 FILLER_36_448 ();
 sg13g2_decap_8 FILLER_36_455 ();
 sg13g2_decap_8 FILLER_36_462 ();
 sg13g2_decap_8 FILLER_36_469 ();
 sg13g2_decap_8 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_483 ();
 sg13g2_decap_8 FILLER_36_490 ();
 sg13g2_decap_8 FILLER_36_497 ();
 sg13g2_decap_8 FILLER_36_504 ();
 sg13g2_decap_8 FILLER_36_511 ();
 sg13g2_decap_8 FILLER_36_518 ();
 sg13g2_decap_8 FILLER_36_525 ();
 sg13g2_decap_8 FILLER_36_532 ();
 sg13g2_decap_8 FILLER_36_539 ();
 sg13g2_decap_8 FILLER_36_546 ();
 sg13g2_decap_8 FILLER_36_553 ();
 sg13g2_decap_8 FILLER_36_560 ();
 sg13g2_decap_8 FILLER_36_567 ();
 sg13g2_decap_8 FILLER_36_574 ();
 sg13g2_decap_8 FILLER_36_581 ();
 sg13g2_decap_8 FILLER_36_588 ();
 sg13g2_decap_8 FILLER_36_595 ();
 sg13g2_decap_8 FILLER_36_602 ();
 sg13g2_decap_8 FILLER_36_609 ();
 sg13g2_decap_8 FILLER_36_616 ();
 sg13g2_decap_8 FILLER_36_623 ();
 sg13g2_decap_8 FILLER_36_630 ();
 sg13g2_decap_8 FILLER_36_637 ();
 sg13g2_decap_8 FILLER_36_644 ();
 sg13g2_decap_8 FILLER_36_651 ();
 sg13g2_decap_8 FILLER_36_658 ();
 sg13g2_decap_8 FILLER_36_665 ();
 sg13g2_decap_8 FILLER_36_672 ();
 sg13g2_decap_8 FILLER_36_679 ();
 sg13g2_decap_8 FILLER_36_686 ();
 sg13g2_decap_8 FILLER_36_693 ();
 sg13g2_decap_8 FILLER_36_700 ();
 sg13g2_decap_8 FILLER_36_707 ();
 sg13g2_decap_8 FILLER_36_714 ();
 sg13g2_decap_8 FILLER_36_721 ();
 sg13g2_decap_8 FILLER_36_728 ();
 sg13g2_decap_8 FILLER_36_735 ();
 sg13g2_decap_8 FILLER_36_742 ();
 sg13g2_decap_8 FILLER_36_749 ();
 sg13g2_decap_8 FILLER_36_756 ();
 sg13g2_decap_8 FILLER_36_763 ();
 sg13g2_decap_8 FILLER_36_770 ();
 sg13g2_decap_8 FILLER_36_777 ();
 sg13g2_decap_8 FILLER_36_784 ();
 sg13g2_decap_8 FILLER_36_791 ();
 sg13g2_decap_8 FILLER_36_798 ();
 sg13g2_decap_8 FILLER_36_805 ();
 sg13g2_decap_8 FILLER_36_812 ();
 sg13g2_decap_8 FILLER_36_819 ();
 sg13g2_decap_8 FILLER_36_826 ();
 sg13g2_decap_8 FILLER_36_833 ();
 sg13g2_fill_1 FILLER_36_840 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_497 ();
 sg13g2_decap_8 FILLER_37_504 ();
 sg13g2_decap_8 FILLER_37_511 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_525 ();
 sg13g2_decap_8 FILLER_37_532 ();
 sg13g2_decap_8 FILLER_37_539 ();
 sg13g2_decap_8 FILLER_37_546 ();
 sg13g2_decap_8 FILLER_37_553 ();
 sg13g2_decap_8 FILLER_37_560 ();
 sg13g2_decap_8 FILLER_37_567 ();
 sg13g2_decap_8 FILLER_37_574 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_595 ();
 sg13g2_decap_8 FILLER_37_602 ();
 sg13g2_decap_8 FILLER_37_609 ();
 sg13g2_decap_8 FILLER_37_616 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_decap_8 FILLER_37_651 ();
 sg13g2_decap_8 FILLER_37_658 ();
 sg13g2_decap_8 FILLER_37_665 ();
 sg13g2_decap_8 FILLER_37_672 ();
 sg13g2_decap_8 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_721 ();
 sg13g2_decap_8 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_742 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_fill_1 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_decap_8 FILLER_38_427 ();
 sg13g2_decap_8 FILLER_38_434 ();
 sg13g2_decap_8 FILLER_38_441 ();
 sg13g2_decap_8 FILLER_38_448 ();
 sg13g2_decap_8 FILLER_38_455 ();
 sg13g2_decap_8 FILLER_38_462 ();
 sg13g2_decap_8 FILLER_38_469 ();
 sg13g2_decap_8 FILLER_38_476 ();
 sg13g2_decap_8 FILLER_38_483 ();
 sg13g2_decap_8 FILLER_38_490 ();
 sg13g2_decap_8 FILLER_38_497 ();
 sg13g2_decap_8 FILLER_38_504 ();
 sg13g2_decap_8 FILLER_38_511 ();
 sg13g2_decap_8 FILLER_38_518 ();
 sg13g2_decap_8 FILLER_38_525 ();
 sg13g2_decap_8 FILLER_38_532 ();
 sg13g2_decap_8 FILLER_38_539 ();
 sg13g2_decap_8 FILLER_38_546 ();
 sg13g2_decap_8 FILLER_38_553 ();
 sg13g2_decap_8 FILLER_38_560 ();
 sg13g2_decap_8 FILLER_38_567 ();
 sg13g2_decap_8 FILLER_38_574 ();
 sg13g2_decap_8 FILLER_38_581 ();
 sg13g2_decap_8 FILLER_38_588 ();
 sg13g2_decap_8 FILLER_38_595 ();
 sg13g2_decap_8 FILLER_38_602 ();
 sg13g2_decap_8 FILLER_38_609 ();
 sg13g2_decap_8 FILLER_38_616 ();
 sg13g2_decap_8 FILLER_38_623 ();
 sg13g2_decap_8 FILLER_38_630 ();
 sg13g2_decap_8 FILLER_38_637 ();
 sg13g2_decap_8 FILLER_38_644 ();
 sg13g2_decap_8 FILLER_38_651 ();
 sg13g2_decap_8 FILLER_38_658 ();
 sg13g2_decap_8 FILLER_38_665 ();
 sg13g2_decap_8 FILLER_38_672 ();
 sg13g2_decap_8 FILLER_38_679 ();
 sg13g2_decap_8 FILLER_38_686 ();
 sg13g2_decap_8 FILLER_38_693 ();
 sg13g2_decap_8 FILLER_38_700 ();
 sg13g2_decap_8 FILLER_38_707 ();
 sg13g2_decap_8 FILLER_38_714 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_decap_8 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_decap_8 FILLER_38_756 ();
 sg13g2_decap_8 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_770 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_8 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_826 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_fill_1 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_decap_8 FILLER_39_427 ();
 sg13g2_decap_8 FILLER_39_434 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_decap_8 FILLER_39_462 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_decap_8 FILLER_39_476 ();
 sg13g2_decap_8 FILLER_39_483 ();
 sg13g2_decap_8 FILLER_39_490 ();
 sg13g2_decap_8 FILLER_39_497 ();
 sg13g2_decap_8 FILLER_39_504 ();
 sg13g2_decap_8 FILLER_39_511 ();
 sg13g2_decap_8 FILLER_39_518 ();
 sg13g2_decap_8 FILLER_39_525 ();
 sg13g2_decap_8 FILLER_39_532 ();
 sg13g2_decap_8 FILLER_39_539 ();
 sg13g2_decap_8 FILLER_39_546 ();
 sg13g2_decap_8 FILLER_39_553 ();
 sg13g2_decap_8 FILLER_39_560 ();
 sg13g2_decap_8 FILLER_39_567 ();
 sg13g2_decap_8 FILLER_39_574 ();
 sg13g2_decap_8 FILLER_39_581 ();
 sg13g2_decap_8 FILLER_39_588 ();
 sg13g2_decap_8 FILLER_39_595 ();
 sg13g2_decap_8 FILLER_39_602 ();
 sg13g2_decap_8 FILLER_39_609 ();
 sg13g2_decap_8 FILLER_39_616 ();
 sg13g2_decap_8 FILLER_39_623 ();
 sg13g2_decap_8 FILLER_39_630 ();
 sg13g2_decap_8 FILLER_39_637 ();
 sg13g2_decap_8 FILLER_39_644 ();
 sg13g2_decap_8 FILLER_39_651 ();
 sg13g2_decap_8 FILLER_39_658 ();
 sg13g2_decap_8 FILLER_39_665 ();
 sg13g2_decap_8 FILLER_39_672 ();
 sg13g2_decap_8 FILLER_39_679 ();
 sg13g2_decap_8 FILLER_39_686 ();
 sg13g2_decap_8 FILLER_39_693 ();
 sg13g2_decap_8 FILLER_39_700 ();
 sg13g2_decap_8 FILLER_39_707 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_decap_8 FILLER_39_721 ();
 sg13g2_decap_8 FILLER_39_728 ();
 sg13g2_decap_8 FILLER_39_735 ();
 sg13g2_decap_8 FILLER_39_742 ();
 sg13g2_decap_8 FILLER_39_749 ();
 sg13g2_decap_8 FILLER_39_756 ();
 sg13g2_decap_8 FILLER_39_763 ();
 sg13g2_decap_8 FILLER_39_770 ();
 sg13g2_decap_8 FILLER_39_777 ();
 sg13g2_decap_8 FILLER_39_784 ();
 sg13g2_decap_8 FILLER_39_791 ();
 sg13g2_decap_8 FILLER_39_798 ();
 sg13g2_decap_8 FILLER_39_805 ();
 sg13g2_decap_8 FILLER_39_812 ();
 sg13g2_decap_8 FILLER_39_819 ();
 sg13g2_decap_8 FILLER_39_826 ();
 sg13g2_decap_8 FILLER_39_833 ();
 sg13g2_fill_1 FILLER_39_840 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_497 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_decap_8 FILLER_40_511 ();
 sg13g2_decap_8 FILLER_40_518 ();
 sg13g2_decap_8 FILLER_40_525 ();
 sg13g2_decap_8 FILLER_40_532 ();
 sg13g2_decap_8 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_546 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_decap_8 FILLER_40_560 ();
 sg13g2_decap_8 FILLER_40_567 ();
 sg13g2_decap_8 FILLER_40_574 ();
 sg13g2_decap_8 FILLER_40_581 ();
 sg13g2_decap_8 FILLER_40_588 ();
 sg13g2_decap_8 FILLER_40_595 ();
 sg13g2_decap_8 FILLER_40_602 ();
 sg13g2_decap_8 FILLER_40_609 ();
 sg13g2_decap_8 FILLER_40_616 ();
 sg13g2_decap_8 FILLER_40_623 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_decap_8 FILLER_40_644 ();
 sg13g2_decap_8 FILLER_40_651 ();
 sg13g2_decap_8 FILLER_40_658 ();
 sg13g2_decap_8 FILLER_40_665 ();
 sg13g2_decap_8 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_679 ();
 sg13g2_decap_8 FILLER_40_686 ();
 sg13g2_decap_8 FILLER_40_693 ();
 sg13g2_decap_8 FILLER_40_700 ();
 sg13g2_decap_8 FILLER_40_707 ();
 sg13g2_decap_8 FILLER_40_714 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_decap_8 FILLER_40_728 ();
 sg13g2_decap_8 FILLER_40_735 ();
 sg13g2_decap_8 FILLER_40_742 ();
 sg13g2_decap_8 FILLER_40_749 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_791 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_805 ();
 sg13g2_decap_8 FILLER_40_812 ();
 sg13g2_decap_8 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_decap_8 FILLER_40_833 ();
 sg13g2_fill_1 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_8 FILLER_41_441 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_decap_8 FILLER_41_455 ();
 sg13g2_decap_8 FILLER_41_462 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_8 FILLER_41_497 ();
 sg13g2_decap_8 FILLER_41_504 ();
 sg13g2_decap_8 FILLER_41_511 ();
 sg13g2_decap_8 FILLER_41_518 ();
 sg13g2_decap_8 FILLER_41_525 ();
 sg13g2_decap_8 FILLER_41_532 ();
 sg13g2_decap_8 FILLER_41_539 ();
 sg13g2_decap_8 FILLER_41_546 ();
 sg13g2_decap_8 FILLER_41_553 ();
 sg13g2_decap_8 FILLER_41_560 ();
 sg13g2_decap_8 FILLER_41_567 ();
 sg13g2_decap_8 FILLER_41_574 ();
 sg13g2_decap_8 FILLER_41_581 ();
 sg13g2_decap_8 FILLER_41_588 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_decap_8 FILLER_41_602 ();
 sg13g2_decap_8 FILLER_41_609 ();
 sg13g2_decap_8 FILLER_41_616 ();
 sg13g2_decap_8 FILLER_41_623 ();
 sg13g2_decap_8 FILLER_41_630 ();
 sg13g2_decap_8 FILLER_41_637 ();
 sg13g2_decap_8 FILLER_41_644 ();
 sg13g2_decap_8 FILLER_41_651 ();
 sg13g2_decap_8 FILLER_41_658 ();
 sg13g2_decap_8 FILLER_41_665 ();
 sg13g2_decap_8 FILLER_41_672 ();
 sg13g2_decap_8 FILLER_41_679 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_8 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_707 ();
 sg13g2_decap_8 FILLER_41_714 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_728 ();
 sg13g2_decap_8 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_fill_1 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_decap_8 FILLER_42_196 ();
 sg13g2_decap_8 FILLER_42_203 ();
 sg13g2_decap_8 FILLER_42_210 ();
 sg13g2_decap_8 FILLER_42_217 ();
 sg13g2_decap_8 FILLER_42_224 ();
 sg13g2_decap_8 FILLER_42_231 ();
 sg13g2_decap_8 FILLER_42_238 ();
 sg13g2_decap_8 FILLER_42_245 ();
 sg13g2_decap_8 FILLER_42_252 ();
 sg13g2_decap_8 FILLER_42_259 ();
 sg13g2_decap_8 FILLER_42_266 ();
 sg13g2_decap_8 FILLER_42_273 ();
 sg13g2_decap_8 FILLER_42_280 ();
 sg13g2_decap_8 FILLER_42_287 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_decap_8 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_315 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_8 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_decap_8 FILLER_42_406 ();
 sg13g2_decap_8 FILLER_42_413 ();
 sg13g2_decap_8 FILLER_42_420 ();
 sg13g2_decap_8 FILLER_42_427 ();
 sg13g2_decap_8 FILLER_42_434 ();
 sg13g2_decap_8 FILLER_42_441 ();
 sg13g2_decap_8 FILLER_42_448 ();
 sg13g2_decap_8 FILLER_42_455 ();
 sg13g2_decap_8 FILLER_42_462 ();
 sg13g2_decap_8 FILLER_42_469 ();
 sg13g2_decap_8 FILLER_42_476 ();
 sg13g2_decap_8 FILLER_42_483 ();
 sg13g2_decap_8 FILLER_42_490 ();
 sg13g2_decap_8 FILLER_42_497 ();
 sg13g2_decap_8 FILLER_42_504 ();
 sg13g2_decap_8 FILLER_42_511 ();
 sg13g2_decap_8 FILLER_42_518 ();
 sg13g2_decap_8 FILLER_42_525 ();
 sg13g2_decap_8 FILLER_42_532 ();
 sg13g2_decap_8 FILLER_42_539 ();
 sg13g2_decap_8 FILLER_42_546 ();
 sg13g2_decap_8 FILLER_42_553 ();
 sg13g2_decap_8 FILLER_42_560 ();
 sg13g2_decap_8 FILLER_42_567 ();
 sg13g2_decap_8 FILLER_42_574 ();
 sg13g2_decap_8 FILLER_42_581 ();
 sg13g2_decap_8 FILLER_42_588 ();
 sg13g2_decap_8 FILLER_42_595 ();
 sg13g2_decap_8 FILLER_42_602 ();
 sg13g2_decap_8 FILLER_42_609 ();
 sg13g2_decap_8 FILLER_42_616 ();
 sg13g2_decap_8 FILLER_42_623 ();
 sg13g2_decap_8 FILLER_42_630 ();
 sg13g2_decap_8 FILLER_42_637 ();
 sg13g2_decap_8 FILLER_42_644 ();
 sg13g2_decap_8 FILLER_42_651 ();
 sg13g2_decap_8 FILLER_42_658 ();
 sg13g2_decap_8 FILLER_42_665 ();
 sg13g2_decap_8 FILLER_42_672 ();
 sg13g2_decap_8 FILLER_42_679 ();
 sg13g2_decap_8 FILLER_42_686 ();
 sg13g2_decap_8 FILLER_42_693 ();
 sg13g2_decap_8 FILLER_42_700 ();
 sg13g2_decap_8 FILLER_42_707 ();
 sg13g2_decap_8 FILLER_42_714 ();
 sg13g2_decap_8 FILLER_42_721 ();
 sg13g2_decap_8 FILLER_42_728 ();
 sg13g2_decap_8 FILLER_42_735 ();
 sg13g2_decap_8 FILLER_42_742 ();
 sg13g2_decap_8 FILLER_42_749 ();
 sg13g2_decap_8 FILLER_42_756 ();
 sg13g2_decap_8 FILLER_42_763 ();
 sg13g2_decap_8 FILLER_42_770 ();
 sg13g2_decap_8 FILLER_42_777 ();
 sg13g2_decap_8 FILLER_42_784 ();
 sg13g2_decap_8 FILLER_42_791 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_decap_8 FILLER_42_819 ();
 sg13g2_decap_8 FILLER_42_826 ();
 sg13g2_decap_8 FILLER_42_833 ();
 sg13g2_fill_1 FILLER_42_840 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_decap_8 FILLER_43_476 ();
 sg13g2_decap_8 FILLER_43_483 ();
 sg13g2_decap_8 FILLER_43_490 ();
 sg13g2_decap_8 FILLER_43_497 ();
 sg13g2_decap_8 FILLER_43_504 ();
 sg13g2_decap_8 FILLER_43_511 ();
 sg13g2_decap_8 FILLER_43_518 ();
 sg13g2_decap_8 FILLER_43_525 ();
 sg13g2_decap_8 FILLER_43_532 ();
 sg13g2_decap_8 FILLER_43_539 ();
 sg13g2_decap_8 FILLER_43_546 ();
 sg13g2_decap_8 FILLER_43_553 ();
 sg13g2_decap_8 FILLER_43_560 ();
 sg13g2_decap_8 FILLER_43_567 ();
 sg13g2_decap_8 FILLER_43_574 ();
 sg13g2_decap_8 FILLER_43_581 ();
 sg13g2_decap_8 FILLER_43_588 ();
 sg13g2_decap_8 FILLER_43_595 ();
 sg13g2_decap_8 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_609 ();
 sg13g2_decap_8 FILLER_43_616 ();
 sg13g2_decap_8 FILLER_43_623 ();
 sg13g2_decap_8 FILLER_43_630 ();
 sg13g2_decap_8 FILLER_43_637 ();
 sg13g2_decap_8 FILLER_43_644 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_decap_8 FILLER_43_665 ();
 sg13g2_decap_8 FILLER_43_672 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_decap_8 FILLER_43_686 ();
 sg13g2_decap_8 FILLER_43_693 ();
 sg13g2_decap_8 FILLER_43_700 ();
 sg13g2_decap_8 FILLER_43_707 ();
 sg13g2_decap_8 FILLER_43_714 ();
 sg13g2_decap_8 FILLER_43_721 ();
 sg13g2_decap_8 FILLER_43_728 ();
 sg13g2_decap_8 FILLER_43_735 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_decap_8 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_756 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_fill_1 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_8 FILLER_44_203 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_decap_8 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_224 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_decap_8 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_decap_8 FILLER_44_252 ();
 sg13g2_decap_8 FILLER_44_259 ();
 sg13g2_decap_8 FILLER_44_266 ();
 sg13g2_decap_8 FILLER_44_273 ();
 sg13g2_decap_8 FILLER_44_280 ();
 sg13g2_decap_8 FILLER_44_287 ();
 sg13g2_decap_8 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_301 ();
 sg13g2_decap_8 FILLER_44_308 ();
 sg13g2_decap_8 FILLER_44_315 ();
 sg13g2_decap_8 FILLER_44_322 ();
 sg13g2_decap_8 FILLER_44_329 ();
 sg13g2_decap_8 FILLER_44_336 ();
 sg13g2_decap_8 FILLER_44_343 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_decap_8 FILLER_44_406 ();
 sg13g2_decap_8 FILLER_44_413 ();
 sg13g2_decap_8 FILLER_44_420 ();
 sg13g2_decap_8 FILLER_44_427 ();
 sg13g2_decap_8 FILLER_44_434 ();
 sg13g2_decap_8 FILLER_44_441 ();
 sg13g2_decap_8 FILLER_44_448 ();
 sg13g2_decap_8 FILLER_44_455 ();
 sg13g2_decap_8 FILLER_44_462 ();
 sg13g2_decap_8 FILLER_44_469 ();
 sg13g2_decap_8 FILLER_44_476 ();
 sg13g2_decap_8 FILLER_44_483 ();
 sg13g2_decap_8 FILLER_44_490 ();
 sg13g2_decap_8 FILLER_44_497 ();
 sg13g2_decap_8 FILLER_44_504 ();
 sg13g2_decap_8 FILLER_44_511 ();
 sg13g2_decap_8 FILLER_44_518 ();
 sg13g2_decap_8 FILLER_44_525 ();
 sg13g2_decap_8 FILLER_44_532 ();
 sg13g2_decap_8 FILLER_44_539 ();
 sg13g2_decap_8 FILLER_44_546 ();
 sg13g2_decap_8 FILLER_44_553 ();
 sg13g2_decap_8 FILLER_44_560 ();
 sg13g2_decap_8 FILLER_44_567 ();
 sg13g2_decap_8 FILLER_44_574 ();
 sg13g2_decap_8 FILLER_44_581 ();
 sg13g2_decap_8 FILLER_44_588 ();
 sg13g2_decap_8 FILLER_44_595 ();
 sg13g2_decap_8 FILLER_44_602 ();
 sg13g2_decap_8 FILLER_44_609 ();
 sg13g2_decap_8 FILLER_44_616 ();
 sg13g2_decap_8 FILLER_44_623 ();
 sg13g2_decap_8 FILLER_44_630 ();
 sg13g2_decap_8 FILLER_44_637 ();
 sg13g2_decap_8 FILLER_44_644 ();
 sg13g2_decap_8 FILLER_44_651 ();
 sg13g2_decap_8 FILLER_44_658 ();
 sg13g2_decap_8 FILLER_44_665 ();
 sg13g2_decap_8 FILLER_44_672 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_decap_8 FILLER_44_686 ();
 sg13g2_decap_8 FILLER_44_693 ();
 sg13g2_decap_8 FILLER_44_700 ();
 sg13g2_decap_8 FILLER_44_707 ();
 sg13g2_decap_8 FILLER_44_714 ();
 sg13g2_decap_8 FILLER_44_721 ();
 sg13g2_decap_8 FILLER_44_728 ();
 sg13g2_decap_8 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_742 ();
 sg13g2_decap_8 FILLER_44_749 ();
 sg13g2_decap_8 FILLER_44_756 ();
 sg13g2_decap_8 FILLER_44_763 ();
 sg13g2_decap_8 FILLER_44_770 ();
 sg13g2_decap_8 FILLER_44_777 ();
 sg13g2_decap_8 FILLER_44_784 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_812 ();
 sg13g2_decap_8 FILLER_44_819 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_decap_8 FILLER_44_833 ();
 sg13g2_fill_1 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_469 ();
 sg13g2_decap_8 FILLER_45_476 ();
 sg13g2_decap_8 FILLER_45_483 ();
 sg13g2_decap_8 FILLER_45_490 ();
 sg13g2_decap_8 FILLER_45_497 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_decap_8 FILLER_45_511 ();
 sg13g2_decap_8 FILLER_45_518 ();
 sg13g2_decap_8 FILLER_45_525 ();
 sg13g2_decap_8 FILLER_45_532 ();
 sg13g2_decap_8 FILLER_45_539 ();
 sg13g2_decap_8 FILLER_45_546 ();
 sg13g2_decap_8 FILLER_45_553 ();
 sg13g2_decap_8 FILLER_45_560 ();
 sg13g2_decap_8 FILLER_45_567 ();
 sg13g2_decap_8 FILLER_45_574 ();
 sg13g2_decap_8 FILLER_45_581 ();
 sg13g2_decap_8 FILLER_45_588 ();
 sg13g2_decap_8 FILLER_45_595 ();
 sg13g2_decap_8 FILLER_45_602 ();
 sg13g2_decap_8 FILLER_45_609 ();
 sg13g2_decap_8 FILLER_45_616 ();
 sg13g2_decap_8 FILLER_45_623 ();
 sg13g2_decap_8 FILLER_45_630 ();
 sg13g2_decap_8 FILLER_45_637 ();
 sg13g2_decap_8 FILLER_45_644 ();
 sg13g2_decap_8 FILLER_45_651 ();
 sg13g2_decap_8 FILLER_45_658 ();
 sg13g2_decap_8 FILLER_45_665 ();
 sg13g2_decap_8 FILLER_45_672 ();
 sg13g2_decap_8 FILLER_45_679 ();
 sg13g2_decap_8 FILLER_45_686 ();
 sg13g2_decap_8 FILLER_45_693 ();
 sg13g2_decap_8 FILLER_45_700 ();
 sg13g2_decap_8 FILLER_45_707 ();
 sg13g2_decap_8 FILLER_45_714 ();
 sg13g2_decap_8 FILLER_45_721 ();
 sg13g2_decap_8 FILLER_45_728 ();
 sg13g2_decap_8 FILLER_45_735 ();
 sg13g2_decap_8 FILLER_45_742 ();
 sg13g2_decap_8 FILLER_45_749 ();
 sg13g2_decap_8 FILLER_45_756 ();
 sg13g2_decap_8 FILLER_45_763 ();
 sg13g2_decap_8 FILLER_45_770 ();
 sg13g2_decap_8 FILLER_45_777 ();
 sg13g2_decap_8 FILLER_45_784 ();
 sg13g2_decap_8 FILLER_45_791 ();
 sg13g2_decap_8 FILLER_45_798 ();
 sg13g2_decap_8 FILLER_45_805 ();
 sg13g2_decap_8 FILLER_45_812 ();
 sg13g2_decap_8 FILLER_45_819 ();
 sg13g2_decap_8 FILLER_45_826 ();
 sg13g2_decap_8 FILLER_45_833 ();
 sg13g2_fill_1 FILLER_45_840 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_8 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_8 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_decap_8 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_602 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_8 FILLER_46_637 ();
 sg13g2_decap_8 FILLER_46_644 ();
 sg13g2_decap_8 FILLER_46_651 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_665 ();
 sg13g2_decap_8 FILLER_46_672 ();
 sg13g2_decap_8 FILLER_46_679 ();
 sg13g2_decap_8 FILLER_46_686 ();
 sg13g2_decap_8 FILLER_46_693 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_8 FILLER_46_721 ();
 sg13g2_decap_8 FILLER_46_728 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_756 ();
 sg13g2_decap_8 FILLER_46_763 ();
 sg13g2_decap_8 FILLER_46_770 ();
 sg13g2_decap_8 FILLER_46_777 ();
 sg13g2_decap_8 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_decap_8 FILLER_46_798 ();
 sg13g2_decap_8 FILLER_46_805 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_decap_8 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_fill_1 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_8 FILLER_47_574 ();
 sg13g2_decap_8 FILLER_47_581 ();
 sg13g2_decap_8 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_8 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_8 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_fill_1 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_609 ();
 sg13g2_decap_8 FILLER_48_616 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_decap_8 FILLER_48_630 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_decap_8 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_8 FILLER_48_700 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_735 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_fill_1 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_406 ();
 sg13g2_decap_8 FILLER_49_413 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_decap_8 FILLER_49_427 ();
 sg13g2_decap_8 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_8 FILLER_49_455 ();
 sg13g2_decap_8 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_469 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_8 FILLER_49_483 ();
 sg13g2_decap_8 FILLER_49_490 ();
 sg13g2_decap_8 FILLER_49_497 ();
 sg13g2_decap_8 FILLER_49_504 ();
 sg13g2_decap_8 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_574 ();
 sg13g2_decap_8 FILLER_49_581 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_644 ();
 sg13g2_decap_8 FILLER_49_651 ();
 sg13g2_decap_8 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_decap_8 FILLER_49_672 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_decap_8 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_decap_8 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_8 FILLER_49_784 ();
 sg13g2_decap_8 FILLER_49_791 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_fill_1 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_147 ();
 sg13g2_decap_8 FILLER_50_154 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_decap_8 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_175 ();
 sg13g2_decap_8 FILLER_50_182 ();
 sg13g2_decap_8 FILLER_50_189 ();
 sg13g2_decap_8 FILLER_50_196 ();
 sg13g2_decap_8 FILLER_50_203 ();
 sg13g2_decap_8 FILLER_50_210 ();
 sg13g2_decap_8 FILLER_50_217 ();
 sg13g2_decap_8 FILLER_50_224 ();
 sg13g2_decap_8 FILLER_50_231 ();
 sg13g2_decap_8 FILLER_50_238 ();
 sg13g2_decap_8 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_252 ();
 sg13g2_decap_8 FILLER_50_259 ();
 sg13g2_decap_8 FILLER_50_266 ();
 sg13g2_decap_8 FILLER_50_273 ();
 sg13g2_decap_8 FILLER_50_280 ();
 sg13g2_decap_8 FILLER_50_287 ();
 sg13g2_decap_8 FILLER_50_294 ();
 sg13g2_decap_8 FILLER_50_301 ();
 sg13g2_decap_8 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_315 ();
 sg13g2_decap_8 FILLER_50_322 ();
 sg13g2_decap_8 FILLER_50_329 ();
 sg13g2_decap_8 FILLER_50_336 ();
 sg13g2_decap_8 FILLER_50_343 ();
 sg13g2_decap_8 FILLER_50_350 ();
 sg13g2_decap_8 FILLER_50_357 ();
 sg13g2_decap_8 FILLER_50_364 ();
 sg13g2_decap_8 FILLER_50_371 ();
 sg13g2_decap_8 FILLER_50_378 ();
 sg13g2_decap_8 FILLER_50_385 ();
 sg13g2_decap_8 FILLER_50_392 ();
 sg13g2_decap_8 FILLER_50_399 ();
 sg13g2_decap_8 FILLER_50_406 ();
 sg13g2_decap_8 FILLER_50_413 ();
 sg13g2_decap_8 FILLER_50_420 ();
 sg13g2_decap_8 FILLER_50_427 ();
 sg13g2_decap_8 FILLER_50_434 ();
 sg13g2_decap_8 FILLER_50_441 ();
 sg13g2_decap_8 FILLER_50_448 ();
 sg13g2_decap_8 FILLER_50_455 ();
 sg13g2_decap_8 FILLER_50_462 ();
 sg13g2_decap_8 FILLER_50_469 ();
 sg13g2_decap_8 FILLER_50_476 ();
 sg13g2_decap_8 FILLER_50_483 ();
 sg13g2_decap_8 FILLER_50_490 ();
 sg13g2_decap_8 FILLER_50_497 ();
 sg13g2_decap_8 FILLER_50_504 ();
 sg13g2_decap_8 FILLER_50_511 ();
 sg13g2_decap_8 FILLER_50_518 ();
 sg13g2_decap_8 FILLER_50_525 ();
 sg13g2_decap_8 FILLER_50_532 ();
 sg13g2_decap_8 FILLER_50_539 ();
 sg13g2_decap_8 FILLER_50_546 ();
 sg13g2_decap_8 FILLER_50_553 ();
 sg13g2_decap_8 FILLER_50_560 ();
 sg13g2_decap_8 FILLER_50_567 ();
 sg13g2_decap_8 FILLER_50_574 ();
 sg13g2_decap_8 FILLER_50_581 ();
 sg13g2_decap_8 FILLER_50_588 ();
 sg13g2_decap_8 FILLER_50_595 ();
 sg13g2_decap_8 FILLER_50_602 ();
 sg13g2_decap_8 FILLER_50_609 ();
 sg13g2_decap_8 FILLER_50_616 ();
 sg13g2_decap_8 FILLER_50_623 ();
 sg13g2_decap_8 FILLER_50_630 ();
 sg13g2_decap_8 FILLER_50_637 ();
 sg13g2_decap_8 FILLER_50_644 ();
 sg13g2_decap_8 FILLER_50_651 ();
 sg13g2_decap_8 FILLER_50_658 ();
 sg13g2_decap_8 FILLER_50_665 ();
 sg13g2_decap_8 FILLER_50_672 ();
 sg13g2_decap_8 FILLER_50_679 ();
 sg13g2_decap_8 FILLER_50_686 ();
 sg13g2_decap_8 FILLER_50_693 ();
 sg13g2_decap_8 FILLER_50_700 ();
 sg13g2_decap_8 FILLER_50_707 ();
 sg13g2_decap_8 FILLER_50_714 ();
 sg13g2_decap_8 FILLER_50_721 ();
 sg13g2_decap_8 FILLER_50_728 ();
 sg13g2_decap_8 FILLER_50_735 ();
 sg13g2_decap_8 FILLER_50_742 ();
 sg13g2_decap_8 FILLER_50_749 ();
 sg13g2_decap_8 FILLER_50_756 ();
 sg13g2_decap_8 FILLER_50_763 ();
 sg13g2_decap_8 FILLER_50_770 ();
 sg13g2_decap_8 FILLER_50_777 ();
 sg13g2_decap_8 FILLER_50_784 ();
 sg13g2_decap_8 FILLER_50_791 ();
 sg13g2_decap_8 FILLER_50_798 ();
 sg13g2_decap_8 FILLER_50_805 ();
 sg13g2_decap_8 FILLER_50_812 ();
 sg13g2_decap_8 FILLER_50_819 ();
 sg13g2_decap_8 FILLER_50_826 ();
 sg13g2_decap_8 FILLER_50_833 ();
 sg13g2_fill_1 FILLER_50_840 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_175 ();
 sg13g2_decap_8 FILLER_51_182 ();
 sg13g2_decap_8 FILLER_51_189 ();
 sg13g2_decap_8 FILLER_51_196 ();
 sg13g2_decap_8 FILLER_51_203 ();
 sg13g2_decap_8 FILLER_51_210 ();
 sg13g2_decap_8 FILLER_51_217 ();
 sg13g2_decap_8 FILLER_51_224 ();
 sg13g2_decap_8 FILLER_51_231 ();
 sg13g2_decap_8 FILLER_51_238 ();
 sg13g2_decap_8 FILLER_51_245 ();
 sg13g2_decap_8 FILLER_51_252 ();
 sg13g2_decap_8 FILLER_51_259 ();
 sg13g2_decap_8 FILLER_51_266 ();
 sg13g2_decap_8 FILLER_51_273 ();
 sg13g2_decap_8 FILLER_51_280 ();
 sg13g2_decap_8 FILLER_51_287 ();
 sg13g2_decap_8 FILLER_51_294 ();
 sg13g2_decap_8 FILLER_51_301 ();
 sg13g2_decap_8 FILLER_51_308 ();
 sg13g2_decap_8 FILLER_51_315 ();
 sg13g2_decap_8 FILLER_51_322 ();
 sg13g2_decap_8 FILLER_51_329 ();
 sg13g2_decap_8 FILLER_51_336 ();
 sg13g2_decap_8 FILLER_51_343 ();
 sg13g2_decap_8 FILLER_51_350 ();
 sg13g2_decap_8 FILLER_51_357 ();
 sg13g2_decap_8 FILLER_51_364 ();
 sg13g2_decap_8 FILLER_51_371 ();
 sg13g2_decap_8 FILLER_51_378 ();
 sg13g2_decap_8 FILLER_51_385 ();
 sg13g2_decap_8 FILLER_51_392 ();
 sg13g2_decap_8 FILLER_51_399 ();
 sg13g2_decap_8 FILLER_51_406 ();
 sg13g2_decap_8 FILLER_51_413 ();
 sg13g2_decap_8 FILLER_51_420 ();
 sg13g2_decap_8 FILLER_51_427 ();
 sg13g2_decap_8 FILLER_51_434 ();
 sg13g2_decap_8 FILLER_51_441 ();
 sg13g2_decap_8 FILLER_51_448 ();
 sg13g2_decap_8 FILLER_51_455 ();
 sg13g2_decap_8 FILLER_51_462 ();
 sg13g2_decap_8 FILLER_51_469 ();
 sg13g2_decap_8 FILLER_51_476 ();
 sg13g2_decap_8 FILLER_51_483 ();
 sg13g2_decap_8 FILLER_51_490 ();
 sg13g2_decap_8 FILLER_51_497 ();
 sg13g2_decap_8 FILLER_51_504 ();
 sg13g2_decap_8 FILLER_51_511 ();
 sg13g2_decap_8 FILLER_51_518 ();
 sg13g2_decap_8 FILLER_51_525 ();
 sg13g2_decap_8 FILLER_51_532 ();
 sg13g2_decap_8 FILLER_51_539 ();
 sg13g2_decap_8 FILLER_51_546 ();
 sg13g2_decap_8 FILLER_51_553 ();
 sg13g2_decap_8 FILLER_51_560 ();
 sg13g2_decap_8 FILLER_51_567 ();
 sg13g2_decap_8 FILLER_51_574 ();
 sg13g2_decap_8 FILLER_51_581 ();
 sg13g2_decap_8 FILLER_51_588 ();
 sg13g2_decap_8 FILLER_51_595 ();
 sg13g2_decap_8 FILLER_51_602 ();
 sg13g2_decap_8 FILLER_51_609 ();
 sg13g2_decap_8 FILLER_51_616 ();
 sg13g2_decap_8 FILLER_51_623 ();
 sg13g2_decap_8 FILLER_51_630 ();
 sg13g2_decap_8 FILLER_51_637 ();
 sg13g2_decap_8 FILLER_51_644 ();
 sg13g2_decap_8 FILLER_51_651 ();
 sg13g2_decap_8 FILLER_51_658 ();
 sg13g2_decap_8 FILLER_51_665 ();
 sg13g2_decap_8 FILLER_51_672 ();
 sg13g2_decap_8 FILLER_51_679 ();
 sg13g2_decap_8 FILLER_51_686 ();
 sg13g2_decap_8 FILLER_51_693 ();
 sg13g2_decap_8 FILLER_51_700 ();
 sg13g2_decap_8 FILLER_51_707 ();
 sg13g2_decap_8 FILLER_51_714 ();
 sg13g2_decap_8 FILLER_51_721 ();
 sg13g2_decap_8 FILLER_51_728 ();
 sg13g2_decap_8 FILLER_51_735 ();
 sg13g2_decap_8 FILLER_51_742 ();
 sg13g2_decap_8 FILLER_51_749 ();
 sg13g2_decap_8 FILLER_51_756 ();
 sg13g2_decap_8 FILLER_51_763 ();
 sg13g2_decap_8 FILLER_51_770 ();
 sg13g2_decap_8 FILLER_51_777 ();
 sg13g2_decap_8 FILLER_51_784 ();
 sg13g2_decap_8 FILLER_51_791 ();
 sg13g2_decap_8 FILLER_51_798 ();
 sg13g2_decap_8 FILLER_51_805 ();
 sg13g2_decap_8 FILLER_51_812 ();
 sg13g2_decap_8 FILLER_51_819 ();
 sg13g2_decap_8 FILLER_51_826 ();
 sg13g2_decap_8 FILLER_51_833 ();
 sg13g2_fill_1 FILLER_51_840 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_168 ();
 sg13g2_decap_8 FILLER_52_175 ();
 sg13g2_decap_8 FILLER_52_182 ();
 sg13g2_decap_8 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_196 ();
 sg13g2_decap_8 FILLER_52_203 ();
 sg13g2_decap_8 FILLER_52_210 ();
 sg13g2_decap_8 FILLER_52_217 ();
 sg13g2_decap_8 FILLER_52_224 ();
 sg13g2_decap_8 FILLER_52_231 ();
 sg13g2_decap_8 FILLER_52_238 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_decap_8 FILLER_52_252 ();
 sg13g2_decap_8 FILLER_52_259 ();
 sg13g2_decap_8 FILLER_52_266 ();
 sg13g2_decap_8 FILLER_52_273 ();
 sg13g2_decap_8 FILLER_52_280 ();
 sg13g2_decap_8 FILLER_52_287 ();
 sg13g2_decap_8 FILLER_52_294 ();
 sg13g2_decap_8 FILLER_52_301 ();
 sg13g2_decap_8 FILLER_52_308 ();
 sg13g2_decap_8 FILLER_52_315 ();
 sg13g2_decap_8 FILLER_52_322 ();
 sg13g2_decap_8 FILLER_52_329 ();
 sg13g2_decap_8 FILLER_52_336 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_decap_8 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_decap_8 FILLER_52_364 ();
 sg13g2_decap_8 FILLER_52_371 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_413 ();
 sg13g2_decap_8 FILLER_52_420 ();
 sg13g2_decap_8 FILLER_52_427 ();
 sg13g2_decap_8 FILLER_52_434 ();
 sg13g2_decap_8 FILLER_52_441 ();
 sg13g2_decap_8 FILLER_52_448 ();
 sg13g2_decap_8 FILLER_52_455 ();
 sg13g2_decap_8 FILLER_52_462 ();
 sg13g2_decap_8 FILLER_52_469 ();
 sg13g2_decap_8 FILLER_52_476 ();
 sg13g2_decap_8 FILLER_52_483 ();
 sg13g2_decap_8 FILLER_52_490 ();
 sg13g2_decap_8 FILLER_52_497 ();
 sg13g2_decap_8 FILLER_52_504 ();
 sg13g2_decap_8 FILLER_52_511 ();
 sg13g2_decap_8 FILLER_52_518 ();
 sg13g2_decap_8 FILLER_52_525 ();
 sg13g2_decap_8 FILLER_52_532 ();
 sg13g2_decap_8 FILLER_52_539 ();
 sg13g2_decap_8 FILLER_52_546 ();
 sg13g2_decap_8 FILLER_52_553 ();
 sg13g2_decap_8 FILLER_52_560 ();
 sg13g2_decap_8 FILLER_52_567 ();
 sg13g2_decap_8 FILLER_52_574 ();
 sg13g2_decap_8 FILLER_52_581 ();
 sg13g2_decap_8 FILLER_52_588 ();
 sg13g2_decap_8 FILLER_52_595 ();
 sg13g2_decap_8 FILLER_52_602 ();
 sg13g2_decap_8 FILLER_52_609 ();
 sg13g2_decap_8 FILLER_52_616 ();
 sg13g2_decap_8 FILLER_52_623 ();
 sg13g2_decap_8 FILLER_52_630 ();
 sg13g2_decap_8 FILLER_52_637 ();
 sg13g2_decap_8 FILLER_52_644 ();
 sg13g2_decap_8 FILLER_52_651 ();
 sg13g2_decap_8 FILLER_52_658 ();
 sg13g2_decap_8 FILLER_52_665 ();
 sg13g2_decap_8 FILLER_52_672 ();
 sg13g2_decap_8 FILLER_52_679 ();
 sg13g2_decap_8 FILLER_52_686 ();
 sg13g2_decap_8 FILLER_52_693 ();
 sg13g2_decap_8 FILLER_52_700 ();
 sg13g2_decap_8 FILLER_52_707 ();
 sg13g2_decap_8 FILLER_52_714 ();
 sg13g2_decap_8 FILLER_52_721 ();
 sg13g2_decap_8 FILLER_52_728 ();
 sg13g2_decap_8 FILLER_52_735 ();
 sg13g2_decap_8 FILLER_52_742 ();
 sg13g2_decap_8 FILLER_52_749 ();
 sg13g2_decap_8 FILLER_52_756 ();
 sg13g2_decap_8 FILLER_52_763 ();
 sg13g2_decap_8 FILLER_52_770 ();
 sg13g2_decap_8 FILLER_52_777 ();
 sg13g2_decap_8 FILLER_52_784 ();
 sg13g2_decap_8 FILLER_52_791 ();
 sg13g2_decap_8 FILLER_52_798 ();
 sg13g2_decap_8 FILLER_52_805 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_decap_8 FILLER_52_833 ();
 sg13g2_fill_1 FILLER_52_840 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_decap_8 FILLER_53_161 ();
 sg13g2_decap_8 FILLER_53_168 ();
 sg13g2_decap_8 FILLER_53_175 ();
 sg13g2_decap_8 FILLER_53_182 ();
 sg13g2_decap_8 FILLER_53_189 ();
 sg13g2_decap_8 FILLER_53_196 ();
 sg13g2_decap_8 FILLER_53_203 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_224 ();
 sg13g2_decap_8 FILLER_53_231 ();
 sg13g2_decap_8 FILLER_53_238 ();
 sg13g2_decap_8 FILLER_53_245 ();
 sg13g2_decap_8 FILLER_53_252 ();
 sg13g2_decap_8 FILLER_53_259 ();
 sg13g2_decap_8 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_273 ();
 sg13g2_decap_8 FILLER_53_280 ();
 sg13g2_decap_8 FILLER_53_287 ();
 sg13g2_decap_8 FILLER_53_294 ();
 sg13g2_decap_8 FILLER_53_301 ();
 sg13g2_decap_8 FILLER_53_308 ();
 sg13g2_decap_8 FILLER_53_315 ();
 sg13g2_decap_8 FILLER_53_322 ();
 sg13g2_decap_8 FILLER_53_329 ();
 sg13g2_decap_8 FILLER_53_336 ();
 sg13g2_decap_8 FILLER_53_343 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_decap_8 FILLER_53_357 ();
 sg13g2_decap_8 FILLER_53_364 ();
 sg13g2_decap_8 FILLER_53_371 ();
 sg13g2_decap_8 FILLER_53_378 ();
 sg13g2_decap_8 FILLER_53_385 ();
 sg13g2_decap_8 FILLER_53_392 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_decap_8 FILLER_53_406 ();
 sg13g2_decap_8 FILLER_53_413 ();
 sg13g2_decap_8 FILLER_53_420 ();
 sg13g2_decap_8 FILLER_53_427 ();
 sg13g2_decap_8 FILLER_53_434 ();
 sg13g2_decap_8 FILLER_53_441 ();
 sg13g2_decap_8 FILLER_53_448 ();
 sg13g2_decap_8 FILLER_53_455 ();
 sg13g2_decap_8 FILLER_53_462 ();
 sg13g2_decap_8 FILLER_53_469 ();
 sg13g2_decap_8 FILLER_53_476 ();
 sg13g2_decap_8 FILLER_53_483 ();
 sg13g2_decap_8 FILLER_53_490 ();
 sg13g2_decap_8 FILLER_53_497 ();
 sg13g2_decap_8 FILLER_53_504 ();
 sg13g2_decap_8 FILLER_53_511 ();
 sg13g2_decap_8 FILLER_53_518 ();
 sg13g2_decap_8 FILLER_53_525 ();
 sg13g2_decap_8 FILLER_53_532 ();
 sg13g2_decap_8 FILLER_53_539 ();
 sg13g2_decap_8 FILLER_53_546 ();
 sg13g2_decap_8 FILLER_53_553 ();
 sg13g2_decap_8 FILLER_53_560 ();
 sg13g2_decap_8 FILLER_53_567 ();
 sg13g2_decap_8 FILLER_53_574 ();
 sg13g2_decap_8 FILLER_53_581 ();
 sg13g2_decap_8 FILLER_53_588 ();
 sg13g2_decap_8 FILLER_53_595 ();
 sg13g2_decap_8 FILLER_53_602 ();
 sg13g2_decap_8 FILLER_53_609 ();
 sg13g2_decap_8 FILLER_53_616 ();
 sg13g2_decap_8 FILLER_53_623 ();
 sg13g2_decap_8 FILLER_53_630 ();
 sg13g2_decap_8 FILLER_53_637 ();
 sg13g2_decap_8 FILLER_53_644 ();
 sg13g2_decap_8 FILLER_53_651 ();
 sg13g2_decap_8 FILLER_53_658 ();
 sg13g2_decap_8 FILLER_53_665 ();
 sg13g2_decap_8 FILLER_53_672 ();
 sg13g2_decap_8 FILLER_53_679 ();
 sg13g2_decap_8 FILLER_53_686 ();
 sg13g2_decap_8 FILLER_53_693 ();
 sg13g2_decap_8 FILLER_53_700 ();
 sg13g2_decap_8 FILLER_53_707 ();
 sg13g2_decap_8 FILLER_53_714 ();
 sg13g2_decap_8 FILLER_53_721 ();
 sg13g2_decap_8 FILLER_53_728 ();
 sg13g2_decap_8 FILLER_53_735 ();
 sg13g2_decap_8 FILLER_53_742 ();
 sg13g2_decap_8 FILLER_53_749 ();
 sg13g2_decap_8 FILLER_53_756 ();
 sg13g2_decap_8 FILLER_53_763 ();
 sg13g2_decap_8 FILLER_53_770 ();
 sg13g2_decap_8 FILLER_53_777 ();
 sg13g2_decap_8 FILLER_53_784 ();
 sg13g2_decap_8 FILLER_53_791 ();
 sg13g2_decap_8 FILLER_53_798 ();
 sg13g2_decap_8 FILLER_53_805 ();
 sg13g2_decap_8 FILLER_53_812 ();
 sg13g2_decap_8 FILLER_53_819 ();
 sg13g2_decap_8 FILLER_53_826 ();
 sg13g2_decap_8 FILLER_53_833 ();
 sg13g2_fill_1 FILLER_53_840 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_8 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_decap_8 FILLER_54_168 ();
 sg13g2_decap_8 FILLER_54_175 ();
 sg13g2_decap_8 FILLER_54_182 ();
 sg13g2_decap_8 FILLER_54_189 ();
 sg13g2_decap_8 FILLER_54_196 ();
 sg13g2_decap_8 FILLER_54_203 ();
 sg13g2_decap_8 FILLER_54_210 ();
 sg13g2_decap_8 FILLER_54_217 ();
 sg13g2_decap_8 FILLER_54_224 ();
 sg13g2_decap_8 FILLER_54_231 ();
 sg13g2_decap_8 FILLER_54_238 ();
 sg13g2_decap_8 FILLER_54_245 ();
 sg13g2_decap_8 FILLER_54_252 ();
 sg13g2_decap_8 FILLER_54_259 ();
 sg13g2_decap_8 FILLER_54_266 ();
 sg13g2_decap_8 FILLER_54_273 ();
 sg13g2_decap_8 FILLER_54_280 ();
 sg13g2_decap_8 FILLER_54_287 ();
 sg13g2_decap_8 FILLER_54_294 ();
 sg13g2_decap_8 FILLER_54_301 ();
 sg13g2_decap_8 FILLER_54_308 ();
 sg13g2_decap_8 FILLER_54_315 ();
 sg13g2_decap_8 FILLER_54_322 ();
 sg13g2_decap_8 FILLER_54_329 ();
 sg13g2_decap_8 FILLER_54_336 ();
 sg13g2_decap_8 FILLER_54_343 ();
 sg13g2_decap_8 FILLER_54_350 ();
 sg13g2_decap_8 FILLER_54_357 ();
 sg13g2_decap_8 FILLER_54_364 ();
 sg13g2_decap_8 FILLER_54_371 ();
 sg13g2_decap_8 FILLER_54_378 ();
 sg13g2_decap_8 FILLER_54_385 ();
 sg13g2_decap_8 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_399 ();
 sg13g2_decap_8 FILLER_54_406 ();
 sg13g2_decap_8 FILLER_54_413 ();
 sg13g2_decap_8 FILLER_54_420 ();
 sg13g2_decap_8 FILLER_54_427 ();
 sg13g2_decap_8 FILLER_54_434 ();
 sg13g2_decap_8 FILLER_54_441 ();
 sg13g2_decap_8 FILLER_54_448 ();
 sg13g2_decap_8 FILLER_54_455 ();
 sg13g2_decap_8 FILLER_54_462 ();
 sg13g2_decap_8 FILLER_54_469 ();
 sg13g2_decap_8 FILLER_54_476 ();
 sg13g2_decap_8 FILLER_54_483 ();
 sg13g2_decap_8 FILLER_54_490 ();
 sg13g2_decap_8 FILLER_54_497 ();
 sg13g2_decap_8 FILLER_54_504 ();
 sg13g2_decap_8 FILLER_54_511 ();
 sg13g2_decap_8 FILLER_54_518 ();
 sg13g2_decap_8 FILLER_54_525 ();
 sg13g2_decap_8 FILLER_54_532 ();
 sg13g2_decap_8 FILLER_54_539 ();
 sg13g2_decap_8 FILLER_54_546 ();
 sg13g2_decap_8 FILLER_54_553 ();
 sg13g2_decap_8 FILLER_54_560 ();
 sg13g2_decap_8 FILLER_54_567 ();
 sg13g2_decap_8 FILLER_54_574 ();
 sg13g2_decap_8 FILLER_54_581 ();
 sg13g2_decap_8 FILLER_54_588 ();
 sg13g2_decap_8 FILLER_54_595 ();
 sg13g2_decap_8 FILLER_54_602 ();
 sg13g2_decap_8 FILLER_54_609 ();
 sg13g2_decap_8 FILLER_54_616 ();
 sg13g2_decap_8 FILLER_54_623 ();
 sg13g2_decap_8 FILLER_54_630 ();
 sg13g2_decap_8 FILLER_54_637 ();
 sg13g2_decap_8 FILLER_54_644 ();
 sg13g2_decap_8 FILLER_54_651 ();
 sg13g2_decap_8 FILLER_54_658 ();
 sg13g2_decap_8 FILLER_54_665 ();
 sg13g2_decap_8 FILLER_54_672 ();
 sg13g2_decap_8 FILLER_54_679 ();
 sg13g2_decap_8 FILLER_54_686 ();
 sg13g2_decap_8 FILLER_54_693 ();
 sg13g2_decap_8 FILLER_54_700 ();
 sg13g2_decap_8 FILLER_54_707 ();
 sg13g2_decap_8 FILLER_54_714 ();
 sg13g2_decap_8 FILLER_54_721 ();
 sg13g2_decap_8 FILLER_54_728 ();
 sg13g2_decap_8 FILLER_54_735 ();
 sg13g2_decap_8 FILLER_54_742 ();
 sg13g2_decap_8 FILLER_54_749 ();
 sg13g2_decap_8 FILLER_54_756 ();
 sg13g2_decap_8 FILLER_54_763 ();
 sg13g2_decap_8 FILLER_54_770 ();
 sg13g2_decap_8 FILLER_54_777 ();
 sg13g2_decap_8 FILLER_54_784 ();
 sg13g2_decap_8 FILLER_54_791 ();
 sg13g2_decap_8 FILLER_54_798 ();
 sg13g2_decap_8 FILLER_54_805 ();
 sg13g2_decap_8 FILLER_54_812 ();
 sg13g2_decap_8 FILLER_54_819 ();
 sg13g2_decap_8 FILLER_54_826 ();
 sg13g2_decap_8 FILLER_54_833 ();
 sg13g2_fill_1 FILLER_54_840 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_168 ();
 sg13g2_decap_8 FILLER_55_175 ();
 sg13g2_decap_8 FILLER_55_182 ();
 sg13g2_decap_8 FILLER_55_189 ();
 sg13g2_decap_8 FILLER_55_196 ();
 sg13g2_decap_8 FILLER_55_203 ();
 sg13g2_decap_8 FILLER_55_210 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_decap_8 FILLER_55_224 ();
 sg13g2_decap_8 FILLER_55_231 ();
 sg13g2_decap_8 FILLER_55_238 ();
 sg13g2_decap_8 FILLER_55_245 ();
 sg13g2_decap_8 FILLER_55_252 ();
 sg13g2_decap_8 FILLER_55_259 ();
 sg13g2_decap_8 FILLER_55_266 ();
 sg13g2_decap_8 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_8 FILLER_55_287 ();
 sg13g2_decap_8 FILLER_55_294 ();
 sg13g2_decap_8 FILLER_55_301 ();
 sg13g2_decap_8 FILLER_55_308 ();
 sg13g2_decap_8 FILLER_55_315 ();
 sg13g2_decap_8 FILLER_55_322 ();
 sg13g2_decap_8 FILLER_55_329 ();
 sg13g2_decap_8 FILLER_55_336 ();
 sg13g2_decap_8 FILLER_55_343 ();
 sg13g2_decap_8 FILLER_55_350 ();
 sg13g2_decap_8 FILLER_55_357 ();
 sg13g2_decap_8 FILLER_55_364 ();
 sg13g2_decap_8 FILLER_55_371 ();
 sg13g2_decap_8 FILLER_55_378 ();
 sg13g2_decap_8 FILLER_55_385 ();
 sg13g2_decap_8 FILLER_55_392 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_decap_8 FILLER_55_406 ();
 sg13g2_decap_8 FILLER_55_413 ();
 sg13g2_decap_8 FILLER_55_420 ();
 sg13g2_decap_8 FILLER_55_427 ();
 sg13g2_decap_8 FILLER_55_434 ();
 sg13g2_decap_8 FILLER_55_441 ();
 sg13g2_decap_8 FILLER_55_448 ();
 sg13g2_decap_8 FILLER_55_455 ();
 sg13g2_decap_8 FILLER_55_462 ();
 sg13g2_decap_8 FILLER_55_469 ();
 sg13g2_decap_8 FILLER_55_476 ();
 sg13g2_decap_8 FILLER_55_483 ();
 sg13g2_decap_8 FILLER_55_490 ();
 sg13g2_decap_8 FILLER_55_497 ();
 sg13g2_decap_8 FILLER_55_504 ();
 sg13g2_decap_8 FILLER_55_511 ();
 sg13g2_decap_8 FILLER_55_518 ();
 sg13g2_decap_8 FILLER_55_525 ();
 sg13g2_decap_8 FILLER_55_532 ();
 sg13g2_decap_8 FILLER_55_539 ();
 sg13g2_decap_8 FILLER_55_546 ();
 sg13g2_decap_8 FILLER_55_553 ();
 sg13g2_decap_8 FILLER_55_560 ();
 sg13g2_decap_8 FILLER_55_567 ();
 sg13g2_decap_8 FILLER_55_574 ();
 sg13g2_decap_8 FILLER_55_581 ();
 sg13g2_decap_8 FILLER_55_588 ();
 sg13g2_decap_8 FILLER_55_595 ();
 sg13g2_decap_8 FILLER_55_602 ();
 sg13g2_decap_8 FILLER_55_609 ();
 sg13g2_decap_8 FILLER_55_616 ();
 sg13g2_decap_8 FILLER_55_623 ();
 sg13g2_decap_8 FILLER_55_630 ();
 sg13g2_decap_8 FILLER_55_637 ();
 sg13g2_decap_8 FILLER_55_644 ();
 sg13g2_decap_8 FILLER_55_651 ();
 sg13g2_decap_8 FILLER_55_658 ();
 sg13g2_decap_8 FILLER_55_665 ();
 sg13g2_decap_8 FILLER_55_672 ();
 sg13g2_decap_8 FILLER_55_679 ();
 sg13g2_decap_8 FILLER_55_686 ();
 sg13g2_decap_8 FILLER_55_693 ();
 sg13g2_decap_8 FILLER_55_700 ();
 sg13g2_decap_8 FILLER_55_707 ();
 sg13g2_decap_8 FILLER_55_714 ();
 sg13g2_decap_8 FILLER_55_721 ();
 sg13g2_decap_8 FILLER_55_728 ();
 sg13g2_decap_8 FILLER_55_735 ();
 sg13g2_decap_8 FILLER_55_742 ();
 sg13g2_decap_8 FILLER_55_749 ();
 sg13g2_decap_8 FILLER_55_756 ();
 sg13g2_decap_8 FILLER_55_763 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_decap_8 FILLER_55_777 ();
 sg13g2_decap_8 FILLER_55_784 ();
 sg13g2_decap_8 FILLER_55_791 ();
 sg13g2_decap_8 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_805 ();
 sg13g2_decap_8 FILLER_55_812 ();
 sg13g2_decap_8 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_826 ();
 sg13g2_decap_8 FILLER_55_833 ();
 sg13g2_fill_1 FILLER_55_840 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_decap_8 FILLER_56_182 ();
 sg13g2_decap_8 FILLER_56_189 ();
 sg13g2_decap_8 FILLER_56_196 ();
 sg13g2_decap_8 FILLER_56_203 ();
 sg13g2_decap_8 FILLER_56_210 ();
 sg13g2_decap_8 FILLER_56_217 ();
 sg13g2_decap_8 FILLER_56_224 ();
 sg13g2_decap_8 FILLER_56_231 ();
 sg13g2_decap_8 FILLER_56_238 ();
 sg13g2_decap_8 FILLER_56_245 ();
 sg13g2_decap_8 FILLER_56_252 ();
 sg13g2_decap_8 FILLER_56_259 ();
 sg13g2_decap_8 FILLER_56_266 ();
 sg13g2_decap_8 FILLER_56_273 ();
 sg13g2_decap_8 FILLER_56_280 ();
 sg13g2_decap_8 FILLER_56_287 ();
 sg13g2_decap_8 FILLER_56_294 ();
 sg13g2_decap_8 FILLER_56_301 ();
 sg13g2_decap_8 FILLER_56_308 ();
 sg13g2_decap_8 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_322 ();
 sg13g2_decap_8 FILLER_56_329 ();
 sg13g2_decap_8 FILLER_56_336 ();
 sg13g2_decap_8 FILLER_56_343 ();
 sg13g2_decap_8 FILLER_56_350 ();
 sg13g2_decap_8 FILLER_56_357 ();
 sg13g2_decap_8 FILLER_56_364 ();
 sg13g2_decap_8 FILLER_56_371 ();
 sg13g2_decap_8 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_385 ();
 sg13g2_decap_8 FILLER_56_392 ();
 sg13g2_decap_8 FILLER_56_399 ();
 sg13g2_decap_8 FILLER_56_406 ();
 sg13g2_decap_8 FILLER_56_413 ();
 sg13g2_decap_8 FILLER_56_420 ();
 sg13g2_decap_8 FILLER_56_427 ();
 sg13g2_decap_8 FILLER_56_434 ();
 sg13g2_decap_8 FILLER_56_441 ();
 sg13g2_decap_8 FILLER_56_448 ();
 sg13g2_decap_8 FILLER_56_455 ();
 sg13g2_decap_8 FILLER_56_462 ();
 sg13g2_decap_8 FILLER_56_469 ();
 sg13g2_decap_8 FILLER_56_476 ();
 sg13g2_decap_8 FILLER_56_483 ();
 sg13g2_decap_8 FILLER_56_490 ();
 sg13g2_decap_8 FILLER_56_497 ();
 sg13g2_decap_8 FILLER_56_504 ();
 sg13g2_decap_8 FILLER_56_511 ();
 sg13g2_decap_8 FILLER_56_518 ();
 sg13g2_decap_8 FILLER_56_525 ();
 sg13g2_decap_8 FILLER_56_532 ();
 sg13g2_decap_8 FILLER_56_539 ();
 sg13g2_decap_8 FILLER_56_546 ();
 sg13g2_decap_8 FILLER_56_553 ();
 sg13g2_decap_8 FILLER_56_560 ();
 sg13g2_decap_8 FILLER_56_567 ();
 sg13g2_decap_8 FILLER_56_574 ();
 sg13g2_decap_8 FILLER_56_581 ();
 sg13g2_decap_8 FILLER_56_588 ();
 sg13g2_decap_8 FILLER_56_595 ();
 sg13g2_decap_8 FILLER_56_602 ();
 sg13g2_decap_8 FILLER_56_609 ();
 sg13g2_decap_8 FILLER_56_616 ();
 sg13g2_decap_8 FILLER_56_623 ();
 sg13g2_decap_8 FILLER_56_630 ();
 sg13g2_decap_8 FILLER_56_637 ();
 sg13g2_decap_8 FILLER_56_644 ();
 sg13g2_decap_8 FILLER_56_651 ();
 sg13g2_decap_8 FILLER_56_658 ();
 sg13g2_decap_8 FILLER_56_665 ();
 sg13g2_decap_8 FILLER_56_672 ();
 sg13g2_decap_8 FILLER_56_679 ();
 sg13g2_decap_8 FILLER_56_686 ();
 sg13g2_decap_8 FILLER_56_693 ();
 sg13g2_decap_8 FILLER_56_700 ();
 sg13g2_decap_8 FILLER_56_707 ();
 sg13g2_decap_8 FILLER_56_714 ();
 sg13g2_decap_8 FILLER_56_721 ();
 sg13g2_decap_8 FILLER_56_728 ();
 sg13g2_decap_8 FILLER_56_735 ();
 sg13g2_decap_8 FILLER_56_742 ();
 sg13g2_decap_8 FILLER_56_749 ();
 sg13g2_decap_8 FILLER_56_756 ();
 sg13g2_decap_8 FILLER_56_763 ();
 sg13g2_decap_8 FILLER_56_770 ();
 sg13g2_decap_8 FILLER_56_777 ();
 sg13g2_decap_8 FILLER_56_784 ();
 sg13g2_decap_8 FILLER_56_791 ();
 sg13g2_decap_8 FILLER_56_798 ();
 sg13g2_decap_8 FILLER_56_805 ();
 sg13g2_decap_8 FILLER_56_812 ();
 sg13g2_decap_8 FILLER_56_819 ();
 sg13g2_decap_8 FILLER_56_826 ();
 sg13g2_decap_8 FILLER_56_833 ();
 sg13g2_fill_1 FILLER_56_840 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_decap_8 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_189 ();
 sg13g2_decap_8 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_231 ();
 sg13g2_decap_8 FILLER_57_238 ();
 sg13g2_decap_8 FILLER_57_245 ();
 sg13g2_decap_8 FILLER_57_252 ();
 sg13g2_decap_8 FILLER_57_259 ();
 sg13g2_decap_8 FILLER_57_266 ();
 sg13g2_decap_8 FILLER_57_273 ();
 sg13g2_decap_8 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_287 ();
 sg13g2_decap_8 FILLER_57_294 ();
 sg13g2_decap_8 FILLER_57_301 ();
 sg13g2_decap_8 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_315 ();
 sg13g2_decap_8 FILLER_57_322 ();
 sg13g2_decap_8 FILLER_57_329 ();
 sg13g2_decap_8 FILLER_57_336 ();
 sg13g2_decap_8 FILLER_57_343 ();
 sg13g2_decap_8 FILLER_57_350 ();
 sg13g2_decap_8 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_364 ();
 sg13g2_decap_8 FILLER_57_371 ();
 sg13g2_decap_8 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_385 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_57_406 ();
 sg13g2_decap_8 FILLER_57_413 ();
 sg13g2_decap_8 FILLER_57_420 ();
 sg13g2_decap_8 FILLER_57_427 ();
 sg13g2_decap_8 FILLER_57_434 ();
 sg13g2_decap_8 FILLER_57_441 ();
 sg13g2_decap_8 FILLER_57_448 ();
 sg13g2_decap_8 FILLER_57_455 ();
 sg13g2_decap_8 FILLER_57_462 ();
 sg13g2_decap_8 FILLER_57_469 ();
 sg13g2_decap_8 FILLER_57_476 ();
 sg13g2_decap_8 FILLER_57_483 ();
 sg13g2_decap_8 FILLER_57_490 ();
 sg13g2_decap_8 FILLER_57_497 ();
 sg13g2_decap_8 FILLER_57_504 ();
 sg13g2_decap_8 FILLER_57_511 ();
 sg13g2_decap_8 FILLER_57_518 ();
 sg13g2_decap_8 FILLER_57_525 ();
 sg13g2_decap_8 FILLER_57_532 ();
 sg13g2_decap_8 FILLER_57_539 ();
 sg13g2_decap_8 FILLER_57_546 ();
 sg13g2_decap_8 FILLER_57_553 ();
 sg13g2_decap_8 FILLER_57_560 ();
 sg13g2_decap_8 FILLER_57_567 ();
 sg13g2_decap_8 FILLER_57_574 ();
 sg13g2_decap_8 FILLER_57_581 ();
 sg13g2_decap_8 FILLER_57_588 ();
 sg13g2_decap_8 FILLER_57_595 ();
 sg13g2_decap_8 FILLER_57_602 ();
 sg13g2_decap_8 FILLER_57_609 ();
 sg13g2_decap_8 FILLER_57_616 ();
 sg13g2_decap_8 FILLER_57_623 ();
 sg13g2_decap_8 FILLER_57_630 ();
 sg13g2_decap_8 FILLER_57_637 ();
 sg13g2_decap_8 FILLER_57_644 ();
 sg13g2_decap_8 FILLER_57_651 ();
 sg13g2_decap_8 FILLER_57_658 ();
 sg13g2_decap_8 FILLER_57_665 ();
 sg13g2_decap_8 FILLER_57_672 ();
 sg13g2_decap_8 FILLER_57_679 ();
 sg13g2_decap_8 FILLER_57_686 ();
 sg13g2_decap_8 FILLER_57_693 ();
 sg13g2_decap_8 FILLER_57_700 ();
 sg13g2_decap_8 FILLER_57_707 ();
 sg13g2_decap_8 FILLER_57_714 ();
 sg13g2_decap_8 FILLER_57_721 ();
 sg13g2_decap_8 FILLER_57_728 ();
 sg13g2_decap_8 FILLER_57_735 ();
 sg13g2_decap_8 FILLER_57_742 ();
 sg13g2_decap_8 FILLER_57_749 ();
 sg13g2_decap_8 FILLER_57_756 ();
 sg13g2_decap_8 FILLER_57_763 ();
 sg13g2_decap_8 FILLER_57_770 ();
 sg13g2_decap_8 FILLER_57_777 ();
 sg13g2_decap_8 FILLER_57_784 ();
 sg13g2_decap_8 FILLER_57_791 ();
 sg13g2_decap_8 FILLER_57_798 ();
 sg13g2_decap_8 FILLER_57_805 ();
 sg13g2_decap_8 FILLER_57_812 ();
 sg13g2_decap_8 FILLER_57_819 ();
 sg13g2_decap_8 FILLER_57_826 ();
 sg13g2_decap_8 FILLER_57_833 ();
 sg13g2_fill_1 FILLER_57_840 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_210 ();
 sg13g2_decap_8 FILLER_58_217 ();
 sg13g2_decap_8 FILLER_58_224 ();
 sg13g2_decap_8 FILLER_58_231 ();
 sg13g2_decap_8 FILLER_58_238 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_decap_8 FILLER_58_252 ();
 sg13g2_decap_8 FILLER_58_259 ();
 sg13g2_decap_8 FILLER_58_266 ();
 sg13g2_decap_8 FILLER_58_273 ();
 sg13g2_decap_8 FILLER_58_280 ();
 sg13g2_decap_8 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_8 FILLER_58_301 ();
 sg13g2_decap_8 FILLER_58_308 ();
 sg13g2_decap_8 FILLER_58_315 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_329 ();
 sg13g2_decap_8 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_343 ();
 sg13g2_decap_8 FILLER_58_350 ();
 sg13g2_decap_8 FILLER_58_357 ();
 sg13g2_decap_8 FILLER_58_364 ();
 sg13g2_decap_8 FILLER_58_371 ();
 sg13g2_decap_8 FILLER_58_378 ();
 sg13g2_decap_8 FILLER_58_385 ();
 sg13g2_decap_8 FILLER_58_392 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_decap_8 FILLER_58_406 ();
 sg13g2_decap_8 FILLER_58_413 ();
 sg13g2_decap_8 FILLER_58_420 ();
 sg13g2_decap_8 FILLER_58_427 ();
 sg13g2_decap_8 FILLER_58_434 ();
 sg13g2_decap_8 FILLER_58_441 ();
 sg13g2_decap_8 FILLER_58_448 ();
 sg13g2_decap_8 FILLER_58_455 ();
 sg13g2_decap_8 FILLER_58_462 ();
 sg13g2_decap_8 FILLER_58_469 ();
 sg13g2_decap_8 FILLER_58_476 ();
 sg13g2_decap_8 FILLER_58_483 ();
 sg13g2_decap_8 FILLER_58_490 ();
 sg13g2_decap_8 FILLER_58_497 ();
 sg13g2_decap_8 FILLER_58_504 ();
 sg13g2_decap_8 FILLER_58_511 ();
 sg13g2_decap_8 FILLER_58_518 ();
 sg13g2_decap_8 FILLER_58_525 ();
 sg13g2_decap_8 FILLER_58_532 ();
 sg13g2_decap_8 FILLER_58_539 ();
 sg13g2_decap_8 FILLER_58_546 ();
 sg13g2_decap_8 FILLER_58_553 ();
 sg13g2_decap_8 FILLER_58_560 ();
 sg13g2_decap_8 FILLER_58_567 ();
 sg13g2_decap_8 FILLER_58_574 ();
 sg13g2_decap_8 FILLER_58_581 ();
 sg13g2_decap_8 FILLER_58_588 ();
 sg13g2_decap_8 FILLER_58_595 ();
 sg13g2_decap_8 FILLER_58_602 ();
 sg13g2_decap_8 FILLER_58_609 ();
 sg13g2_decap_8 FILLER_58_616 ();
 sg13g2_decap_8 FILLER_58_623 ();
 sg13g2_decap_8 FILLER_58_630 ();
 sg13g2_decap_8 FILLER_58_637 ();
 sg13g2_decap_8 FILLER_58_644 ();
 sg13g2_decap_8 FILLER_58_651 ();
 sg13g2_decap_8 FILLER_58_658 ();
 sg13g2_decap_8 FILLER_58_665 ();
 sg13g2_decap_8 FILLER_58_672 ();
 sg13g2_decap_8 FILLER_58_679 ();
 sg13g2_decap_8 FILLER_58_686 ();
 sg13g2_decap_8 FILLER_58_693 ();
 sg13g2_decap_8 FILLER_58_700 ();
 sg13g2_decap_8 FILLER_58_707 ();
 sg13g2_decap_8 FILLER_58_714 ();
 sg13g2_decap_8 FILLER_58_721 ();
 sg13g2_decap_8 FILLER_58_728 ();
 sg13g2_decap_8 FILLER_58_735 ();
 sg13g2_decap_8 FILLER_58_742 ();
 sg13g2_decap_8 FILLER_58_749 ();
 sg13g2_decap_8 FILLER_58_756 ();
 sg13g2_decap_8 FILLER_58_763 ();
 sg13g2_decap_8 FILLER_58_770 ();
 sg13g2_decap_8 FILLER_58_777 ();
 sg13g2_decap_8 FILLER_58_784 ();
 sg13g2_decap_8 FILLER_58_791 ();
 sg13g2_decap_8 FILLER_58_798 ();
 sg13g2_decap_8 FILLER_58_805 ();
 sg13g2_decap_8 FILLER_58_812 ();
 sg13g2_decap_8 FILLER_58_819 ();
 sg13g2_decap_8 FILLER_58_826 ();
 sg13g2_decap_8 FILLER_58_833 ();
 sg13g2_fill_1 FILLER_58_840 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_decap_8 FILLER_59_175 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_decap_8 FILLER_59_203 ();
 sg13g2_decap_8 FILLER_59_210 ();
 sg13g2_decap_8 FILLER_59_217 ();
 sg13g2_decap_8 FILLER_59_224 ();
 sg13g2_decap_8 FILLER_59_231 ();
 sg13g2_decap_8 FILLER_59_238 ();
 sg13g2_decap_8 FILLER_59_245 ();
 sg13g2_decap_8 FILLER_59_252 ();
 sg13g2_decap_8 FILLER_59_259 ();
 sg13g2_decap_8 FILLER_59_266 ();
 sg13g2_decap_8 FILLER_59_273 ();
 sg13g2_decap_8 FILLER_59_280 ();
 sg13g2_decap_8 FILLER_59_287 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_decap_8 FILLER_59_301 ();
 sg13g2_decap_8 FILLER_59_308 ();
 sg13g2_decap_8 FILLER_59_315 ();
 sg13g2_decap_8 FILLER_59_322 ();
 sg13g2_decap_8 FILLER_59_329 ();
 sg13g2_decap_8 FILLER_59_336 ();
 sg13g2_decap_8 FILLER_59_343 ();
 sg13g2_decap_8 FILLER_59_350 ();
 sg13g2_decap_8 FILLER_59_357 ();
 sg13g2_decap_8 FILLER_59_364 ();
 sg13g2_decap_8 FILLER_59_371 ();
 sg13g2_decap_8 FILLER_59_378 ();
 sg13g2_decap_8 FILLER_59_385 ();
 sg13g2_decap_8 FILLER_59_392 ();
 sg13g2_decap_8 FILLER_59_399 ();
 sg13g2_decap_8 FILLER_59_406 ();
 sg13g2_decap_8 FILLER_59_413 ();
 sg13g2_decap_8 FILLER_59_420 ();
 sg13g2_decap_8 FILLER_59_427 ();
 sg13g2_decap_8 FILLER_59_434 ();
 sg13g2_decap_8 FILLER_59_441 ();
 sg13g2_decap_8 FILLER_59_448 ();
 sg13g2_decap_8 FILLER_59_455 ();
 sg13g2_decap_8 FILLER_59_462 ();
 sg13g2_decap_8 FILLER_59_469 ();
 sg13g2_decap_8 FILLER_59_476 ();
 sg13g2_decap_8 FILLER_59_483 ();
 sg13g2_decap_8 FILLER_59_490 ();
 sg13g2_decap_8 FILLER_59_497 ();
 sg13g2_decap_8 FILLER_59_504 ();
 sg13g2_decap_8 FILLER_59_511 ();
 sg13g2_decap_8 FILLER_59_518 ();
 sg13g2_decap_8 FILLER_59_525 ();
 sg13g2_decap_8 FILLER_59_532 ();
 sg13g2_decap_8 FILLER_59_539 ();
 sg13g2_decap_8 FILLER_59_546 ();
 sg13g2_decap_8 FILLER_59_553 ();
 sg13g2_decap_8 FILLER_59_560 ();
 sg13g2_decap_8 FILLER_59_567 ();
 sg13g2_decap_8 FILLER_59_574 ();
 sg13g2_decap_8 FILLER_59_581 ();
 sg13g2_decap_8 FILLER_59_588 ();
 sg13g2_decap_8 FILLER_59_595 ();
 sg13g2_decap_8 FILLER_59_602 ();
 sg13g2_decap_8 FILLER_59_609 ();
 sg13g2_decap_8 FILLER_59_616 ();
 sg13g2_decap_8 FILLER_59_623 ();
 sg13g2_decap_8 FILLER_59_630 ();
 sg13g2_decap_8 FILLER_59_637 ();
 sg13g2_decap_8 FILLER_59_644 ();
 sg13g2_decap_8 FILLER_59_651 ();
 sg13g2_decap_8 FILLER_59_658 ();
 sg13g2_decap_8 FILLER_59_665 ();
 sg13g2_decap_8 FILLER_59_672 ();
 sg13g2_decap_8 FILLER_59_679 ();
 sg13g2_decap_8 FILLER_59_686 ();
 sg13g2_decap_8 FILLER_59_693 ();
 sg13g2_decap_8 FILLER_59_700 ();
 sg13g2_decap_8 FILLER_59_707 ();
 sg13g2_decap_8 FILLER_59_714 ();
 sg13g2_decap_8 FILLER_59_721 ();
 sg13g2_decap_8 FILLER_59_728 ();
 sg13g2_decap_8 FILLER_59_735 ();
 sg13g2_decap_8 FILLER_59_742 ();
 sg13g2_decap_8 FILLER_59_749 ();
 sg13g2_decap_8 FILLER_59_756 ();
 sg13g2_decap_8 FILLER_59_763 ();
 sg13g2_decap_8 FILLER_59_770 ();
 sg13g2_decap_8 FILLER_59_777 ();
 sg13g2_decap_8 FILLER_59_784 ();
 sg13g2_decap_8 FILLER_59_791 ();
 sg13g2_decap_8 FILLER_59_798 ();
 sg13g2_decap_8 FILLER_59_805 ();
 sg13g2_decap_8 FILLER_59_812 ();
 sg13g2_decap_8 FILLER_59_819 ();
 sg13g2_decap_8 FILLER_59_826 ();
 sg13g2_decap_8 FILLER_59_833 ();
 sg13g2_fill_1 FILLER_59_840 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_196 ();
 sg13g2_decap_8 FILLER_60_203 ();
 sg13g2_decap_8 FILLER_60_210 ();
 sg13g2_decap_8 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_decap_8 FILLER_60_231 ();
 sg13g2_decap_8 FILLER_60_238 ();
 sg13g2_decap_8 FILLER_60_245 ();
 sg13g2_decap_8 FILLER_60_252 ();
 sg13g2_decap_8 FILLER_60_259 ();
 sg13g2_decap_8 FILLER_60_266 ();
 sg13g2_decap_8 FILLER_60_273 ();
 sg13g2_decap_8 FILLER_60_280 ();
 sg13g2_decap_8 FILLER_60_287 ();
 sg13g2_decap_8 FILLER_60_294 ();
 sg13g2_decap_8 FILLER_60_301 ();
 sg13g2_decap_8 FILLER_60_308 ();
 sg13g2_decap_8 FILLER_60_315 ();
 sg13g2_decap_8 FILLER_60_322 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_decap_8 FILLER_60_336 ();
 sg13g2_decap_8 FILLER_60_343 ();
 sg13g2_decap_8 FILLER_60_350 ();
 sg13g2_decap_8 FILLER_60_357 ();
 sg13g2_decap_8 FILLER_60_364 ();
 sg13g2_decap_8 FILLER_60_371 ();
 sg13g2_decap_8 FILLER_60_378 ();
 sg13g2_decap_8 FILLER_60_385 ();
 sg13g2_decap_8 FILLER_60_392 ();
 sg13g2_decap_8 FILLER_60_399 ();
 sg13g2_decap_8 FILLER_60_406 ();
 sg13g2_decap_8 FILLER_60_413 ();
 sg13g2_decap_8 FILLER_60_420 ();
 sg13g2_decap_8 FILLER_60_427 ();
 sg13g2_decap_8 FILLER_60_434 ();
 sg13g2_decap_8 FILLER_60_441 ();
 sg13g2_decap_8 FILLER_60_448 ();
 sg13g2_decap_8 FILLER_60_455 ();
 sg13g2_decap_8 FILLER_60_462 ();
 sg13g2_decap_8 FILLER_60_469 ();
 sg13g2_decap_8 FILLER_60_476 ();
 sg13g2_decap_8 FILLER_60_483 ();
 sg13g2_decap_8 FILLER_60_490 ();
 sg13g2_decap_8 FILLER_60_497 ();
 sg13g2_decap_8 FILLER_60_504 ();
 sg13g2_decap_8 FILLER_60_511 ();
 sg13g2_decap_8 FILLER_60_518 ();
 sg13g2_decap_8 FILLER_60_525 ();
 sg13g2_decap_8 FILLER_60_532 ();
 sg13g2_decap_8 FILLER_60_539 ();
 sg13g2_decap_8 FILLER_60_546 ();
 sg13g2_decap_8 FILLER_60_553 ();
 sg13g2_decap_8 FILLER_60_560 ();
 sg13g2_decap_8 FILLER_60_567 ();
 sg13g2_decap_8 FILLER_60_574 ();
 sg13g2_decap_8 FILLER_60_581 ();
 sg13g2_decap_8 FILLER_60_588 ();
 sg13g2_decap_8 FILLER_60_595 ();
 sg13g2_decap_8 FILLER_60_602 ();
 sg13g2_decap_8 FILLER_60_609 ();
 sg13g2_decap_8 FILLER_60_616 ();
 sg13g2_decap_8 FILLER_60_623 ();
 sg13g2_decap_8 FILLER_60_630 ();
 sg13g2_decap_8 FILLER_60_637 ();
 sg13g2_decap_8 FILLER_60_644 ();
 sg13g2_decap_8 FILLER_60_651 ();
 sg13g2_decap_8 FILLER_60_658 ();
 sg13g2_decap_8 FILLER_60_665 ();
 sg13g2_decap_8 FILLER_60_672 ();
 sg13g2_decap_8 FILLER_60_679 ();
 sg13g2_decap_8 FILLER_60_686 ();
 sg13g2_decap_8 FILLER_60_693 ();
 sg13g2_decap_8 FILLER_60_700 ();
 sg13g2_decap_8 FILLER_60_707 ();
 sg13g2_decap_8 FILLER_60_714 ();
 sg13g2_decap_8 FILLER_60_721 ();
 sg13g2_decap_8 FILLER_60_728 ();
 sg13g2_decap_8 FILLER_60_735 ();
 sg13g2_decap_8 FILLER_60_742 ();
 sg13g2_decap_8 FILLER_60_749 ();
 sg13g2_decap_8 FILLER_60_756 ();
 sg13g2_decap_8 FILLER_60_763 ();
 sg13g2_decap_8 FILLER_60_770 ();
 sg13g2_decap_8 FILLER_60_777 ();
 sg13g2_decap_8 FILLER_60_784 ();
 sg13g2_decap_8 FILLER_60_791 ();
 sg13g2_decap_8 FILLER_60_798 ();
 sg13g2_decap_8 FILLER_60_805 ();
 sg13g2_decap_8 FILLER_60_812 ();
 sg13g2_decap_8 FILLER_60_819 ();
 sg13g2_decap_8 FILLER_60_826 ();
 sg13g2_decap_8 FILLER_60_833 ();
 sg13g2_fill_1 FILLER_60_840 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_decap_8 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_182 ();
 sg13g2_decap_8 FILLER_61_189 ();
 sg13g2_decap_8 FILLER_61_196 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_decap_8 FILLER_61_217 ();
 sg13g2_decap_8 FILLER_61_224 ();
 sg13g2_decap_8 FILLER_61_231 ();
 sg13g2_decap_8 FILLER_61_238 ();
 sg13g2_decap_8 FILLER_61_245 ();
 sg13g2_decap_8 FILLER_61_252 ();
 sg13g2_decap_8 FILLER_61_259 ();
 sg13g2_decap_8 FILLER_61_266 ();
 sg13g2_decap_8 FILLER_61_273 ();
 sg13g2_decap_8 FILLER_61_280 ();
 sg13g2_decap_8 FILLER_61_287 ();
 sg13g2_decap_8 FILLER_61_294 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_308 ();
 sg13g2_decap_8 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_322 ();
 sg13g2_decap_8 FILLER_61_329 ();
 sg13g2_decap_8 FILLER_61_336 ();
 sg13g2_decap_8 FILLER_61_343 ();
 sg13g2_decap_8 FILLER_61_350 ();
 sg13g2_decap_8 FILLER_61_357 ();
 sg13g2_decap_8 FILLER_61_364 ();
 sg13g2_decap_8 FILLER_61_371 ();
 sg13g2_decap_8 FILLER_61_378 ();
 sg13g2_decap_8 FILLER_61_385 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_decap_8 FILLER_61_406 ();
 sg13g2_decap_8 FILLER_61_413 ();
 sg13g2_decap_8 FILLER_61_420 ();
 sg13g2_decap_8 FILLER_61_427 ();
 sg13g2_decap_8 FILLER_61_434 ();
 sg13g2_decap_8 FILLER_61_441 ();
 sg13g2_decap_8 FILLER_61_448 ();
 sg13g2_decap_8 FILLER_61_455 ();
 sg13g2_decap_8 FILLER_61_462 ();
 sg13g2_decap_8 FILLER_61_469 ();
 sg13g2_decap_8 FILLER_61_476 ();
 sg13g2_decap_8 FILLER_61_483 ();
 sg13g2_decap_8 FILLER_61_490 ();
 sg13g2_decap_8 FILLER_61_497 ();
 sg13g2_decap_8 FILLER_61_504 ();
 sg13g2_decap_8 FILLER_61_511 ();
 sg13g2_decap_8 FILLER_61_518 ();
 sg13g2_decap_8 FILLER_61_525 ();
 sg13g2_decap_8 FILLER_61_532 ();
 sg13g2_decap_8 FILLER_61_539 ();
 sg13g2_decap_8 FILLER_61_546 ();
 sg13g2_decap_8 FILLER_61_553 ();
 sg13g2_decap_8 FILLER_61_560 ();
 sg13g2_decap_8 FILLER_61_567 ();
 sg13g2_decap_8 FILLER_61_574 ();
 sg13g2_decap_8 FILLER_61_581 ();
 sg13g2_decap_8 FILLER_61_588 ();
 sg13g2_decap_8 FILLER_61_595 ();
 sg13g2_decap_8 FILLER_61_602 ();
 sg13g2_decap_8 FILLER_61_609 ();
 sg13g2_decap_8 FILLER_61_616 ();
 sg13g2_decap_8 FILLER_61_623 ();
 sg13g2_decap_8 FILLER_61_630 ();
 sg13g2_decap_8 FILLER_61_637 ();
 sg13g2_decap_8 FILLER_61_644 ();
 sg13g2_decap_8 FILLER_61_651 ();
 sg13g2_decap_8 FILLER_61_658 ();
 sg13g2_decap_8 FILLER_61_665 ();
 sg13g2_decap_8 FILLER_61_672 ();
 sg13g2_decap_8 FILLER_61_679 ();
 sg13g2_decap_8 FILLER_61_686 ();
 sg13g2_decap_8 FILLER_61_693 ();
 sg13g2_decap_8 FILLER_61_700 ();
 sg13g2_decap_8 FILLER_61_707 ();
 sg13g2_decap_8 FILLER_61_714 ();
 sg13g2_decap_8 FILLER_61_721 ();
 sg13g2_decap_8 FILLER_61_728 ();
 sg13g2_decap_8 FILLER_61_735 ();
 sg13g2_decap_8 FILLER_61_742 ();
 sg13g2_decap_8 FILLER_61_749 ();
 sg13g2_decap_8 FILLER_61_756 ();
 sg13g2_decap_8 FILLER_61_763 ();
 sg13g2_decap_8 FILLER_61_770 ();
 sg13g2_decap_8 FILLER_61_777 ();
 sg13g2_decap_8 FILLER_61_784 ();
 sg13g2_decap_8 FILLER_61_791 ();
 sg13g2_decap_8 FILLER_61_798 ();
 sg13g2_decap_8 FILLER_61_805 ();
 sg13g2_decap_8 FILLER_61_812 ();
 sg13g2_decap_8 FILLER_61_819 ();
 sg13g2_decap_8 FILLER_61_826 ();
 sg13g2_decap_8 FILLER_61_833 ();
 sg13g2_fill_1 FILLER_61_840 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_189 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_decap_8 FILLER_62_217 ();
 sg13g2_decap_8 FILLER_62_224 ();
 sg13g2_decap_8 FILLER_62_231 ();
 sg13g2_decap_8 FILLER_62_238 ();
 sg13g2_decap_8 FILLER_62_245 ();
 sg13g2_decap_8 FILLER_62_252 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_decap_8 FILLER_62_266 ();
 sg13g2_decap_8 FILLER_62_273 ();
 sg13g2_decap_8 FILLER_62_280 ();
 sg13g2_decap_8 FILLER_62_287 ();
 sg13g2_decap_8 FILLER_62_294 ();
 sg13g2_decap_8 FILLER_62_301 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_decap_8 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_329 ();
 sg13g2_decap_8 FILLER_62_336 ();
 sg13g2_decap_8 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_8 FILLER_62_385 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_decap_8 FILLER_62_406 ();
 sg13g2_decap_8 FILLER_62_413 ();
 sg13g2_decap_8 FILLER_62_420 ();
 sg13g2_decap_8 FILLER_62_427 ();
 sg13g2_decap_8 FILLER_62_434 ();
 sg13g2_decap_8 FILLER_62_441 ();
 sg13g2_decap_8 FILLER_62_448 ();
 sg13g2_decap_8 FILLER_62_455 ();
 sg13g2_decap_8 FILLER_62_462 ();
 sg13g2_decap_8 FILLER_62_469 ();
 sg13g2_decap_8 FILLER_62_476 ();
 sg13g2_decap_8 FILLER_62_483 ();
 sg13g2_decap_8 FILLER_62_490 ();
 sg13g2_decap_8 FILLER_62_497 ();
 sg13g2_decap_8 FILLER_62_504 ();
 sg13g2_decap_8 FILLER_62_511 ();
 sg13g2_decap_8 FILLER_62_518 ();
 sg13g2_decap_8 FILLER_62_525 ();
 sg13g2_decap_8 FILLER_62_532 ();
 sg13g2_decap_8 FILLER_62_539 ();
 sg13g2_decap_8 FILLER_62_546 ();
 sg13g2_decap_8 FILLER_62_553 ();
 sg13g2_decap_8 FILLER_62_560 ();
 sg13g2_decap_8 FILLER_62_567 ();
 sg13g2_decap_8 FILLER_62_574 ();
 sg13g2_decap_8 FILLER_62_581 ();
 sg13g2_decap_8 FILLER_62_588 ();
 sg13g2_decap_8 FILLER_62_595 ();
 sg13g2_decap_8 FILLER_62_602 ();
 sg13g2_decap_8 FILLER_62_609 ();
 sg13g2_decap_8 FILLER_62_616 ();
 sg13g2_decap_8 FILLER_62_623 ();
 sg13g2_decap_8 FILLER_62_630 ();
 sg13g2_decap_8 FILLER_62_637 ();
 sg13g2_decap_8 FILLER_62_644 ();
 sg13g2_decap_8 FILLER_62_651 ();
 sg13g2_decap_8 FILLER_62_658 ();
 sg13g2_decap_8 FILLER_62_665 ();
 sg13g2_decap_8 FILLER_62_672 ();
 sg13g2_decap_8 FILLER_62_679 ();
 sg13g2_decap_8 FILLER_62_686 ();
 sg13g2_decap_8 FILLER_62_693 ();
 sg13g2_decap_8 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_707 ();
 sg13g2_decap_8 FILLER_62_714 ();
 sg13g2_decap_8 FILLER_62_721 ();
 sg13g2_decap_8 FILLER_62_728 ();
 sg13g2_decap_8 FILLER_62_735 ();
 sg13g2_decap_8 FILLER_62_742 ();
 sg13g2_decap_8 FILLER_62_749 ();
 sg13g2_decap_8 FILLER_62_756 ();
 sg13g2_decap_8 FILLER_62_763 ();
 sg13g2_decap_8 FILLER_62_770 ();
 sg13g2_decap_8 FILLER_62_777 ();
 sg13g2_decap_8 FILLER_62_784 ();
 sg13g2_decap_8 FILLER_62_791 ();
 sg13g2_decap_8 FILLER_62_798 ();
 sg13g2_decap_8 FILLER_62_805 ();
 sg13g2_decap_8 FILLER_62_812 ();
 sg13g2_decap_8 FILLER_62_819 ();
 sg13g2_decap_8 FILLER_62_826 ();
 sg13g2_decap_8 FILLER_62_833 ();
 sg13g2_fill_1 FILLER_62_840 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_8 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_217 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_decap_8 FILLER_63_231 ();
 sg13g2_decap_8 FILLER_63_238 ();
 sg13g2_decap_8 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_252 ();
 sg13g2_decap_8 FILLER_63_259 ();
 sg13g2_decap_8 FILLER_63_266 ();
 sg13g2_decap_8 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_280 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_decap_8 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_301 ();
 sg13g2_decap_8 FILLER_63_308 ();
 sg13g2_decap_8 FILLER_63_315 ();
 sg13g2_decap_8 FILLER_63_322 ();
 sg13g2_decap_8 FILLER_63_329 ();
 sg13g2_decap_8 FILLER_63_336 ();
 sg13g2_decap_8 FILLER_63_343 ();
 sg13g2_decap_8 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_decap_8 FILLER_63_364 ();
 sg13g2_decap_8 FILLER_63_371 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_8 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_decap_8 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_63_406 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_decap_8 FILLER_63_427 ();
 sg13g2_decap_8 FILLER_63_434 ();
 sg13g2_decap_8 FILLER_63_441 ();
 sg13g2_decap_8 FILLER_63_448 ();
 sg13g2_decap_8 FILLER_63_455 ();
 sg13g2_decap_8 FILLER_63_462 ();
 sg13g2_decap_8 FILLER_63_469 ();
 sg13g2_decap_8 FILLER_63_476 ();
 sg13g2_decap_8 FILLER_63_483 ();
 sg13g2_decap_8 FILLER_63_490 ();
 sg13g2_decap_8 FILLER_63_497 ();
 sg13g2_decap_8 FILLER_63_504 ();
 sg13g2_decap_8 FILLER_63_511 ();
 sg13g2_decap_8 FILLER_63_518 ();
 sg13g2_decap_8 FILLER_63_525 ();
 sg13g2_decap_8 FILLER_63_532 ();
 sg13g2_decap_8 FILLER_63_539 ();
 sg13g2_decap_8 FILLER_63_546 ();
 sg13g2_decap_8 FILLER_63_553 ();
 sg13g2_decap_8 FILLER_63_560 ();
 sg13g2_decap_8 FILLER_63_567 ();
 sg13g2_decap_8 FILLER_63_574 ();
 sg13g2_decap_8 FILLER_63_581 ();
 sg13g2_decap_8 FILLER_63_588 ();
 sg13g2_decap_8 FILLER_63_595 ();
 sg13g2_decap_8 FILLER_63_602 ();
 sg13g2_decap_8 FILLER_63_609 ();
 sg13g2_decap_8 FILLER_63_616 ();
 sg13g2_decap_8 FILLER_63_623 ();
 sg13g2_decap_8 FILLER_63_630 ();
 sg13g2_decap_8 FILLER_63_637 ();
 sg13g2_decap_8 FILLER_63_644 ();
 sg13g2_decap_8 FILLER_63_651 ();
 sg13g2_decap_8 FILLER_63_658 ();
 sg13g2_decap_8 FILLER_63_665 ();
 sg13g2_decap_8 FILLER_63_672 ();
 sg13g2_decap_8 FILLER_63_679 ();
 sg13g2_decap_8 FILLER_63_686 ();
 sg13g2_decap_8 FILLER_63_693 ();
 sg13g2_decap_8 FILLER_63_700 ();
 sg13g2_decap_8 FILLER_63_707 ();
 sg13g2_decap_8 FILLER_63_714 ();
 sg13g2_decap_8 FILLER_63_721 ();
 sg13g2_decap_8 FILLER_63_728 ();
 sg13g2_decap_8 FILLER_63_735 ();
 sg13g2_decap_8 FILLER_63_742 ();
 sg13g2_decap_8 FILLER_63_749 ();
 sg13g2_decap_8 FILLER_63_756 ();
 sg13g2_decap_8 FILLER_63_763 ();
 sg13g2_decap_8 FILLER_63_770 ();
 sg13g2_decap_8 FILLER_63_777 ();
 sg13g2_decap_8 FILLER_63_784 ();
 sg13g2_decap_8 FILLER_63_791 ();
 sg13g2_decap_8 FILLER_63_798 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_decap_8 FILLER_63_812 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_833 ();
 sg13g2_fill_1 FILLER_63_840 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_168 ();
 sg13g2_decap_8 FILLER_64_175 ();
 sg13g2_decap_8 FILLER_64_182 ();
 sg13g2_decap_8 FILLER_64_189 ();
 sg13g2_decap_8 FILLER_64_196 ();
 sg13g2_decap_8 FILLER_64_203 ();
 sg13g2_decap_8 FILLER_64_210 ();
 sg13g2_decap_8 FILLER_64_217 ();
 sg13g2_decap_8 FILLER_64_224 ();
 sg13g2_decap_8 FILLER_64_231 ();
 sg13g2_decap_8 FILLER_64_238 ();
 sg13g2_decap_8 FILLER_64_245 ();
 sg13g2_decap_8 FILLER_64_252 ();
 sg13g2_decap_8 FILLER_64_259 ();
 sg13g2_decap_8 FILLER_64_266 ();
 sg13g2_decap_8 FILLER_64_273 ();
 sg13g2_decap_8 FILLER_64_280 ();
 sg13g2_decap_8 FILLER_64_287 ();
 sg13g2_decap_8 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_301 ();
 sg13g2_decap_8 FILLER_64_308 ();
 sg13g2_decap_8 FILLER_64_315 ();
 sg13g2_decap_8 FILLER_64_322 ();
 sg13g2_decap_8 FILLER_64_329 ();
 sg13g2_decap_8 FILLER_64_336 ();
 sg13g2_decap_8 FILLER_64_343 ();
 sg13g2_decap_8 FILLER_64_350 ();
 sg13g2_decap_8 FILLER_64_357 ();
 sg13g2_decap_8 FILLER_64_364 ();
 sg13g2_decap_8 FILLER_64_371 ();
 sg13g2_decap_8 FILLER_64_378 ();
 sg13g2_decap_8 FILLER_64_385 ();
 sg13g2_decap_8 FILLER_64_392 ();
 sg13g2_decap_8 FILLER_64_399 ();
 sg13g2_decap_8 FILLER_64_406 ();
 sg13g2_decap_8 FILLER_64_413 ();
 sg13g2_decap_8 FILLER_64_420 ();
 sg13g2_decap_8 FILLER_64_427 ();
 sg13g2_decap_8 FILLER_64_434 ();
 sg13g2_decap_8 FILLER_64_441 ();
 sg13g2_decap_8 FILLER_64_448 ();
 sg13g2_decap_8 FILLER_64_455 ();
 sg13g2_decap_8 FILLER_64_462 ();
 sg13g2_decap_8 FILLER_64_469 ();
 sg13g2_decap_8 FILLER_64_476 ();
 sg13g2_decap_8 FILLER_64_483 ();
 sg13g2_decap_8 FILLER_64_490 ();
 sg13g2_decap_8 FILLER_64_497 ();
 sg13g2_decap_8 FILLER_64_504 ();
 sg13g2_decap_8 FILLER_64_511 ();
 sg13g2_decap_8 FILLER_64_518 ();
 sg13g2_decap_8 FILLER_64_525 ();
 sg13g2_decap_8 FILLER_64_532 ();
 sg13g2_decap_8 FILLER_64_539 ();
 sg13g2_decap_8 FILLER_64_546 ();
 sg13g2_decap_8 FILLER_64_553 ();
 sg13g2_decap_8 FILLER_64_560 ();
 sg13g2_decap_8 FILLER_64_567 ();
 sg13g2_decap_8 FILLER_64_574 ();
 sg13g2_decap_8 FILLER_64_581 ();
 sg13g2_decap_8 FILLER_64_588 ();
 sg13g2_decap_8 FILLER_64_595 ();
 sg13g2_decap_8 FILLER_64_602 ();
 sg13g2_decap_8 FILLER_64_609 ();
 sg13g2_decap_8 FILLER_64_616 ();
 sg13g2_decap_8 FILLER_64_623 ();
 sg13g2_decap_8 FILLER_64_630 ();
 sg13g2_decap_8 FILLER_64_637 ();
 sg13g2_decap_8 FILLER_64_644 ();
 sg13g2_decap_8 FILLER_64_651 ();
 sg13g2_decap_8 FILLER_64_658 ();
 sg13g2_decap_8 FILLER_64_665 ();
 sg13g2_decap_8 FILLER_64_672 ();
 sg13g2_decap_8 FILLER_64_679 ();
 sg13g2_decap_8 FILLER_64_686 ();
 sg13g2_decap_8 FILLER_64_693 ();
 sg13g2_decap_8 FILLER_64_700 ();
 sg13g2_decap_8 FILLER_64_707 ();
 sg13g2_decap_8 FILLER_64_714 ();
 sg13g2_decap_8 FILLER_64_721 ();
 sg13g2_decap_8 FILLER_64_728 ();
 sg13g2_decap_8 FILLER_64_735 ();
 sg13g2_decap_8 FILLER_64_742 ();
 sg13g2_decap_8 FILLER_64_749 ();
 sg13g2_decap_8 FILLER_64_756 ();
 sg13g2_decap_8 FILLER_64_763 ();
 sg13g2_decap_8 FILLER_64_770 ();
 sg13g2_decap_8 FILLER_64_777 ();
 sg13g2_decap_8 FILLER_64_784 ();
 sg13g2_decap_8 FILLER_64_791 ();
 sg13g2_decap_8 FILLER_64_798 ();
 sg13g2_decap_8 FILLER_64_805 ();
 sg13g2_decap_8 FILLER_64_812 ();
 sg13g2_decap_8 FILLER_64_819 ();
 sg13g2_decap_8 FILLER_64_826 ();
 sg13g2_decap_8 FILLER_64_833 ();
 sg13g2_fill_1 FILLER_64_840 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_189 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_8 FILLER_65_203 ();
 sg13g2_decap_8 FILLER_65_210 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_238 ();
 sg13g2_decap_8 FILLER_65_245 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_decap_8 FILLER_65_259 ();
 sg13g2_decap_8 FILLER_65_266 ();
 sg13g2_decap_8 FILLER_65_273 ();
 sg13g2_decap_8 FILLER_65_280 ();
 sg13g2_decap_8 FILLER_65_287 ();
 sg13g2_decap_8 FILLER_65_294 ();
 sg13g2_decap_8 FILLER_65_301 ();
 sg13g2_decap_8 FILLER_65_308 ();
 sg13g2_decap_8 FILLER_65_315 ();
 sg13g2_decap_8 FILLER_65_322 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_decap_8 FILLER_65_336 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_350 ();
 sg13g2_decap_8 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_decap_8 FILLER_65_406 ();
 sg13g2_decap_8 FILLER_65_413 ();
 sg13g2_decap_8 FILLER_65_420 ();
 sg13g2_decap_8 FILLER_65_427 ();
 sg13g2_decap_8 FILLER_65_434 ();
 sg13g2_decap_8 FILLER_65_441 ();
 sg13g2_decap_8 FILLER_65_448 ();
 sg13g2_decap_8 FILLER_65_455 ();
 sg13g2_decap_8 FILLER_65_462 ();
 sg13g2_decap_8 FILLER_65_469 ();
 sg13g2_decap_8 FILLER_65_476 ();
 sg13g2_decap_8 FILLER_65_483 ();
 sg13g2_decap_8 FILLER_65_490 ();
 sg13g2_decap_8 FILLER_65_497 ();
 sg13g2_decap_8 FILLER_65_504 ();
 sg13g2_decap_8 FILLER_65_511 ();
 sg13g2_decap_8 FILLER_65_518 ();
 sg13g2_decap_8 FILLER_65_525 ();
 sg13g2_decap_8 FILLER_65_532 ();
 sg13g2_decap_8 FILLER_65_539 ();
 sg13g2_decap_8 FILLER_65_546 ();
 sg13g2_decap_8 FILLER_65_553 ();
 sg13g2_decap_8 FILLER_65_560 ();
 sg13g2_decap_8 FILLER_65_567 ();
 sg13g2_decap_8 FILLER_65_574 ();
 sg13g2_decap_8 FILLER_65_581 ();
 sg13g2_decap_8 FILLER_65_588 ();
 sg13g2_decap_8 FILLER_65_595 ();
 sg13g2_decap_8 FILLER_65_602 ();
 sg13g2_decap_8 FILLER_65_609 ();
 sg13g2_decap_8 FILLER_65_616 ();
 sg13g2_decap_8 FILLER_65_623 ();
 sg13g2_decap_8 FILLER_65_630 ();
 sg13g2_decap_8 FILLER_65_637 ();
 sg13g2_decap_8 FILLER_65_644 ();
 sg13g2_decap_8 FILLER_65_651 ();
 sg13g2_decap_8 FILLER_65_658 ();
 sg13g2_decap_8 FILLER_65_665 ();
 sg13g2_decap_8 FILLER_65_672 ();
 sg13g2_decap_8 FILLER_65_679 ();
 sg13g2_decap_8 FILLER_65_686 ();
 sg13g2_decap_8 FILLER_65_693 ();
 sg13g2_decap_8 FILLER_65_700 ();
 sg13g2_decap_8 FILLER_65_707 ();
 sg13g2_decap_8 FILLER_65_714 ();
 sg13g2_decap_8 FILLER_65_721 ();
 sg13g2_decap_8 FILLER_65_728 ();
 sg13g2_decap_8 FILLER_65_735 ();
 sg13g2_decap_8 FILLER_65_742 ();
 sg13g2_decap_8 FILLER_65_749 ();
 sg13g2_decap_8 FILLER_65_756 ();
 sg13g2_decap_8 FILLER_65_763 ();
 sg13g2_decap_8 FILLER_65_770 ();
 sg13g2_decap_8 FILLER_65_777 ();
 sg13g2_decap_8 FILLER_65_784 ();
 sg13g2_decap_8 FILLER_65_791 ();
 sg13g2_decap_8 FILLER_65_798 ();
 sg13g2_decap_8 FILLER_65_805 ();
 sg13g2_decap_8 FILLER_65_812 ();
 sg13g2_decap_8 FILLER_65_819 ();
 sg13g2_decap_8 FILLER_65_826 ();
 sg13g2_decap_8 FILLER_65_833 ();
 sg13g2_fill_1 FILLER_65_840 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_8 FILLER_66_182 ();
 sg13g2_decap_8 FILLER_66_189 ();
 sg13g2_decap_8 FILLER_66_196 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_217 ();
 sg13g2_decap_8 FILLER_66_224 ();
 sg13g2_decap_8 FILLER_66_231 ();
 sg13g2_decap_8 FILLER_66_238 ();
 sg13g2_decap_8 FILLER_66_245 ();
 sg13g2_decap_8 FILLER_66_252 ();
 sg13g2_decap_8 FILLER_66_259 ();
 sg13g2_decap_8 FILLER_66_266 ();
 sg13g2_decap_8 FILLER_66_273 ();
 sg13g2_decap_8 FILLER_66_280 ();
 sg13g2_decap_8 FILLER_66_287 ();
 sg13g2_decap_8 FILLER_66_294 ();
 sg13g2_decap_8 FILLER_66_301 ();
 sg13g2_decap_8 FILLER_66_308 ();
 sg13g2_decap_8 FILLER_66_315 ();
 sg13g2_decap_8 FILLER_66_322 ();
 sg13g2_decap_8 FILLER_66_329 ();
 sg13g2_decap_8 FILLER_66_336 ();
 sg13g2_decap_8 FILLER_66_343 ();
 sg13g2_decap_8 FILLER_66_350 ();
 sg13g2_decap_8 FILLER_66_357 ();
 sg13g2_decap_8 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_371 ();
 sg13g2_decap_8 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_385 ();
 sg13g2_decap_8 FILLER_66_392 ();
 sg13g2_decap_8 FILLER_66_399 ();
 sg13g2_decap_8 FILLER_66_406 ();
 sg13g2_decap_8 FILLER_66_413 ();
 sg13g2_decap_8 FILLER_66_420 ();
 sg13g2_decap_8 FILLER_66_427 ();
 sg13g2_decap_8 FILLER_66_434 ();
 sg13g2_decap_8 FILLER_66_441 ();
 sg13g2_decap_8 FILLER_66_448 ();
 sg13g2_decap_8 FILLER_66_455 ();
 sg13g2_decap_8 FILLER_66_462 ();
 sg13g2_decap_8 FILLER_66_469 ();
 sg13g2_decap_8 FILLER_66_476 ();
 sg13g2_decap_8 FILLER_66_483 ();
 sg13g2_decap_8 FILLER_66_490 ();
 sg13g2_decap_8 FILLER_66_497 ();
 sg13g2_decap_8 FILLER_66_504 ();
 sg13g2_decap_8 FILLER_66_511 ();
 sg13g2_decap_8 FILLER_66_518 ();
 sg13g2_decap_8 FILLER_66_525 ();
 sg13g2_decap_8 FILLER_66_532 ();
 sg13g2_decap_8 FILLER_66_539 ();
 sg13g2_decap_8 FILLER_66_546 ();
 sg13g2_decap_8 FILLER_66_553 ();
 sg13g2_decap_8 FILLER_66_560 ();
 sg13g2_decap_8 FILLER_66_567 ();
 sg13g2_decap_8 FILLER_66_574 ();
 sg13g2_decap_8 FILLER_66_581 ();
 sg13g2_decap_8 FILLER_66_588 ();
 sg13g2_decap_8 FILLER_66_595 ();
 sg13g2_decap_8 FILLER_66_602 ();
 sg13g2_decap_8 FILLER_66_609 ();
 sg13g2_decap_8 FILLER_66_616 ();
 sg13g2_decap_8 FILLER_66_623 ();
 sg13g2_decap_8 FILLER_66_630 ();
 sg13g2_decap_8 FILLER_66_637 ();
 sg13g2_decap_8 FILLER_66_644 ();
 sg13g2_decap_8 FILLER_66_651 ();
 sg13g2_decap_8 FILLER_66_658 ();
 sg13g2_decap_8 FILLER_66_665 ();
 sg13g2_decap_8 FILLER_66_672 ();
 sg13g2_decap_8 FILLER_66_679 ();
 sg13g2_decap_8 FILLER_66_686 ();
 sg13g2_decap_8 FILLER_66_693 ();
 sg13g2_decap_8 FILLER_66_700 ();
 sg13g2_decap_8 FILLER_66_707 ();
 sg13g2_decap_8 FILLER_66_714 ();
 sg13g2_decap_8 FILLER_66_721 ();
 sg13g2_decap_8 FILLER_66_728 ();
 sg13g2_decap_8 FILLER_66_735 ();
 sg13g2_decap_8 FILLER_66_742 ();
 sg13g2_decap_8 FILLER_66_749 ();
 sg13g2_decap_8 FILLER_66_756 ();
 sg13g2_decap_8 FILLER_66_763 ();
 sg13g2_decap_8 FILLER_66_770 ();
 sg13g2_decap_8 FILLER_66_777 ();
 sg13g2_decap_8 FILLER_66_784 ();
 sg13g2_decap_8 FILLER_66_791 ();
 sg13g2_decap_8 FILLER_66_798 ();
 sg13g2_decap_8 FILLER_66_805 ();
 sg13g2_decap_8 FILLER_66_812 ();
 sg13g2_decap_8 FILLER_66_819 ();
 sg13g2_decap_8 FILLER_66_826 ();
 sg13g2_decap_8 FILLER_66_833 ();
 sg13g2_fill_1 FILLER_66_840 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_decap_8 FILLER_67_252 ();
 sg13g2_decap_8 FILLER_67_259 ();
 sg13g2_decap_8 FILLER_67_266 ();
 sg13g2_decap_8 FILLER_67_273 ();
 sg13g2_decap_8 FILLER_67_280 ();
 sg13g2_decap_8 FILLER_67_287 ();
 sg13g2_decap_8 FILLER_67_294 ();
 sg13g2_decap_8 FILLER_67_301 ();
 sg13g2_decap_8 FILLER_67_308 ();
 sg13g2_decap_8 FILLER_67_315 ();
 sg13g2_decap_8 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_329 ();
 sg13g2_decap_8 FILLER_67_336 ();
 sg13g2_decap_8 FILLER_67_343 ();
 sg13g2_decap_8 FILLER_67_350 ();
 sg13g2_decap_8 FILLER_67_357 ();
 sg13g2_decap_8 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_67_378 ();
 sg13g2_decap_8 FILLER_67_385 ();
 sg13g2_decap_8 FILLER_67_392 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_decap_8 FILLER_67_406 ();
 sg13g2_decap_8 FILLER_67_413 ();
 sg13g2_decap_8 FILLER_67_420 ();
 sg13g2_decap_8 FILLER_67_427 ();
 sg13g2_decap_8 FILLER_67_434 ();
 sg13g2_decap_8 FILLER_67_441 ();
 sg13g2_decap_8 FILLER_67_448 ();
 sg13g2_decap_8 FILLER_67_455 ();
 sg13g2_decap_8 FILLER_67_462 ();
 sg13g2_decap_8 FILLER_67_469 ();
 sg13g2_decap_8 FILLER_67_476 ();
 sg13g2_decap_8 FILLER_67_483 ();
 sg13g2_decap_8 FILLER_67_490 ();
 sg13g2_decap_8 FILLER_67_497 ();
 sg13g2_decap_8 FILLER_67_504 ();
 sg13g2_decap_8 FILLER_67_511 ();
 sg13g2_decap_8 FILLER_67_518 ();
 sg13g2_decap_8 FILLER_67_525 ();
 sg13g2_decap_8 FILLER_67_532 ();
 sg13g2_decap_8 FILLER_67_539 ();
 sg13g2_decap_8 FILLER_67_546 ();
 sg13g2_decap_8 FILLER_67_553 ();
 sg13g2_decap_8 FILLER_67_560 ();
 sg13g2_decap_8 FILLER_67_567 ();
 sg13g2_decap_8 FILLER_67_574 ();
 sg13g2_decap_8 FILLER_67_581 ();
 sg13g2_decap_8 FILLER_67_588 ();
 sg13g2_decap_8 FILLER_67_595 ();
 sg13g2_decap_8 FILLER_67_602 ();
 sg13g2_decap_8 FILLER_67_609 ();
 sg13g2_decap_8 FILLER_67_616 ();
 sg13g2_decap_8 FILLER_67_623 ();
 sg13g2_decap_8 FILLER_67_630 ();
 sg13g2_decap_8 FILLER_67_637 ();
 sg13g2_decap_8 FILLER_67_644 ();
 sg13g2_decap_8 FILLER_67_651 ();
 sg13g2_decap_8 FILLER_67_658 ();
 sg13g2_decap_8 FILLER_67_665 ();
 sg13g2_decap_8 FILLER_67_672 ();
 sg13g2_decap_8 FILLER_67_679 ();
 sg13g2_decap_8 FILLER_67_686 ();
 sg13g2_decap_8 FILLER_67_693 ();
 sg13g2_decap_8 FILLER_67_700 ();
 sg13g2_decap_8 FILLER_67_707 ();
 sg13g2_decap_8 FILLER_67_714 ();
 sg13g2_decap_8 FILLER_67_721 ();
 sg13g2_decap_8 FILLER_67_728 ();
 sg13g2_decap_8 FILLER_67_735 ();
 sg13g2_decap_8 FILLER_67_742 ();
 sg13g2_decap_8 FILLER_67_749 ();
 sg13g2_decap_8 FILLER_67_756 ();
 sg13g2_decap_8 FILLER_67_763 ();
 sg13g2_decap_8 FILLER_67_770 ();
 sg13g2_decap_8 FILLER_67_777 ();
 sg13g2_decap_8 FILLER_67_784 ();
 sg13g2_decap_8 FILLER_67_791 ();
 sg13g2_decap_8 FILLER_67_798 ();
 sg13g2_decap_8 FILLER_67_805 ();
 sg13g2_decap_8 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_819 ();
 sg13g2_decap_8 FILLER_67_826 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_fill_1 FILLER_67_840 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_decap_8 FILLER_68_189 ();
 sg13g2_decap_8 FILLER_68_196 ();
 sg13g2_decap_8 FILLER_68_203 ();
 sg13g2_decap_8 FILLER_68_210 ();
 sg13g2_decap_8 FILLER_68_217 ();
 sg13g2_decap_8 FILLER_68_224 ();
 sg13g2_decap_8 FILLER_68_231 ();
 sg13g2_decap_8 FILLER_68_238 ();
 sg13g2_decap_8 FILLER_68_245 ();
 sg13g2_decap_8 FILLER_68_252 ();
 sg13g2_decap_8 FILLER_68_259 ();
 sg13g2_decap_8 FILLER_68_266 ();
 sg13g2_decap_8 FILLER_68_273 ();
 sg13g2_decap_8 FILLER_68_280 ();
 sg13g2_decap_8 FILLER_68_287 ();
 sg13g2_decap_8 FILLER_68_294 ();
 sg13g2_decap_8 FILLER_68_301 ();
 sg13g2_decap_8 FILLER_68_308 ();
 sg13g2_decap_8 FILLER_68_315 ();
 sg13g2_decap_8 FILLER_68_322 ();
 sg13g2_decap_8 FILLER_68_329 ();
 sg13g2_decap_8 FILLER_68_336 ();
 sg13g2_decap_8 FILLER_68_343 ();
 sg13g2_decap_8 FILLER_68_350 ();
 sg13g2_decap_8 FILLER_68_357 ();
 sg13g2_decap_8 FILLER_68_364 ();
 sg13g2_decap_8 FILLER_68_371 ();
 sg13g2_decap_8 FILLER_68_378 ();
 sg13g2_decap_8 FILLER_68_385 ();
 sg13g2_decap_8 FILLER_68_392 ();
 sg13g2_decap_8 FILLER_68_399 ();
 sg13g2_decap_8 FILLER_68_406 ();
 sg13g2_decap_8 FILLER_68_413 ();
 sg13g2_decap_8 FILLER_68_420 ();
 sg13g2_decap_8 FILLER_68_427 ();
 sg13g2_decap_8 FILLER_68_434 ();
 sg13g2_decap_8 FILLER_68_441 ();
 sg13g2_decap_8 FILLER_68_448 ();
 sg13g2_decap_8 FILLER_68_455 ();
 sg13g2_decap_8 FILLER_68_462 ();
 sg13g2_decap_8 FILLER_68_469 ();
 sg13g2_decap_8 FILLER_68_476 ();
 sg13g2_decap_8 FILLER_68_483 ();
 sg13g2_decap_8 FILLER_68_490 ();
 sg13g2_decap_8 FILLER_68_497 ();
 sg13g2_decap_8 FILLER_68_504 ();
 sg13g2_decap_8 FILLER_68_511 ();
 sg13g2_decap_8 FILLER_68_518 ();
 sg13g2_decap_8 FILLER_68_525 ();
 sg13g2_decap_8 FILLER_68_532 ();
 sg13g2_decap_8 FILLER_68_539 ();
 sg13g2_decap_8 FILLER_68_546 ();
 sg13g2_decap_8 FILLER_68_553 ();
 sg13g2_decap_8 FILLER_68_560 ();
 sg13g2_decap_8 FILLER_68_567 ();
 sg13g2_decap_8 FILLER_68_574 ();
 sg13g2_decap_8 FILLER_68_581 ();
 sg13g2_decap_8 FILLER_68_588 ();
 sg13g2_decap_8 FILLER_68_595 ();
 sg13g2_decap_8 FILLER_68_602 ();
 sg13g2_decap_8 FILLER_68_609 ();
 sg13g2_decap_8 FILLER_68_616 ();
 sg13g2_decap_8 FILLER_68_623 ();
 sg13g2_decap_8 FILLER_68_630 ();
 sg13g2_decap_8 FILLER_68_637 ();
 sg13g2_decap_8 FILLER_68_644 ();
 sg13g2_decap_8 FILLER_68_651 ();
 sg13g2_decap_8 FILLER_68_658 ();
 sg13g2_decap_8 FILLER_68_665 ();
 sg13g2_decap_8 FILLER_68_672 ();
 sg13g2_decap_8 FILLER_68_679 ();
 sg13g2_decap_8 FILLER_68_686 ();
 sg13g2_decap_8 FILLER_68_693 ();
 sg13g2_decap_8 FILLER_68_700 ();
 sg13g2_decap_8 FILLER_68_707 ();
 sg13g2_decap_8 FILLER_68_714 ();
 sg13g2_decap_8 FILLER_68_721 ();
 sg13g2_decap_8 FILLER_68_728 ();
 sg13g2_decap_8 FILLER_68_735 ();
 sg13g2_decap_8 FILLER_68_742 ();
 sg13g2_decap_8 FILLER_68_749 ();
 sg13g2_decap_8 FILLER_68_756 ();
 sg13g2_decap_8 FILLER_68_763 ();
 sg13g2_decap_8 FILLER_68_770 ();
 sg13g2_decap_8 FILLER_68_777 ();
 sg13g2_decap_8 FILLER_68_784 ();
 sg13g2_decap_8 FILLER_68_791 ();
 sg13g2_decap_8 FILLER_68_798 ();
 sg13g2_decap_8 FILLER_68_805 ();
 sg13g2_decap_8 FILLER_68_812 ();
 sg13g2_decap_8 FILLER_68_819 ();
 sg13g2_decap_8 FILLER_68_826 ();
 sg13g2_decap_8 FILLER_68_833 ();
 sg13g2_fill_1 FILLER_68_840 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_decap_8 FILLER_69_168 ();
 sg13g2_decap_8 FILLER_69_175 ();
 sg13g2_decap_8 FILLER_69_182 ();
 sg13g2_decap_8 FILLER_69_189 ();
 sg13g2_decap_8 FILLER_69_196 ();
 sg13g2_decap_8 FILLER_69_203 ();
 sg13g2_decap_8 FILLER_69_210 ();
 sg13g2_decap_8 FILLER_69_217 ();
 sg13g2_decap_8 FILLER_69_224 ();
 sg13g2_decap_8 FILLER_69_231 ();
 sg13g2_decap_8 FILLER_69_238 ();
 sg13g2_decap_8 FILLER_69_245 ();
 sg13g2_decap_8 FILLER_69_252 ();
 sg13g2_decap_8 FILLER_69_259 ();
 sg13g2_decap_8 FILLER_69_266 ();
 sg13g2_decap_8 FILLER_69_273 ();
 sg13g2_decap_8 FILLER_69_280 ();
 sg13g2_decap_8 FILLER_69_287 ();
 sg13g2_decap_8 FILLER_69_294 ();
 sg13g2_decap_8 FILLER_69_301 ();
 sg13g2_decap_8 FILLER_69_308 ();
 sg13g2_decap_8 FILLER_69_315 ();
 sg13g2_decap_8 FILLER_69_322 ();
 sg13g2_decap_8 FILLER_69_329 ();
 sg13g2_decap_8 FILLER_69_336 ();
 sg13g2_decap_8 FILLER_69_343 ();
 sg13g2_decap_8 FILLER_69_350 ();
 sg13g2_decap_8 FILLER_69_357 ();
 sg13g2_decap_8 FILLER_69_364 ();
 sg13g2_decap_8 FILLER_69_371 ();
 sg13g2_decap_8 FILLER_69_378 ();
 sg13g2_decap_8 FILLER_69_385 ();
 sg13g2_decap_8 FILLER_69_392 ();
 sg13g2_decap_8 FILLER_69_399 ();
 sg13g2_decap_8 FILLER_69_406 ();
 sg13g2_decap_8 FILLER_69_413 ();
 sg13g2_decap_8 FILLER_69_420 ();
 sg13g2_decap_8 FILLER_69_427 ();
 sg13g2_decap_8 FILLER_69_434 ();
 sg13g2_decap_8 FILLER_69_441 ();
 sg13g2_decap_8 FILLER_69_448 ();
 sg13g2_decap_8 FILLER_69_455 ();
 sg13g2_decap_8 FILLER_69_462 ();
 sg13g2_decap_8 FILLER_69_469 ();
 sg13g2_decap_8 FILLER_69_476 ();
 sg13g2_decap_8 FILLER_69_483 ();
 sg13g2_decap_8 FILLER_69_490 ();
 sg13g2_decap_8 FILLER_69_497 ();
 sg13g2_decap_8 FILLER_69_504 ();
 sg13g2_decap_8 FILLER_69_511 ();
 sg13g2_decap_8 FILLER_69_518 ();
 sg13g2_decap_8 FILLER_69_525 ();
 sg13g2_decap_8 FILLER_69_532 ();
 sg13g2_decap_8 FILLER_69_539 ();
 sg13g2_decap_8 FILLER_69_546 ();
 sg13g2_decap_8 FILLER_69_553 ();
 sg13g2_decap_8 FILLER_69_560 ();
 sg13g2_decap_8 FILLER_69_567 ();
 sg13g2_decap_8 FILLER_69_574 ();
 sg13g2_decap_8 FILLER_69_581 ();
 sg13g2_decap_8 FILLER_69_588 ();
 sg13g2_decap_8 FILLER_69_595 ();
 sg13g2_decap_8 FILLER_69_602 ();
 sg13g2_decap_8 FILLER_69_609 ();
 sg13g2_decap_8 FILLER_69_616 ();
 sg13g2_decap_8 FILLER_69_623 ();
 sg13g2_decap_8 FILLER_69_630 ();
 sg13g2_decap_8 FILLER_69_637 ();
 sg13g2_decap_8 FILLER_69_644 ();
 sg13g2_decap_8 FILLER_69_651 ();
 sg13g2_decap_8 FILLER_69_658 ();
 sg13g2_decap_8 FILLER_69_665 ();
 sg13g2_decap_8 FILLER_69_672 ();
 sg13g2_decap_8 FILLER_69_679 ();
 sg13g2_decap_8 FILLER_69_686 ();
 sg13g2_decap_8 FILLER_69_693 ();
 sg13g2_decap_8 FILLER_69_700 ();
 sg13g2_decap_8 FILLER_69_707 ();
 sg13g2_decap_8 FILLER_69_714 ();
 sg13g2_decap_8 FILLER_69_721 ();
 sg13g2_decap_8 FILLER_69_728 ();
 sg13g2_decap_8 FILLER_69_735 ();
 sg13g2_decap_8 FILLER_69_742 ();
 sg13g2_decap_8 FILLER_69_749 ();
 sg13g2_decap_8 FILLER_69_756 ();
 sg13g2_decap_8 FILLER_69_763 ();
 sg13g2_decap_8 FILLER_69_770 ();
 sg13g2_decap_8 FILLER_69_777 ();
 sg13g2_decap_8 FILLER_69_784 ();
 sg13g2_decap_8 FILLER_69_791 ();
 sg13g2_decap_8 FILLER_69_798 ();
 sg13g2_decap_8 FILLER_69_805 ();
 sg13g2_decap_8 FILLER_69_812 ();
 sg13g2_decap_8 FILLER_69_819 ();
 sg13g2_decap_8 FILLER_69_826 ();
 sg13g2_decap_8 FILLER_69_833 ();
 sg13g2_fill_1 FILLER_69_840 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_decap_8 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_196 ();
 sg13g2_decap_8 FILLER_70_203 ();
 sg13g2_decap_8 FILLER_70_210 ();
 sg13g2_decap_8 FILLER_70_217 ();
 sg13g2_decap_8 FILLER_70_224 ();
 sg13g2_decap_8 FILLER_70_231 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_decap_8 FILLER_70_245 ();
 sg13g2_decap_8 FILLER_70_252 ();
 sg13g2_decap_8 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_266 ();
 sg13g2_decap_8 FILLER_70_273 ();
 sg13g2_decap_8 FILLER_70_280 ();
 sg13g2_decap_8 FILLER_70_287 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_decap_8 FILLER_70_301 ();
 sg13g2_decap_8 FILLER_70_308 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_322 ();
 sg13g2_decap_8 FILLER_70_329 ();
 sg13g2_decap_8 FILLER_70_336 ();
 sg13g2_decap_8 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_decap_8 FILLER_70_357 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_decap_8 FILLER_70_371 ();
 sg13g2_decap_8 FILLER_70_378 ();
 sg13g2_decap_8 FILLER_70_385 ();
 sg13g2_decap_8 FILLER_70_392 ();
 sg13g2_decap_8 FILLER_70_399 ();
 sg13g2_decap_8 FILLER_70_406 ();
 sg13g2_decap_8 FILLER_70_413 ();
 sg13g2_decap_8 FILLER_70_420 ();
 sg13g2_decap_8 FILLER_70_427 ();
 sg13g2_decap_8 FILLER_70_434 ();
 sg13g2_decap_8 FILLER_70_441 ();
 sg13g2_decap_8 FILLER_70_448 ();
 sg13g2_decap_8 FILLER_70_455 ();
 sg13g2_decap_8 FILLER_70_462 ();
 sg13g2_decap_8 FILLER_70_469 ();
 sg13g2_decap_8 FILLER_70_476 ();
 sg13g2_decap_8 FILLER_70_483 ();
 sg13g2_decap_8 FILLER_70_490 ();
 sg13g2_decap_8 FILLER_70_497 ();
 sg13g2_decap_8 FILLER_70_504 ();
 sg13g2_decap_8 FILLER_70_511 ();
 sg13g2_decap_8 FILLER_70_518 ();
 sg13g2_decap_8 FILLER_70_525 ();
 sg13g2_decap_8 FILLER_70_532 ();
 sg13g2_decap_8 FILLER_70_539 ();
 sg13g2_decap_8 FILLER_70_546 ();
 sg13g2_decap_8 FILLER_70_553 ();
 sg13g2_decap_8 FILLER_70_560 ();
 sg13g2_decap_8 FILLER_70_567 ();
 sg13g2_decap_8 FILLER_70_574 ();
 sg13g2_decap_8 FILLER_70_581 ();
 sg13g2_decap_8 FILLER_70_588 ();
 sg13g2_decap_8 FILLER_70_595 ();
 sg13g2_decap_8 FILLER_70_602 ();
 sg13g2_decap_8 FILLER_70_609 ();
 sg13g2_decap_8 FILLER_70_616 ();
 sg13g2_decap_8 FILLER_70_623 ();
 sg13g2_decap_8 FILLER_70_630 ();
 sg13g2_decap_8 FILLER_70_637 ();
 sg13g2_decap_8 FILLER_70_644 ();
 sg13g2_decap_8 FILLER_70_651 ();
 sg13g2_decap_8 FILLER_70_658 ();
 sg13g2_decap_8 FILLER_70_665 ();
 sg13g2_decap_8 FILLER_70_672 ();
 sg13g2_decap_8 FILLER_70_679 ();
 sg13g2_decap_8 FILLER_70_686 ();
 sg13g2_decap_8 FILLER_70_693 ();
 sg13g2_decap_8 FILLER_70_700 ();
 sg13g2_decap_8 FILLER_70_707 ();
 sg13g2_decap_8 FILLER_70_714 ();
 sg13g2_decap_8 FILLER_70_721 ();
 sg13g2_decap_8 FILLER_70_728 ();
 sg13g2_decap_8 FILLER_70_735 ();
 sg13g2_decap_8 FILLER_70_742 ();
 sg13g2_decap_8 FILLER_70_749 ();
 sg13g2_decap_8 FILLER_70_756 ();
 sg13g2_decap_8 FILLER_70_763 ();
 sg13g2_decap_8 FILLER_70_770 ();
 sg13g2_decap_8 FILLER_70_777 ();
 sg13g2_decap_8 FILLER_70_784 ();
 sg13g2_decap_8 FILLER_70_791 ();
 sg13g2_decap_8 FILLER_70_798 ();
 sg13g2_decap_8 FILLER_70_805 ();
 sg13g2_decap_8 FILLER_70_812 ();
 sg13g2_decap_8 FILLER_70_819 ();
 sg13g2_decap_8 FILLER_70_826 ();
 sg13g2_decap_8 FILLER_70_833 ();
 sg13g2_fill_1 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_decap_8 FILLER_71_182 ();
 sg13g2_decap_8 FILLER_71_189 ();
 sg13g2_decap_8 FILLER_71_196 ();
 sg13g2_decap_8 FILLER_71_203 ();
 sg13g2_decap_8 FILLER_71_210 ();
 sg13g2_decap_8 FILLER_71_217 ();
 sg13g2_decap_8 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_231 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_245 ();
 sg13g2_decap_8 FILLER_71_252 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_decap_8 FILLER_71_266 ();
 sg13g2_decap_8 FILLER_71_273 ();
 sg13g2_decap_8 FILLER_71_280 ();
 sg13g2_decap_8 FILLER_71_287 ();
 sg13g2_decap_8 FILLER_71_294 ();
 sg13g2_decap_8 FILLER_71_301 ();
 sg13g2_decap_8 FILLER_71_308 ();
 sg13g2_decap_8 FILLER_71_315 ();
 sg13g2_decap_8 FILLER_71_322 ();
 sg13g2_decap_8 FILLER_71_329 ();
 sg13g2_decap_8 FILLER_71_336 ();
 sg13g2_decap_8 FILLER_71_343 ();
 sg13g2_decap_8 FILLER_71_350 ();
 sg13g2_decap_8 FILLER_71_357 ();
 sg13g2_decap_8 FILLER_71_364 ();
 sg13g2_decap_8 FILLER_71_371 ();
 sg13g2_decap_8 FILLER_71_378 ();
 sg13g2_decap_8 FILLER_71_385 ();
 sg13g2_decap_8 FILLER_71_392 ();
 sg13g2_decap_8 FILLER_71_399 ();
 sg13g2_decap_8 FILLER_71_406 ();
 sg13g2_decap_8 FILLER_71_413 ();
 sg13g2_decap_8 FILLER_71_420 ();
 sg13g2_decap_8 FILLER_71_427 ();
 sg13g2_decap_8 FILLER_71_434 ();
 sg13g2_decap_8 FILLER_71_441 ();
 sg13g2_decap_8 FILLER_71_448 ();
 sg13g2_decap_8 FILLER_71_455 ();
 sg13g2_decap_8 FILLER_71_462 ();
 sg13g2_decap_8 FILLER_71_469 ();
 sg13g2_decap_8 FILLER_71_476 ();
 sg13g2_decap_8 FILLER_71_483 ();
 sg13g2_decap_8 FILLER_71_490 ();
 sg13g2_decap_8 FILLER_71_497 ();
 sg13g2_decap_8 FILLER_71_504 ();
 sg13g2_decap_8 FILLER_71_511 ();
 sg13g2_decap_8 FILLER_71_518 ();
 sg13g2_decap_8 FILLER_71_525 ();
 sg13g2_decap_8 FILLER_71_532 ();
 sg13g2_decap_8 FILLER_71_539 ();
 sg13g2_decap_8 FILLER_71_546 ();
 sg13g2_decap_8 FILLER_71_553 ();
 sg13g2_decap_8 FILLER_71_560 ();
 sg13g2_decap_8 FILLER_71_567 ();
 sg13g2_decap_8 FILLER_71_574 ();
 sg13g2_decap_8 FILLER_71_581 ();
 sg13g2_decap_8 FILLER_71_588 ();
 sg13g2_decap_8 FILLER_71_595 ();
 sg13g2_decap_8 FILLER_71_602 ();
 sg13g2_decap_8 FILLER_71_609 ();
 sg13g2_decap_8 FILLER_71_616 ();
 sg13g2_decap_8 FILLER_71_623 ();
 sg13g2_decap_8 FILLER_71_630 ();
 sg13g2_decap_8 FILLER_71_637 ();
 sg13g2_decap_8 FILLER_71_644 ();
 sg13g2_decap_8 FILLER_71_651 ();
 sg13g2_decap_8 FILLER_71_658 ();
 sg13g2_decap_8 FILLER_71_665 ();
 sg13g2_decap_8 FILLER_71_672 ();
 sg13g2_decap_8 FILLER_71_679 ();
 sg13g2_decap_8 FILLER_71_686 ();
 sg13g2_decap_8 FILLER_71_693 ();
 sg13g2_decap_8 FILLER_71_700 ();
 sg13g2_decap_8 FILLER_71_707 ();
 sg13g2_decap_8 FILLER_71_714 ();
 sg13g2_decap_8 FILLER_71_721 ();
 sg13g2_decap_8 FILLER_71_728 ();
 sg13g2_decap_8 FILLER_71_735 ();
 sg13g2_decap_8 FILLER_71_742 ();
 sg13g2_decap_8 FILLER_71_749 ();
 sg13g2_decap_8 FILLER_71_756 ();
 sg13g2_decap_8 FILLER_71_763 ();
 sg13g2_decap_8 FILLER_71_770 ();
 sg13g2_decap_8 FILLER_71_777 ();
 sg13g2_decap_8 FILLER_71_784 ();
 sg13g2_decap_8 FILLER_71_791 ();
 sg13g2_decap_8 FILLER_71_798 ();
 sg13g2_decap_8 FILLER_71_805 ();
 sg13g2_decap_8 FILLER_71_812 ();
 sg13g2_decap_8 FILLER_71_819 ();
 sg13g2_decap_8 FILLER_71_826 ();
 sg13g2_decap_8 FILLER_71_833 ();
 sg13g2_fill_1 FILLER_71_840 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_decap_8 FILLER_72_182 ();
 sg13g2_decap_8 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_decap_8 FILLER_72_238 ();
 sg13g2_decap_8 FILLER_72_245 ();
 sg13g2_decap_8 FILLER_72_252 ();
 sg13g2_decap_8 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_266 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_decap_8 FILLER_72_280 ();
 sg13g2_decap_8 FILLER_72_287 ();
 sg13g2_decap_8 FILLER_72_294 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_308 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_decap_8 FILLER_72_322 ();
 sg13g2_decap_8 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_336 ();
 sg13g2_decap_8 FILLER_72_343 ();
 sg13g2_decap_8 FILLER_72_350 ();
 sg13g2_decap_8 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_decap_8 FILLER_72_406 ();
 sg13g2_decap_8 FILLER_72_413 ();
 sg13g2_decap_8 FILLER_72_420 ();
 sg13g2_decap_8 FILLER_72_427 ();
 sg13g2_decap_8 FILLER_72_434 ();
 sg13g2_decap_8 FILLER_72_441 ();
 sg13g2_decap_8 FILLER_72_448 ();
 sg13g2_decap_8 FILLER_72_455 ();
 sg13g2_decap_8 FILLER_72_462 ();
 sg13g2_decap_8 FILLER_72_469 ();
 sg13g2_decap_8 FILLER_72_476 ();
 sg13g2_decap_8 FILLER_72_483 ();
 sg13g2_decap_8 FILLER_72_490 ();
 sg13g2_decap_8 FILLER_72_497 ();
 sg13g2_decap_8 FILLER_72_504 ();
 sg13g2_decap_8 FILLER_72_511 ();
 sg13g2_decap_8 FILLER_72_518 ();
 sg13g2_decap_8 FILLER_72_525 ();
 sg13g2_decap_8 FILLER_72_532 ();
 sg13g2_decap_8 FILLER_72_539 ();
 sg13g2_decap_8 FILLER_72_546 ();
 sg13g2_decap_8 FILLER_72_553 ();
 sg13g2_decap_8 FILLER_72_560 ();
 sg13g2_decap_8 FILLER_72_567 ();
 sg13g2_decap_8 FILLER_72_574 ();
 sg13g2_decap_8 FILLER_72_581 ();
 sg13g2_decap_8 FILLER_72_588 ();
 sg13g2_decap_8 FILLER_72_595 ();
 sg13g2_decap_8 FILLER_72_602 ();
 sg13g2_decap_8 FILLER_72_609 ();
 sg13g2_decap_8 FILLER_72_616 ();
 sg13g2_decap_8 FILLER_72_623 ();
 sg13g2_decap_8 FILLER_72_630 ();
 sg13g2_decap_8 FILLER_72_637 ();
 sg13g2_decap_8 FILLER_72_644 ();
 sg13g2_decap_8 FILLER_72_651 ();
 sg13g2_decap_8 FILLER_72_658 ();
 sg13g2_decap_8 FILLER_72_665 ();
 sg13g2_decap_8 FILLER_72_672 ();
 sg13g2_decap_8 FILLER_72_679 ();
 sg13g2_decap_8 FILLER_72_686 ();
 sg13g2_decap_8 FILLER_72_693 ();
 sg13g2_decap_8 FILLER_72_700 ();
 sg13g2_decap_8 FILLER_72_707 ();
 sg13g2_decap_8 FILLER_72_714 ();
 sg13g2_decap_8 FILLER_72_721 ();
 sg13g2_decap_8 FILLER_72_728 ();
 sg13g2_decap_8 FILLER_72_735 ();
 sg13g2_decap_8 FILLER_72_742 ();
 sg13g2_decap_8 FILLER_72_749 ();
 sg13g2_decap_8 FILLER_72_756 ();
 sg13g2_decap_8 FILLER_72_763 ();
 sg13g2_decap_8 FILLER_72_770 ();
 sg13g2_decap_8 FILLER_72_777 ();
 sg13g2_decap_8 FILLER_72_784 ();
 sg13g2_decap_8 FILLER_72_791 ();
 sg13g2_decap_8 FILLER_72_798 ();
 sg13g2_decap_8 FILLER_72_805 ();
 sg13g2_decap_8 FILLER_72_812 ();
 sg13g2_decap_8 FILLER_72_819 ();
 sg13g2_decap_8 FILLER_72_826 ();
 sg13g2_decap_8 FILLER_72_833 ();
 sg13g2_fill_1 FILLER_72_840 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_8 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_189 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_decap_8 FILLER_73_217 ();
 sg13g2_decap_8 FILLER_73_224 ();
 sg13g2_decap_8 FILLER_73_231 ();
 sg13g2_decap_8 FILLER_73_238 ();
 sg13g2_decap_8 FILLER_73_245 ();
 sg13g2_decap_8 FILLER_73_252 ();
 sg13g2_decap_8 FILLER_73_259 ();
 sg13g2_decap_8 FILLER_73_266 ();
 sg13g2_decap_8 FILLER_73_273 ();
 sg13g2_decap_8 FILLER_73_280 ();
 sg13g2_decap_8 FILLER_73_287 ();
 sg13g2_decap_8 FILLER_73_294 ();
 sg13g2_decap_8 FILLER_73_301 ();
 sg13g2_decap_8 FILLER_73_308 ();
 sg13g2_decap_8 FILLER_73_315 ();
 sg13g2_decap_8 FILLER_73_322 ();
 sg13g2_decap_8 FILLER_73_329 ();
 sg13g2_decap_8 FILLER_73_336 ();
 sg13g2_decap_8 FILLER_73_343 ();
 sg13g2_decap_8 FILLER_73_350 ();
 sg13g2_decap_8 FILLER_73_357 ();
 sg13g2_decap_8 FILLER_73_364 ();
 sg13g2_decap_8 FILLER_73_371 ();
 sg13g2_decap_8 FILLER_73_378 ();
 sg13g2_decap_8 FILLER_73_385 ();
 sg13g2_decap_8 FILLER_73_392 ();
 sg13g2_decap_8 FILLER_73_399 ();
 sg13g2_decap_8 FILLER_73_406 ();
 sg13g2_decap_8 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_420 ();
 sg13g2_decap_8 FILLER_73_427 ();
 sg13g2_decap_8 FILLER_73_434 ();
 sg13g2_decap_8 FILLER_73_441 ();
 sg13g2_decap_8 FILLER_73_448 ();
 sg13g2_decap_8 FILLER_73_455 ();
 sg13g2_decap_8 FILLER_73_462 ();
 sg13g2_decap_8 FILLER_73_469 ();
 sg13g2_decap_8 FILLER_73_476 ();
 sg13g2_decap_8 FILLER_73_483 ();
 sg13g2_decap_8 FILLER_73_490 ();
 sg13g2_decap_8 FILLER_73_497 ();
 sg13g2_decap_8 FILLER_73_504 ();
 sg13g2_decap_8 FILLER_73_511 ();
 sg13g2_decap_8 FILLER_73_518 ();
 sg13g2_decap_8 FILLER_73_525 ();
 sg13g2_decap_8 FILLER_73_532 ();
 sg13g2_decap_8 FILLER_73_539 ();
 sg13g2_decap_8 FILLER_73_546 ();
 sg13g2_decap_8 FILLER_73_553 ();
 sg13g2_decap_8 FILLER_73_560 ();
 sg13g2_decap_8 FILLER_73_567 ();
 sg13g2_decap_8 FILLER_73_574 ();
 sg13g2_decap_8 FILLER_73_581 ();
 sg13g2_decap_8 FILLER_73_588 ();
 sg13g2_decap_8 FILLER_73_595 ();
 sg13g2_decap_8 FILLER_73_602 ();
 sg13g2_decap_8 FILLER_73_609 ();
 sg13g2_decap_8 FILLER_73_616 ();
 sg13g2_decap_8 FILLER_73_623 ();
 sg13g2_decap_8 FILLER_73_630 ();
 sg13g2_decap_8 FILLER_73_637 ();
 sg13g2_decap_8 FILLER_73_644 ();
 sg13g2_decap_8 FILLER_73_651 ();
 sg13g2_decap_8 FILLER_73_658 ();
 sg13g2_decap_8 FILLER_73_665 ();
 sg13g2_decap_8 FILLER_73_672 ();
 sg13g2_decap_8 FILLER_73_679 ();
 sg13g2_decap_8 FILLER_73_686 ();
 sg13g2_decap_8 FILLER_73_693 ();
 sg13g2_decap_8 FILLER_73_700 ();
 sg13g2_decap_8 FILLER_73_707 ();
 sg13g2_decap_8 FILLER_73_714 ();
 sg13g2_decap_8 FILLER_73_721 ();
 sg13g2_decap_8 FILLER_73_728 ();
 sg13g2_decap_8 FILLER_73_735 ();
 sg13g2_decap_8 FILLER_73_742 ();
 sg13g2_decap_8 FILLER_73_749 ();
 sg13g2_decap_8 FILLER_73_756 ();
 sg13g2_decap_8 FILLER_73_763 ();
 sg13g2_decap_8 FILLER_73_770 ();
 sg13g2_decap_8 FILLER_73_777 ();
 sg13g2_decap_8 FILLER_73_784 ();
 sg13g2_decap_8 FILLER_73_791 ();
 sg13g2_decap_8 FILLER_73_798 ();
 sg13g2_decap_8 FILLER_73_805 ();
 sg13g2_decap_8 FILLER_73_812 ();
 sg13g2_decap_8 FILLER_73_819 ();
 sg13g2_decap_8 FILLER_73_826 ();
 sg13g2_decap_8 FILLER_73_833 ();
 sg13g2_fill_1 FILLER_73_840 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_8 FILLER_74_175 ();
 sg13g2_decap_8 FILLER_74_182 ();
 sg13g2_decap_8 FILLER_74_189 ();
 sg13g2_decap_8 FILLER_74_196 ();
 sg13g2_decap_8 FILLER_74_203 ();
 sg13g2_decap_8 FILLER_74_210 ();
 sg13g2_decap_8 FILLER_74_217 ();
 sg13g2_decap_8 FILLER_74_224 ();
 sg13g2_decap_8 FILLER_74_231 ();
 sg13g2_decap_8 FILLER_74_238 ();
 sg13g2_decap_8 FILLER_74_245 ();
 sg13g2_decap_8 FILLER_74_252 ();
 sg13g2_decap_8 FILLER_74_259 ();
 sg13g2_decap_8 FILLER_74_266 ();
 sg13g2_decap_8 FILLER_74_273 ();
 sg13g2_decap_8 FILLER_74_280 ();
 sg13g2_decap_8 FILLER_74_287 ();
 sg13g2_decap_8 FILLER_74_294 ();
 sg13g2_decap_8 FILLER_74_301 ();
 sg13g2_decap_8 FILLER_74_308 ();
 sg13g2_decap_8 FILLER_74_315 ();
 sg13g2_decap_8 FILLER_74_322 ();
 sg13g2_decap_8 FILLER_74_329 ();
 sg13g2_decap_8 FILLER_74_336 ();
 sg13g2_decap_8 FILLER_74_343 ();
 sg13g2_decap_8 FILLER_74_350 ();
 sg13g2_decap_8 FILLER_74_357 ();
 sg13g2_decap_8 FILLER_74_364 ();
 sg13g2_decap_8 FILLER_74_371 ();
 sg13g2_decap_8 FILLER_74_378 ();
 sg13g2_decap_8 FILLER_74_385 ();
 sg13g2_decap_8 FILLER_74_392 ();
 sg13g2_decap_8 FILLER_74_399 ();
 sg13g2_decap_8 FILLER_74_406 ();
 sg13g2_decap_8 FILLER_74_413 ();
 sg13g2_decap_8 FILLER_74_420 ();
 sg13g2_decap_8 FILLER_74_427 ();
 sg13g2_decap_8 FILLER_74_434 ();
 sg13g2_decap_8 FILLER_74_441 ();
 sg13g2_decap_8 FILLER_74_448 ();
 sg13g2_decap_8 FILLER_74_455 ();
 sg13g2_decap_8 FILLER_74_462 ();
 sg13g2_decap_8 FILLER_74_469 ();
 sg13g2_decap_8 FILLER_74_476 ();
 sg13g2_decap_8 FILLER_74_483 ();
 sg13g2_decap_8 FILLER_74_490 ();
 sg13g2_decap_8 FILLER_74_497 ();
 sg13g2_decap_8 FILLER_74_504 ();
 sg13g2_decap_8 FILLER_74_511 ();
 sg13g2_decap_8 FILLER_74_518 ();
 sg13g2_decap_8 FILLER_74_525 ();
 sg13g2_decap_8 FILLER_74_532 ();
 sg13g2_decap_8 FILLER_74_539 ();
 sg13g2_decap_8 FILLER_74_546 ();
 sg13g2_decap_8 FILLER_74_553 ();
 sg13g2_decap_8 FILLER_74_560 ();
 sg13g2_decap_8 FILLER_74_567 ();
 sg13g2_decap_8 FILLER_74_574 ();
 sg13g2_decap_8 FILLER_74_581 ();
 sg13g2_decap_8 FILLER_74_588 ();
 sg13g2_decap_8 FILLER_74_595 ();
 sg13g2_decap_8 FILLER_74_602 ();
 sg13g2_decap_8 FILLER_74_609 ();
 sg13g2_decap_8 FILLER_74_616 ();
 sg13g2_decap_8 FILLER_74_623 ();
 sg13g2_decap_8 FILLER_74_630 ();
 sg13g2_decap_8 FILLER_74_637 ();
 sg13g2_decap_8 FILLER_74_644 ();
 sg13g2_decap_8 FILLER_74_651 ();
 sg13g2_decap_8 FILLER_74_658 ();
 sg13g2_decap_8 FILLER_74_665 ();
 sg13g2_decap_8 FILLER_74_672 ();
 sg13g2_decap_8 FILLER_74_679 ();
 sg13g2_decap_8 FILLER_74_686 ();
 sg13g2_decap_8 FILLER_74_693 ();
 sg13g2_decap_8 FILLER_74_700 ();
 sg13g2_decap_8 FILLER_74_707 ();
 sg13g2_decap_8 FILLER_74_714 ();
 sg13g2_decap_8 FILLER_74_721 ();
 sg13g2_decap_8 FILLER_74_728 ();
 sg13g2_decap_8 FILLER_74_735 ();
 sg13g2_decap_8 FILLER_74_742 ();
 sg13g2_decap_8 FILLER_74_749 ();
 sg13g2_decap_8 FILLER_74_756 ();
 sg13g2_decap_8 FILLER_74_763 ();
 sg13g2_decap_8 FILLER_74_770 ();
 sg13g2_decap_8 FILLER_74_777 ();
 sg13g2_decap_8 FILLER_74_784 ();
 sg13g2_decap_8 FILLER_74_791 ();
 sg13g2_decap_8 FILLER_74_798 ();
 sg13g2_decap_8 FILLER_74_805 ();
 sg13g2_decap_8 FILLER_74_812 ();
 sg13g2_decap_8 FILLER_74_819 ();
 sg13g2_decap_8 FILLER_74_826 ();
 sg13g2_decap_8 FILLER_74_833 ();
 sg13g2_fill_1 FILLER_74_840 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_decap_8 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_75_329 ();
 sg13g2_decap_8 FILLER_75_336 ();
 sg13g2_decap_8 FILLER_75_343 ();
 sg13g2_decap_8 FILLER_75_350 ();
 sg13g2_decap_8 FILLER_75_357 ();
 sg13g2_decap_8 FILLER_75_364 ();
 sg13g2_decap_8 FILLER_75_371 ();
 sg13g2_decap_8 FILLER_75_378 ();
 sg13g2_decap_8 FILLER_75_385 ();
 sg13g2_decap_8 FILLER_75_392 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_decap_8 FILLER_75_406 ();
 sg13g2_decap_8 FILLER_75_413 ();
 sg13g2_decap_8 FILLER_75_420 ();
 sg13g2_decap_8 FILLER_75_427 ();
 sg13g2_decap_8 FILLER_75_434 ();
 sg13g2_decap_8 FILLER_75_441 ();
 sg13g2_decap_8 FILLER_75_448 ();
 sg13g2_decap_8 FILLER_75_455 ();
 sg13g2_decap_8 FILLER_75_462 ();
 sg13g2_decap_8 FILLER_75_469 ();
 sg13g2_decap_8 FILLER_75_476 ();
 sg13g2_decap_8 FILLER_75_483 ();
 sg13g2_decap_8 FILLER_75_490 ();
 sg13g2_decap_8 FILLER_75_497 ();
 sg13g2_decap_8 FILLER_75_504 ();
 sg13g2_decap_8 FILLER_75_511 ();
 sg13g2_decap_8 FILLER_75_518 ();
 sg13g2_decap_8 FILLER_75_525 ();
 sg13g2_decap_8 FILLER_75_532 ();
 sg13g2_decap_8 FILLER_75_539 ();
 sg13g2_decap_8 FILLER_75_546 ();
 sg13g2_decap_8 FILLER_75_553 ();
 sg13g2_decap_8 FILLER_75_560 ();
 sg13g2_decap_8 FILLER_75_567 ();
 sg13g2_decap_8 FILLER_75_574 ();
 sg13g2_decap_8 FILLER_75_581 ();
 sg13g2_decap_8 FILLER_75_588 ();
 sg13g2_decap_8 FILLER_75_595 ();
 sg13g2_decap_8 FILLER_75_602 ();
 sg13g2_decap_8 FILLER_75_609 ();
 sg13g2_decap_8 FILLER_75_616 ();
 sg13g2_decap_8 FILLER_75_623 ();
 sg13g2_decap_8 FILLER_75_630 ();
 sg13g2_decap_8 FILLER_75_637 ();
 sg13g2_decap_8 FILLER_75_644 ();
 sg13g2_decap_8 FILLER_75_651 ();
 sg13g2_decap_8 FILLER_75_658 ();
 sg13g2_decap_8 FILLER_75_665 ();
 sg13g2_decap_8 FILLER_75_672 ();
 sg13g2_decap_8 FILLER_75_679 ();
 sg13g2_decap_8 FILLER_75_686 ();
 sg13g2_decap_8 FILLER_75_693 ();
 sg13g2_decap_8 FILLER_75_700 ();
 sg13g2_decap_8 FILLER_75_707 ();
 sg13g2_decap_8 FILLER_75_714 ();
 sg13g2_decap_8 FILLER_75_721 ();
 sg13g2_decap_8 FILLER_75_728 ();
 sg13g2_decap_8 FILLER_75_735 ();
 sg13g2_decap_8 FILLER_75_742 ();
 sg13g2_decap_8 FILLER_75_749 ();
 sg13g2_decap_8 FILLER_75_756 ();
 sg13g2_decap_8 FILLER_75_763 ();
 sg13g2_decap_8 FILLER_75_770 ();
 sg13g2_decap_8 FILLER_75_777 ();
 sg13g2_decap_8 FILLER_75_784 ();
 sg13g2_decap_8 FILLER_75_791 ();
 sg13g2_decap_8 FILLER_75_798 ();
 sg13g2_decap_8 FILLER_75_805 ();
 sg13g2_decap_8 FILLER_75_812 ();
 sg13g2_decap_8 FILLER_75_819 ();
 sg13g2_decap_8 FILLER_75_826 ();
 sg13g2_decap_8 FILLER_75_833 ();
 sg13g2_fill_1 FILLER_75_840 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_203 ();
 sg13g2_decap_8 FILLER_76_210 ();
 sg13g2_decap_8 FILLER_76_217 ();
 sg13g2_decap_8 FILLER_76_224 ();
 sg13g2_decap_8 FILLER_76_231 ();
 sg13g2_decap_8 FILLER_76_238 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_decap_8 FILLER_76_266 ();
 sg13g2_decap_8 FILLER_76_273 ();
 sg13g2_decap_8 FILLER_76_280 ();
 sg13g2_decap_8 FILLER_76_287 ();
 sg13g2_decap_8 FILLER_76_294 ();
 sg13g2_decap_8 FILLER_76_301 ();
 sg13g2_decap_8 FILLER_76_308 ();
 sg13g2_decap_8 FILLER_76_315 ();
 sg13g2_decap_8 FILLER_76_322 ();
 sg13g2_decap_8 FILLER_76_329 ();
 sg13g2_decap_8 FILLER_76_336 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_8 FILLER_76_357 ();
 sg13g2_decap_8 FILLER_76_364 ();
 sg13g2_decap_8 FILLER_76_371 ();
 sg13g2_decap_8 FILLER_76_378 ();
 sg13g2_decap_8 FILLER_76_385 ();
 sg13g2_decap_8 FILLER_76_392 ();
 sg13g2_decap_8 FILLER_76_399 ();
 sg13g2_decap_8 FILLER_76_406 ();
 sg13g2_decap_8 FILLER_76_413 ();
 sg13g2_decap_8 FILLER_76_420 ();
 sg13g2_decap_8 FILLER_76_427 ();
 sg13g2_decap_8 FILLER_76_434 ();
 sg13g2_decap_8 FILLER_76_441 ();
 sg13g2_decap_8 FILLER_76_448 ();
 sg13g2_decap_8 FILLER_76_455 ();
 sg13g2_decap_8 FILLER_76_462 ();
 sg13g2_decap_8 FILLER_76_469 ();
 sg13g2_decap_8 FILLER_76_476 ();
 sg13g2_decap_8 FILLER_76_483 ();
 sg13g2_decap_8 FILLER_76_490 ();
 sg13g2_decap_8 FILLER_76_497 ();
 sg13g2_decap_8 FILLER_76_504 ();
 sg13g2_decap_8 FILLER_76_511 ();
 sg13g2_decap_8 FILLER_76_518 ();
 sg13g2_decap_8 FILLER_76_525 ();
 sg13g2_decap_8 FILLER_76_532 ();
 sg13g2_decap_8 FILLER_76_539 ();
 sg13g2_decap_8 FILLER_76_546 ();
 sg13g2_decap_8 FILLER_76_553 ();
 sg13g2_decap_8 FILLER_76_560 ();
 sg13g2_decap_8 FILLER_76_567 ();
 sg13g2_decap_8 FILLER_76_574 ();
 sg13g2_decap_8 FILLER_76_581 ();
 sg13g2_decap_8 FILLER_76_588 ();
 sg13g2_decap_8 FILLER_76_595 ();
 sg13g2_decap_8 FILLER_76_602 ();
 sg13g2_decap_8 FILLER_76_609 ();
 sg13g2_decap_8 FILLER_76_616 ();
 sg13g2_decap_8 FILLER_76_623 ();
 sg13g2_decap_8 FILLER_76_630 ();
 sg13g2_decap_8 FILLER_76_637 ();
 sg13g2_decap_8 FILLER_76_644 ();
 sg13g2_decap_8 FILLER_76_651 ();
 sg13g2_decap_8 FILLER_76_658 ();
 sg13g2_decap_8 FILLER_76_665 ();
 sg13g2_decap_8 FILLER_76_672 ();
 sg13g2_decap_8 FILLER_76_679 ();
 sg13g2_decap_8 FILLER_76_686 ();
 sg13g2_decap_8 FILLER_76_693 ();
 sg13g2_decap_8 FILLER_76_700 ();
 sg13g2_decap_8 FILLER_76_707 ();
 sg13g2_decap_8 FILLER_76_714 ();
 sg13g2_decap_8 FILLER_76_721 ();
 sg13g2_decap_8 FILLER_76_728 ();
 sg13g2_decap_8 FILLER_76_735 ();
 sg13g2_decap_8 FILLER_76_742 ();
 sg13g2_decap_8 FILLER_76_749 ();
 sg13g2_decap_8 FILLER_76_756 ();
 sg13g2_decap_8 FILLER_76_763 ();
 sg13g2_decap_8 FILLER_76_770 ();
 sg13g2_decap_8 FILLER_76_777 ();
 sg13g2_decap_8 FILLER_76_784 ();
 sg13g2_decap_8 FILLER_76_791 ();
 sg13g2_decap_8 FILLER_76_798 ();
 sg13g2_decap_8 FILLER_76_805 ();
 sg13g2_decap_8 FILLER_76_812 ();
 sg13g2_decap_8 FILLER_76_819 ();
 sg13g2_decap_8 FILLER_76_826 ();
 sg13g2_decap_8 FILLER_76_833 ();
 sg13g2_fill_1 FILLER_76_840 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_441 ();
 sg13g2_decap_8 FILLER_77_448 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_decap_8 FILLER_77_462 ();
 sg13g2_decap_8 FILLER_77_469 ();
 sg13g2_decap_8 FILLER_77_476 ();
 sg13g2_decap_8 FILLER_77_483 ();
 sg13g2_decap_8 FILLER_77_490 ();
 sg13g2_decap_8 FILLER_77_497 ();
 sg13g2_decap_8 FILLER_77_504 ();
 sg13g2_decap_8 FILLER_77_511 ();
 sg13g2_decap_8 FILLER_77_518 ();
 sg13g2_decap_8 FILLER_77_525 ();
 sg13g2_decap_8 FILLER_77_532 ();
 sg13g2_decap_8 FILLER_77_539 ();
 sg13g2_decap_8 FILLER_77_546 ();
 sg13g2_decap_8 FILLER_77_553 ();
 sg13g2_decap_8 FILLER_77_560 ();
 sg13g2_decap_8 FILLER_77_567 ();
 sg13g2_decap_8 FILLER_77_574 ();
 sg13g2_decap_8 FILLER_77_581 ();
 sg13g2_decap_8 FILLER_77_588 ();
 sg13g2_decap_8 FILLER_77_595 ();
 sg13g2_decap_8 FILLER_77_602 ();
 sg13g2_decap_8 FILLER_77_609 ();
 sg13g2_decap_8 FILLER_77_616 ();
 sg13g2_decap_8 FILLER_77_623 ();
 sg13g2_decap_8 FILLER_77_630 ();
 sg13g2_decap_8 FILLER_77_637 ();
 sg13g2_decap_8 FILLER_77_644 ();
 sg13g2_decap_8 FILLER_77_651 ();
 sg13g2_decap_8 FILLER_77_658 ();
 sg13g2_decap_8 FILLER_77_665 ();
 sg13g2_decap_8 FILLER_77_672 ();
 sg13g2_decap_8 FILLER_77_679 ();
 sg13g2_decap_8 FILLER_77_686 ();
 sg13g2_decap_8 FILLER_77_693 ();
 sg13g2_decap_8 FILLER_77_700 ();
 sg13g2_decap_8 FILLER_77_707 ();
 sg13g2_decap_8 FILLER_77_714 ();
 sg13g2_decap_8 FILLER_77_721 ();
 sg13g2_decap_8 FILLER_77_728 ();
 sg13g2_decap_8 FILLER_77_735 ();
 sg13g2_decap_8 FILLER_77_742 ();
 sg13g2_decap_8 FILLER_77_749 ();
 sg13g2_decap_8 FILLER_77_756 ();
 sg13g2_decap_8 FILLER_77_763 ();
 sg13g2_decap_8 FILLER_77_770 ();
 sg13g2_decap_8 FILLER_77_777 ();
 sg13g2_decap_8 FILLER_77_784 ();
 sg13g2_decap_8 FILLER_77_791 ();
 sg13g2_decap_8 FILLER_77_798 ();
 sg13g2_decap_8 FILLER_77_805 ();
 sg13g2_decap_8 FILLER_77_812 ();
 sg13g2_decap_8 FILLER_77_819 ();
 sg13g2_decap_8 FILLER_77_826 ();
 sg13g2_decap_8 FILLER_77_833 ();
 sg13g2_fill_1 FILLER_77_840 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_decap_8 FILLER_78_84 ();
 sg13g2_decap_8 FILLER_78_91 ();
 sg13g2_decap_8 FILLER_78_98 ();
 sg13g2_decap_8 FILLER_78_105 ();
 sg13g2_decap_8 FILLER_78_112 ();
 sg13g2_decap_8 FILLER_78_119 ();
 sg13g2_decap_8 FILLER_78_126 ();
 sg13g2_decap_8 FILLER_78_133 ();
 sg13g2_decap_8 FILLER_78_140 ();
 sg13g2_decap_8 FILLER_78_147 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_161 ();
 sg13g2_decap_8 FILLER_78_168 ();
 sg13g2_decap_8 FILLER_78_175 ();
 sg13g2_decap_8 FILLER_78_182 ();
 sg13g2_decap_8 FILLER_78_189 ();
 sg13g2_decap_8 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_203 ();
 sg13g2_decap_8 FILLER_78_210 ();
 sg13g2_decap_8 FILLER_78_217 ();
 sg13g2_decap_8 FILLER_78_224 ();
 sg13g2_decap_8 FILLER_78_231 ();
 sg13g2_decap_8 FILLER_78_238 ();
 sg13g2_decap_8 FILLER_78_245 ();
 sg13g2_decap_8 FILLER_78_252 ();
 sg13g2_decap_8 FILLER_78_259 ();
 sg13g2_decap_8 FILLER_78_266 ();
 sg13g2_decap_8 FILLER_78_273 ();
 sg13g2_decap_8 FILLER_78_280 ();
 sg13g2_decap_8 FILLER_78_287 ();
 sg13g2_decap_8 FILLER_78_294 ();
 sg13g2_decap_8 FILLER_78_301 ();
 sg13g2_decap_8 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_315 ();
 sg13g2_decap_8 FILLER_78_322 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_8 FILLER_78_350 ();
 sg13g2_decap_8 FILLER_78_357 ();
 sg13g2_decap_8 FILLER_78_364 ();
 sg13g2_decap_8 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_385 ();
 sg13g2_decap_8 FILLER_78_392 ();
 sg13g2_decap_8 FILLER_78_399 ();
 sg13g2_decap_8 FILLER_78_406 ();
 sg13g2_decap_8 FILLER_78_413 ();
 sg13g2_decap_8 FILLER_78_420 ();
 sg13g2_decap_8 FILLER_78_427 ();
 sg13g2_decap_8 FILLER_78_434 ();
 sg13g2_decap_8 FILLER_78_441 ();
 sg13g2_decap_8 FILLER_78_448 ();
 sg13g2_decap_8 FILLER_78_455 ();
 sg13g2_decap_8 FILLER_78_462 ();
 sg13g2_decap_8 FILLER_78_469 ();
 sg13g2_decap_8 FILLER_78_476 ();
 sg13g2_decap_8 FILLER_78_483 ();
 sg13g2_decap_8 FILLER_78_490 ();
 sg13g2_decap_8 FILLER_78_497 ();
 sg13g2_decap_8 FILLER_78_504 ();
 sg13g2_decap_8 FILLER_78_511 ();
 sg13g2_decap_8 FILLER_78_518 ();
 sg13g2_decap_8 FILLER_78_525 ();
 sg13g2_decap_8 FILLER_78_532 ();
 sg13g2_decap_8 FILLER_78_539 ();
 sg13g2_decap_8 FILLER_78_546 ();
 sg13g2_decap_8 FILLER_78_553 ();
 sg13g2_decap_8 FILLER_78_560 ();
 sg13g2_decap_8 FILLER_78_567 ();
 sg13g2_decap_8 FILLER_78_574 ();
 sg13g2_decap_8 FILLER_78_581 ();
 sg13g2_decap_8 FILLER_78_588 ();
 sg13g2_decap_8 FILLER_78_595 ();
 sg13g2_decap_8 FILLER_78_602 ();
 sg13g2_decap_8 FILLER_78_609 ();
 sg13g2_decap_8 FILLER_78_616 ();
 sg13g2_decap_8 FILLER_78_623 ();
 sg13g2_decap_8 FILLER_78_630 ();
 sg13g2_decap_8 FILLER_78_637 ();
 sg13g2_decap_8 FILLER_78_644 ();
 sg13g2_decap_8 FILLER_78_651 ();
 sg13g2_decap_8 FILLER_78_658 ();
 sg13g2_decap_8 FILLER_78_665 ();
 sg13g2_decap_8 FILLER_78_672 ();
 sg13g2_decap_8 FILLER_78_679 ();
 sg13g2_decap_8 FILLER_78_686 ();
 sg13g2_decap_8 FILLER_78_693 ();
 sg13g2_decap_8 FILLER_78_700 ();
 sg13g2_decap_8 FILLER_78_707 ();
 sg13g2_decap_8 FILLER_78_714 ();
 sg13g2_decap_8 FILLER_78_721 ();
 sg13g2_decap_8 FILLER_78_728 ();
 sg13g2_decap_8 FILLER_78_735 ();
 sg13g2_decap_8 FILLER_78_742 ();
 sg13g2_decap_8 FILLER_78_749 ();
 sg13g2_decap_8 FILLER_78_756 ();
 sg13g2_decap_8 FILLER_78_763 ();
 sg13g2_decap_8 FILLER_78_770 ();
 sg13g2_decap_8 FILLER_78_777 ();
 sg13g2_decap_8 FILLER_78_784 ();
 sg13g2_decap_8 FILLER_78_791 ();
 sg13g2_decap_8 FILLER_78_798 ();
 sg13g2_decap_8 FILLER_78_805 ();
 sg13g2_decap_8 FILLER_78_812 ();
 sg13g2_decap_8 FILLER_78_819 ();
 sg13g2_decap_8 FILLER_78_826 ();
 sg13g2_decap_8 FILLER_78_833 ();
 sg13g2_fill_1 FILLER_78_840 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_decap_8 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_77 ();
 sg13g2_decap_8 FILLER_79_84 ();
 sg13g2_decap_8 FILLER_79_91 ();
 sg13g2_decap_8 FILLER_79_98 ();
 sg13g2_decap_8 FILLER_79_105 ();
 sg13g2_decap_8 FILLER_79_112 ();
 sg13g2_decap_8 FILLER_79_119 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_8 FILLER_79_154 ();
 sg13g2_decap_8 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_168 ();
 sg13g2_decap_8 FILLER_79_175 ();
 sg13g2_decap_8 FILLER_79_182 ();
 sg13g2_decap_8 FILLER_79_189 ();
 sg13g2_decap_8 FILLER_79_196 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_decap_8 FILLER_79_210 ();
 sg13g2_decap_8 FILLER_79_217 ();
 sg13g2_decap_8 FILLER_79_224 ();
 sg13g2_decap_8 FILLER_79_231 ();
 sg13g2_decap_8 FILLER_79_238 ();
 sg13g2_decap_8 FILLER_79_245 ();
 sg13g2_decap_8 FILLER_79_252 ();
 sg13g2_decap_8 FILLER_79_259 ();
 sg13g2_decap_8 FILLER_79_266 ();
 sg13g2_decap_8 FILLER_79_273 ();
 sg13g2_decap_8 FILLER_79_280 ();
 sg13g2_decap_8 FILLER_79_287 ();
 sg13g2_decap_8 FILLER_79_294 ();
 sg13g2_decap_8 FILLER_79_301 ();
 sg13g2_decap_8 FILLER_79_308 ();
 sg13g2_decap_8 FILLER_79_315 ();
 sg13g2_decap_8 FILLER_79_322 ();
 sg13g2_decap_8 FILLER_79_329 ();
 sg13g2_decap_8 FILLER_79_336 ();
 sg13g2_decap_8 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_350 ();
 sg13g2_decap_8 FILLER_79_357 ();
 sg13g2_decap_8 FILLER_79_364 ();
 sg13g2_decap_8 FILLER_79_371 ();
 sg13g2_decap_8 FILLER_79_378 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_decap_8 FILLER_79_406 ();
 sg13g2_decap_8 FILLER_79_413 ();
 sg13g2_decap_8 FILLER_79_420 ();
 sg13g2_decap_8 FILLER_79_427 ();
 sg13g2_decap_8 FILLER_79_434 ();
 sg13g2_decap_8 FILLER_79_441 ();
 sg13g2_decap_8 FILLER_79_448 ();
 sg13g2_decap_8 FILLER_79_455 ();
 sg13g2_decap_8 FILLER_79_462 ();
 sg13g2_decap_8 FILLER_79_469 ();
 sg13g2_decap_8 FILLER_79_476 ();
 sg13g2_decap_8 FILLER_79_483 ();
 sg13g2_decap_8 FILLER_79_490 ();
 sg13g2_decap_8 FILLER_79_497 ();
 sg13g2_decap_8 FILLER_79_504 ();
 sg13g2_decap_8 FILLER_79_511 ();
 sg13g2_decap_8 FILLER_79_518 ();
 sg13g2_decap_8 FILLER_79_525 ();
 sg13g2_decap_8 FILLER_79_532 ();
 sg13g2_decap_8 FILLER_79_539 ();
 sg13g2_decap_8 FILLER_79_546 ();
 sg13g2_decap_8 FILLER_79_553 ();
 sg13g2_decap_8 FILLER_79_560 ();
 sg13g2_decap_8 FILLER_79_567 ();
 sg13g2_decap_8 FILLER_79_574 ();
 sg13g2_decap_8 FILLER_79_581 ();
 sg13g2_decap_8 FILLER_79_588 ();
 sg13g2_decap_8 FILLER_79_595 ();
 sg13g2_decap_8 FILLER_79_602 ();
 sg13g2_decap_8 FILLER_79_609 ();
 sg13g2_decap_8 FILLER_79_616 ();
 sg13g2_decap_8 FILLER_79_623 ();
 sg13g2_decap_8 FILLER_79_630 ();
 sg13g2_decap_8 FILLER_79_637 ();
 sg13g2_decap_8 FILLER_79_644 ();
 sg13g2_decap_8 FILLER_79_651 ();
 sg13g2_decap_8 FILLER_79_658 ();
 sg13g2_decap_8 FILLER_79_665 ();
 sg13g2_decap_8 FILLER_79_672 ();
 sg13g2_decap_8 FILLER_79_679 ();
 sg13g2_decap_8 FILLER_79_686 ();
 sg13g2_decap_8 FILLER_79_693 ();
 sg13g2_decap_8 FILLER_79_700 ();
 sg13g2_decap_8 FILLER_79_707 ();
 sg13g2_decap_8 FILLER_79_714 ();
 sg13g2_decap_8 FILLER_79_721 ();
 sg13g2_decap_8 FILLER_79_728 ();
 sg13g2_decap_8 FILLER_79_735 ();
 sg13g2_decap_8 FILLER_79_742 ();
 sg13g2_decap_8 FILLER_79_749 ();
 sg13g2_decap_8 FILLER_79_756 ();
 sg13g2_decap_8 FILLER_79_763 ();
 sg13g2_decap_8 FILLER_79_770 ();
 sg13g2_decap_8 FILLER_79_777 ();
 sg13g2_decap_8 FILLER_79_784 ();
 sg13g2_decap_8 FILLER_79_791 ();
 sg13g2_decap_8 FILLER_79_798 ();
 sg13g2_decap_8 FILLER_79_805 ();
 sg13g2_decap_8 FILLER_79_812 ();
 sg13g2_decap_8 FILLER_79_819 ();
 sg13g2_decap_8 FILLER_79_826 ();
 sg13g2_decap_8 FILLER_79_833 ();
 sg13g2_fill_1 FILLER_79_840 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_77 ();
 sg13g2_decap_8 FILLER_80_84 ();
 sg13g2_decap_8 FILLER_80_91 ();
 sg13g2_decap_8 FILLER_80_98 ();
 sg13g2_decap_8 FILLER_80_105 ();
 sg13g2_decap_8 FILLER_80_112 ();
 sg13g2_decap_8 FILLER_80_119 ();
 sg13g2_decap_8 FILLER_80_126 ();
 sg13g2_decap_8 FILLER_80_133 ();
 sg13g2_decap_8 FILLER_80_140 ();
 sg13g2_decap_8 FILLER_80_147 ();
 sg13g2_decap_8 FILLER_80_154 ();
 sg13g2_decap_8 FILLER_80_161 ();
 sg13g2_decap_8 FILLER_80_168 ();
 sg13g2_decap_8 FILLER_80_175 ();
 sg13g2_decap_8 FILLER_80_182 ();
 sg13g2_decap_8 FILLER_80_189 ();
 sg13g2_decap_8 FILLER_80_196 ();
 sg13g2_decap_8 FILLER_80_203 ();
 sg13g2_decap_8 FILLER_80_210 ();
 sg13g2_decap_8 FILLER_80_217 ();
 sg13g2_decap_8 FILLER_80_224 ();
 sg13g2_decap_8 FILLER_80_231 ();
 sg13g2_decap_8 FILLER_80_238 ();
 sg13g2_decap_8 FILLER_80_245 ();
 sg13g2_decap_8 FILLER_80_252 ();
 sg13g2_decap_8 FILLER_80_259 ();
 sg13g2_decap_8 FILLER_80_266 ();
 sg13g2_decap_8 FILLER_80_273 ();
 sg13g2_decap_8 FILLER_80_280 ();
 sg13g2_decap_8 FILLER_80_287 ();
 sg13g2_decap_8 FILLER_80_294 ();
 sg13g2_decap_8 FILLER_80_301 ();
 sg13g2_decap_8 FILLER_80_308 ();
 sg13g2_decap_8 FILLER_80_315 ();
 sg13g2_decap_8 FILLER_80_322 ();
 sg13g2_decap_8 FILLER_80_329 ();
 sg13g2_decap_8 FILLER_80_336 ();
 sg13g2_decap_8 FILLER_80_343 ();
 sg13g2_decap_8 FILLER_80_350 ();
 sg13g2_decap_8 FILLER_80_357 ();
 sg13g2_decap_8 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_371 ();
 sg13g2_decap_8 FILLER_80_378 ();
 sg13g2_decap_8 FILLER_80_385 ();
 sg13g2_decap_8 FILLER_80_392 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_decap_8 FILLER_80_406 ();
 sg13g2_decap_8 FILLER_80_413 ();
 sg13g2_decap_8 FILLER_80_420 ();
 sg13g2_decap_8 FILLER_80_427 ();
 sg13g2_decap_8 FILLER_80_434 ();
 sg13g2_decap_8 FILLER_80_441 ();
 sg13g2_decap_8 FILLER_80_448 ();
 sg13g2_decap_8 FILLER_80_455 ();
 sg13g2_decap_8 FILLER_80_462 ();
 sg13g2_decap_8 FILLER_80_469 ();
 sg13g2_decap_8 FILLER_80_476 ();
 sg13g2_decap_8 FILLER_80_483 ();
 sg13g2_decap_8 FILLER_80_490 ();
 sg13g2_decap_8 FILLER_80_497 ();
 sg13g2_decap_8 FILLER_80_504 ();
 sg13g2_decap_8 FILLER_80_511 ();
 sg13g2_decap_8 FILLER_80_518 ();
 sg13g2_decap_8 FILLER_80_525 ();
 sg13g2_decap_8 FILLER_80_532 ();
 sg13g2_decap_8 FILLER_80_539 ();
 sg13g2_decap_8 FILLER_80_546 ();
 sg13g2_decap_8 FILLER_80_553 ();
 sg13g2_decap_8 FILLER_80_560 ();
 sg13g2_decap_8 FILLER_80_567 ();
 sg13g2_decap_8 FILLER_80_574 ();
 sg13g2_decap_8 FILLER_80_581 ();
 sg13g2_decap_8 FILLER_80_588 ();
 sg13g2_decap_8 FILLER_80_595 ();
 sg13g2_decap_8 FILLER_80_602 ();
 sg13g2_decap_8 FILLER_80_609 ();
 sg13g2_decap_8 FILLER_80_616 ();
 sg13g2_decap_8 FILLER_80_623 ();
 sg13g2_decap_8 FILLER_80_630 ();
 sg13g2_decap_8 FILLER_80_637 ();
 sg13g2_decap_8 FILLER_80_644 ();
 sg13g2_decap_8 FILLER_80_651 ();
 sg13g2_decap_8 FILLER_80_658 ();
 sg13g2_decap_8 FILLER_80_665 ();
 sg13g2_decap_8 FILLER_80_672 ();
 sg13g2_decap_8 FILLER_80_679 ();
 sg13g2_decap_8 FILLER_80_686 ();
 sg13g2_decap_8 FILLER_80_693 ();
 sg13g2_decap_8 FILLER_80_700 ();
 sg13g2_decap_8 FILLER_80_707 ();
 sg13g2_decap_8 FILLER_80_714 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_728 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_decap_8 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_decap_8 FILLER_80_770 ();
 sg13g2_decap_8 FILLER_80_777 ();
 sg13g2_decap_8 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_791 ();
 sg13g2_decap_8 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_805 ();
 sg13g2_decap_8 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_8 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_833 ();
 sg13g2_fill_1 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_81_0 ();
 sg13g2_decap_8 FILLER_81_7 ();
 sg13g2_decap_8 FILLER_81_14 ();
 sg13g2_decap_8 FILLER_81_21 ();
 sg13g2_decap_8 FILLER_81_28 ();
 sg13g2_decap_8 FILLER_81_35 ();
 sg13g2_decap_8 FILLER_81_42 ();
 sg13g2_decap_8 FILLER_81_49 ();
 sg13g2_decap_8 FILLER_81_56 ();
 sg13g2_decap_8 FILLER_81_63 ();
 sg13g2_decap_8 FILLER_81_70 ();
 sg13g2_decap_8 FILLER_81_77 ();
 sg13g2_decap_8 FILLER_81_84 ();
 sg13g2_decap_8 FILLER_81_91 ();
 sg13g2_decap_8 FILLER_81_98 ();
 sg13g2_decap_8 FILLER_81_105 ();
 sg13g2_decap_8 FILLER_81_112 ();
 sg13g2_decap_8 FILLER_81_119 ();
 sg13g2_decap_8 FILLER_81_126 ();
 sg13g2_decap_8 FILLER_81_133 ();
 sg13g2_decap_8 FILLER_81_140 ();
 sg13g2_decap_8 FILLER_81_147 ();
 sg13g2_decap_8 FILLER_81_154 ();
 sg13g2_decap_8 FILLER_81_161 ();
 sg13g2_decap_8 FILLER_81_168 ();
 sg13g2_decap_8 FILLER_81_175 ();
 sg13g2_decap_8 FILLER_81_182 ();
 sg13g2_decap_8 FILLER_81_189 ();
 sg13g2_decap_8 FILLER_81_196 ();
 sg13g2_decap_8 FILLER_81_203 ();
 sg13g2_decap_8 FILLER_81_210 ();
 sg13g2_decap_8 FILLER_81_217 ();
 sg13g2_decap_8 FILLER_81_224 ();
 sg13g2_decap_8 FILLER_81_231 ();
 sg13g2_decap_8 FILLER_81_238 ();
 sg13g2_decap_8 FILLER_81_245 ();
 sg13g2_decap_8 FILLER_81_252 ();
 sg13g2_decap_8 FILLER_81_259 ();
 sg13g2_decap_8 FILLER_81_266 ();
 sg13g2_decap_8 FILLER_81_273 ();
 sg13g2_decap_8 FILLER_81_280 ();
 sg13g2_decap_8 FILLER_81_287 ();
 sg13g2_decap_8 FILLER_81_294 ();
 sg13g2_decap_8 FILLER_81_301 ();
 sg13g2_decap_8 FILLER_81_308 ();
 sg13g2_decap_8 FILLER_81_315 ();
 sg13g2_decap_8 FILLER_81_322 ();
 sg13g2_decap_8 FILLER_81_329 ();
 sg13g2_decap_8 FILLER_81_336 ();
 sg13g2_decap_8 FILLER_81_343 ();
 sg13g2_decap_8 FILLER_81_350 ();
 sg13g2_decap_8 FILLER_81_357 ();
 sg13g2_decap_8 FILLER_81_364 ();
 sg13g2_decap_8 FILLER_81_371 ();
 sg13g2_decap_8 FILLER_81_378 ();
 sg13g2_decap_8 FILLER_81_385 ();
 sg13g2_decap_8 FILLER_81_392 ();
 sg13g2_decap_8 FILLER_81_399 ();
 sg13g2_decap_8 FILLER_81_406 ();
 sg13g2_decap_8 FILLER_81_413 ();
 sg13g2_decap_8 FILLER_81_420 ();
 sg13g2_decap_8 FILLER_81_427 ();
 sg13g2_decap_8 FILLER_81_434 ();
 sg13g2_decap_8 FILLER_81_441 ();
 sg13g2_decap_8 FILLER_81_448 ();
 sg13g2_decap_8 FILLER_81_455 ();
 sg13g2_decap_8 FILLER_81_462 ();
 sg13g2_decap_8 FILLER_81_469 ();
 sg13g2_decap_8 FILLER_81_476 ();
 sg13g2_decap_8 FILLER_81_483 ();
 sg13g2_decap_8 FILLER_81_490 ();
 sg13g2_decap_8 FILLER_81_497 ();
 sg13g2_decap_8 FILLER_81_504 ();
 sg13g2_decap_8 FILLER_81_511 ();
 sg13g2_decap_8 FILLER_81_518 ();
 sg13g2_decap_8 FILLER_81_525 ();
 sg13g2_decap_8 FILLER_81_532 ();
 sg13g2_decap_8 FILLER_81_539 ();
 sg13g2_decap_8 FILLER_81_546 ();
 sg13g2_decap_8 FILLER_81_553 ();
 sg13g2_decap_8 FILLER_81_560 ();
 sg13g2_decap_8 FILLER_81_567 ();
 sg13g2_decap_8 FILLER_81_574 ();
 sg13g2_decap_8 FILLER_81_581 ();
 sg13g2_decap_8 FILLER_81_588 ();
 sg13g2_decap_8 FILLER_81_595 ();
 sg13g2_decap_8 FILLER_81_602 ();
 sg13g2_decap_8 FILLER_81_609 ();
 sg13g2_decap_8 FILLER_81_616 ();
 sg13g2_decap_8 FILLER_81_623 ();
 sg13g2_decap_8 FILLER_81_630 ();
 sg13g2_decap_8 FILLER_81_637 ();
 sg13g2_decap_8 FILLER_81_644 ();
 sg13g2_decap_8 FILLER_81_651 ();
 sg13g2_decap_8 FILLER_81_658 ();
 sg13g2_decap_8 FILLER_81_665 ();
 sg13g2_decap_8 FILLER_81_672 ();
 sg13g2_decap_8 FILLER_81_679 ();
 sg13g2_decap_8 FILLER_81_686 ();
 sg13g2_decap_8 FILLER_81_693 ();
 sg13g2_decap_8 FILLER_81_700 ();
 sg13g2_decap_8 FILLER_81_707 ();
 sg13g2_decap_8 FILLER_81_714 ();
 sg13g2_decap_8 FILLER_81_721 ();
 sg13g2_decap_8 FILLER_81_728 ();
 sg13g2_decap_8 FILLER_81_735 ();
 sg13g2_decap_8 FILLER_81_742 ();
 sg13g2_decap_8 FILLER_81_749 ();
 sg13g2_decap_8 FILLER_81_756 ();
 sg13g2_decap_8 FILLER_81_763 ();
 sg13g2_decap_8 FILLER_81_770 ();
 sg13g2_decap_8 FILLER_81_777 ();
 sg13g2_decap_8 FILLER_81_784 ();
 sg13g2_decap_8 FILLER_81_791 ();
 sg13g2_decap_8 FILLER_81_798 ();
 sg13g2_decap_8 FILLER_81_805 ();
 sg13g2_decap_8 FILLER_81_812 ();
 sg13g2_decap_8 FILLER_81_819 ();
 sg13g2_decap_8 FILLER_81_826 ();
 sg13g2_decap_8 FILLER_81_833 ();
 sg13g2_fill_1 FILLER_81_840 ();
 sg13g2_decap_8 FILLER_82_0 ();
 sg13g2_decap_8 FILLER_82_7 ();
 sg13g2_decap_8 FILLER_82_14 ();
 sg13g2_decap_8 FILLER_82_21 ();
 sg13g2_decap_8 FILLER_82_28 ();
 sg13g2_decap_8 FILLER_82_35 ();
 sg13g2_decap_8 FILLER_82_42 ();
 sg13g2_decap_8 FILLER_82_49 ();
 sg13g2_decap_8 FILLER_82_56 ();
 sg13g2_decap_8 FILLER_82_63 ();
 sg13g2_decap_8 FILLER_82_70 ();
 sg13g2_decap_8 FILLER_82_77 ();
 sg13g2_decap_8 FILLER_82_84 ();
 sg13g2_decap_8 FILLER_82_91 ();
 sg13g2_decap_8 FILLER_82_98 ();
 sg13g2_decap_8 FILLER_82_105 ();
 sg13g2_decap_8 FILLER_82_112 ();
 sg13g2_decap_8 FILLER_82_119 ();
 sg13g2_decap_8 FILLER_82_126 ();
 sg13g2_decap_8 FILLER_82_133 ();
 sg13g2_decap_8 FILLER_82_140 ();
 sg13g2_decap_8 FILLER_82_147 ();
 sg13g2_decap_8 FILLER_82_154 ();
 sg13g2_decap_8 FILLER_82_161 ();
 sg13g2_decap_8 FILLER_82_168 ();
 sg13g2_decap_8 FILLER_82_175 ();
 sg13g2_decap_8 FILLER_82_182 ();
 sg13g2_decap_8 FILLER_82_189 ();
 sg13g2_decap_8 FILLER_82_196 ();
 sg13g2_decap_8 FILLER_82_203 ();
 sg13g2_decap_8 FILLER_82_210 ();
 sg13g2_decap_8 FILLER_82_217 ();
 sg13g2_decap_8 FILLER_82_224 ();
 sg13g2_decap_8 FILLER_82_231 ();
 sg13g2_decap_8 FILLER_82_238 ();
 sg13g2_decap_8 FILLER_82_245 ();
 sg13g2_decap_8 FILLER_82_252 ();
 sg13g2_decap_8 FILLER_82_259 ();
 sg13g2_decap_8 FILLER_82_266 ();
 sg13g2_decap_8 FILLER_82_273 ();
 sg13g2_decap_8 FILLER_82_280 ();
 sg13g2_decap_8 FILLER_82_287 ();
 sg13g2_decap_8 FILLER_82_294 ();
 sg13g2_decap_8 FILLER_82_301 ();
 sg13g2_decap_8 FILLER_82_308 ();
 sg13g2_decap_8 FILLER_82_315 ();
 sg13g2_decap_8 FILLER_82_322 ();
 sg13g2_decap_8 FILLER_82_329 ();
 sg13g2_decap_8 FILLER_82_336 ();
 sg13g2_decap_8 FILLER_82_343 ();
 sg13g2_decap_8 FILLER_82_350 ();
 sg13g2_decap_8 FILLER_82_357 ();
 sg13g2_decap_8 FILLER_82_364 ();
 sg13g2_decap_8 FILLER_82_371 ();
 sg13g2_decap_8 FILLER_82_378 ();
 sg13g2_decap_8 FILLER_82_385 ();
 sg13g2_decap_8 FILLER_82_392 ();
 sg13g2_decap_8 FILLER_82_399 ();
 sg13g2_decap_8 FILLER_82_406 ();
 sg13g2_decap_8 FILLER_82_413 ();
 sg13g2_decap_8 FILLER_82_420 ();
 sg13g2_decap_8 FILLER_82_427 ();
 sg13g2_decap_8 FILLER_82_434 ();
 sg13g2_decap_8 FILLER_82_441 ();
 sg13g2_decap_8 FILLER_82_448 ();
 sg13g2_decap_8 FILLER_82_455 ();
 sg13g2_decap_8 FILLER_82_462 ();
 sg13g2_decap_8 FILLER_82_469 ();
 sg13g2_decap_8 FILLER_82_476 ();
 sg13g2_decap_8 FILLER_82_483 ();
 sg13g2_decap_8 FILLER_82_490 ();
 sg13g2_decap_8 FILLER_82_497 ();
 sg13g2_decap_8 FILLER_82_504 ();
 sg13g2_decap_8 FILLER_82_511 ();
 sg13g2_decap_8 FILLER_82_518 ();
 sg13g2_decap_8 FILLER_82_525 ();
 sg13g2_decap_8 FILLER_82_532 ();
 sg13g2_decap_8 FILLER_82_539 ();
 sg13g2_decap_8 FILLER_82_546 ();
 sg13g2_decap_8 FILLER_82_553 ();
 sg13g2_decap_8 FILLER_82_560 ();
 sg13g2_decap_8 FILLER_82_567 ();
 sg13g2_decap_8 FILLER_82_574 ();
 sg13g2_decap_8 FILLER_82_581 ();
 sg13g2_decap_8 FILLER_82_588 ();
 sg13g2_decap_8 FILLER_82_595 ();
 sg13g2_decap_8 FILLER_82_602 ();
 sg13g2_decap_8 FILLER_82_609 ();
 sg13g2_decap_8 FILLER_82_616 ();
 sg13g2_decap_8 FILLER_82_623 ();
 sg13g2_decap_8 FILLER_82_630 ();
 sg13g2_decap_8 FILLER_82_637 ();
 sg13g2_decap_8 FILLER_82_644 ();
 sg13g2_decap_8 FILLER_82_651 ();
 sg13g2_decap_8 FILLER_82_658 ();
 sg13g2_decap_8 FILLER_82_665 ();
 sg13g2_decap_8 FILLER_82_672 ();
 sg13g2_decap_8 FILLER_82_679 ();
 sg13g2_decap_8 FILLER_82_686 ();
 sg13g2_decap_8 FILLER_82_693 ();
 sg13g2_decap_8 FILLER_82_700 ();
 sg13g2_decap_8 FILLER_82_707 ();
 sg13g2_decap_8 FILLER_82_714 ();
 sg13g2_decap_8 FILLER_82_721 ();
 sg13g2_decap_8 FILLER_82_728 ();
 sg13g2_decap_8 FILLER_82_735 ();
 sg13g2_decap_8 FILLER_82_742 ();
 sg13g2_decap_8 FILLER_82_749 ();
 sg13g2_decap_8 FILLER_82_756 ();
 sg13g2_decap_8 FILLER_82_763 ();
 sg13g2_decap_8 FILLER_82_770 ();
 sg13g2_decap_8 FILLER_82_777 ();
 sg13g2_decap_8 FILLER_82_784 ();
 sg13g2_decap_8 FILLER_82_791 ();
 sg13g2_decap_8 FILLER_82_798 ();
 sg13g2_decap_8 FILLER_82_805 ();
 sg13g2_decap_8 FILLER_82_812 ();
 sg13g2_decap_8 FILLER_82_819 ();
 sg13g2_decap_8 FILLER_82_826 ();
 sg13g2_decap_8 FILLER_82_833 ();
 sg13g2_fill_1 FILLER_82_840 ();
 sg13g2_decap_8 FILLER_83_0 ();
 sg13g2_decap_8 FILLER_83_7 ();
 sg13g2_decap_8 FILLER_83_14 ();
 sg13g2_decap_8 FILLER_83_21 ();
 sg13g2_decap_8 FILLER_83_28 ();
 sg13g2_decap_8 FILLER_83_35 ();
 sg13g2_decap_8 FILLER_83_42 ();
 sg13g2_decap_8 FILLER_83_49 ();
 sg13g2_decap_8 FILLER_83_56 ();
 sg13g2_decap_8 FILLER_83_63 ();
 sg13g2_decap_8 FILLER_83_70 ();
 sg13g2_decap_8 FILLER_83_77 ();
 sg13g2_decap_8 FILLER_83_84 ();
 sg13g2_decap_8 FILLER_83_91 ();
 sg13g2_decap_8 FILLER_83_98 ();
 sg13g2_decap_8 FILLER_83_105 ();
 sg13g2_decap_8 FILLER_83_112 ();
 sg13g2_decap_8 FILLER_83_119 ();
 sg13g2_decap_8 FILLER_83_126 ();
 sg13g2_decap_8 FILLER_83_133 ();
 sg13g2_decap_8 FILLER_83_140 ();
 sg13g2_decap_8 FILLER_83_147 ();
 sg13g2_decap_8 FILLER_83_154 ();
 sg13g2_decap_8 FILLER_83_161 ();
 sg13g2_decap_8 FILLER_83_168 ();
 sg13g2_decap_8 FILLER_83_175 ();
 sg13g2_decap_8 FILLER_83_182 ();
 sg13g2_decap_8 FILLER_83_189 ();
 sg13g2_decap_8 FILLER_83_196 ();
 sg13g2_decap_8 FILLER_83_203 ();
 sg13g2_decap_8 FILLER_83_210 ();
 sg13g2_decap_8 FILLER_83_217 ();
 sg13g2_decap_8 FILLER_83_224 ();
 sg13g2_decap_8 FILLER_83_231 ();
 sg13g2_decap_8 FILLER_83_238 ();
 sg13g2_decap_8 FILLER_83_245 ();
 sg13g2_decap_8 FILLER_83_252 ();
 sg13g2_decap_8 FILLER_83_259 ();
 sg13g2_decap_8 FILLER_83_266 ();
 sg13g2_decap_8 FILLER_83_273 ();
 sg13g2_decap_8 FILLER_83_280 ();
 sg13g2_decap_8 FILLER_83_287 ();
 sg13g2_decap_8 FILLER_83_294 ();
 sg13g2_decap_8 FILLER_83_301 ();
 sg13g2_decap_8 FILLER_83_308 ();
 sg13g2_decap_8 FILLER_83_315 ();
 sg13g2_decap_8 FILLER_83_322 ();
 sg13g2_decap_8 FILLER_83_329 ();
 sg13g2_decap_8 FILLER_83_336 ();
 sg13g2_decap_8 FILLER_83_343 ();
 sg13g2_decap_8 FILLER_83_350 ();
 sg13g2_decap_8 FILLER_83_357 ();
 sg13g2_decap_8 FILLER_83_364 ();
 sg13g2_decap_8 FILLER_83_371 ();
 sg13g2_decap_8 FILLER_83_378 ();
 sg13g2_decap_8 FILLER_83_385 ();
 sg13g2_decap_8 FILLER_83_392 ();
 sg13g2_decap_8 FILLER_83_399 ();
 sg13g2_decap_8 FILLER_83_406 ();
 sg13g2_decap_8 FILLER_83_413 ();
 sg13g2_decap_8 FILLER_83_420 ();
 sg13g2_decap_8 FILLER_83_427 ();
 sg13g2_decap_8 FILLER_83_434 ();
 sg13g2_decap_8 FILLER_83_441 ();
 sg13g2_decap_8 FILLER_83_448 ();
 sg13g2_decap_8 FILLER_83_455 ();
 sg13g2_decap_8 FILLER_83_462 ();
 sg13g2_decap_8 FILLER_83_469 ();
 sg13g2_decap_8 FILLER_83_476 ();
 sg13g2_decap_8 FILLER_83_483 ();
 sg13g2_decap_8 FILLER_83_490 ();
 sg13g2_decap_8 FILLER_83_497 ();
 sg13g2_decap_8 FILLER_83_504 ();
 sg13g2_decap_8 FILLER_83_511 ();
 sg13g2_decap_8 FILLER_83_518 ();
 sg13g2_decap_8 FILLER_83_525 ();
 sg13g2_decap_8 FILLER_83_532 ();
 sg13g2_decap_8 FILLER_83_539 ();
 sg13g2_decap_8 FILLER_83_546 ();
 sg13g2_decap_8 FILLER_83_553 ();
 sg13g2_decap_8 FILLER_83_560 ();
 sg13g2_decap_8 FILLER_83_567 ();
 sg13g2_decap_8 FILLER_83_574 ();
 sg13g2_decap_8 FILLER_83_581 ();
 sg13g2_decap_8 FILLER_83_588 ();
 sg13g2_decap_8 FILLER_83_595 ();
 sg13g2_decap_8 FILLER_83_602 ();
 sg13g2_decap_8 FILLER_83_609 ();
 sg13g2_decap_8 FILLER_83_616 ();
 sg13g2_decap_8 FILLER_83_623 ();
 sg13g2_decap_8 FILLER_83_630 ();
 sg13g2_decap_8 FILLER_83_637 ();
 sg13g2_decap_8 FILLER_83_644 ();
 sg13g2_decap_8 FILLER_83_651 ();
 sg13g2_decap_8 FILLER_83_658 ();
 sg13g2_decap_8 FILLER_83_665 ();
 sg13g2_decap_8 FILLER_83_672 ();
 sg13g2_decap_8 FILLER_83_679 ();
 sg13g2_decap_8 FILLER_83_686 ();
 sg13g2_decap_8 FILLER_83_693 ();
 sg13g2_decap_8 FILLER_83_700 ();
 sg13g2_decap_8 FILLER_83_707 ();
 sg13g2_decap_8 FILLER_83_714 ();
 sg13g2_decap_8 FILLER_83_721 ();
 sg13g2_decap_8 FILLER_83_728 ();
 sg13g2_decap_8 FILLER_83_735 ();
 sg13g2_decap_8 FILLER_83_742 ();
 sg13g2_decap_8 FILLER_83_749 ();
 sg13g2_decap_8 FILLER_83_756 ();
 sg13g2_decap_8 FILLER_83_763 ();
 sg13g2_decap_8 FILLER_83_770 ();
 sg13g2_decap_8 FILLER_83_777 ();
 sg13g2_decap_8 FILLER_83_784 ();
 sg13g2_decap_8 FILLER_83_791 ();
 sg13g2_decap_8 FILLER_83_798 ();
 sg13g2_decap_8 FILLER_83_805 ();
 sg13g2_decap_8 FILLER_83_812 ();
 sg13g2_decap_8 FILLER_83_819 ();
 sg13g2_decap_8 FILLER_83_826 ();
 sg13g2_decap_8 FILLER_83_833 ();
 sg13g2_fill_1 FILLER_83_840 ();
 sg13g2_decap_8 FILLER_84_0 ();
 sg13g2_decap_8 FILLER_84_7 ();
 sg13g2_decap_8 FILLER_84_14 ();
 sg13g2_decap_8 FILLER_84_21 ();
 sg13g2_decap_8 FILLER_84_28 ();
 sg13g2_decap_8 FILLER_84_35 ();
 sg13g2_decap_8 FILLER_84_42 ();
 sg13g2_decap_8 FILLER_84_49 ();
 sg13g2_decap_8 FILLER_84_56 ();
 sg13g2_decap_8 FILLER_84_63 ();
 sg13g2_decap_8 FILLER_84_70 ();
 sg13g2_decap_8 FILLER_84_77 ();
 sg13g2_decap_8 FILLER_84_84 ();
 sg13g2_decap_8 FILLER_84_91 ();
 sg13g2_decap_8 FILLER_84_98 ();
 sg13g2_decap_8 FILLER_84_105 ();
 sg13g2_decap_8 FILLER_84_112 ();
 sg13g2_decap_8 FILLER_84_119 ();
 sg13g2_decap_8 FILLER_84_126 ();
 sg13g2_decap_8 FILLER_84_133 ();
 sg13g2_decap_8 FILLER_84_140 ();
 sg13g2_decap_8 FILLER_84_147 ();
 sg13g2_decap_8 FILLER_84_154 ();
 sg13g2_decap_8 FILLER_84_161 ();
 sg13g2_decap_8 FILLER_84_168 ();
 sg13g2_decap_8 FILLER_84_175 ();
 sg13g2_decap_8 FILLER_84_182 ();
 sg13g2_decap_8 FILLER_84_189 ();
 sg13g2_decap_8 FILLER_84_196 ();
 sg13g2_decap_8 FILLER_84_203 ();
 sg13g2_decap_8 FILLER_84_210 ();
 sg13g2_decap_8 FILLER_84_217 ();
 sg13g2_decap_8 FILLER_84_224 ();
 sg13g2_decap_8 FILLER_84_231 ();
 sg13g2_decap_8 FILLER_84_238 ();
 sg13g2_decap_8 FILLER_84_245 ();
 sg13g2_decap_8 FILLER_84_252 ();
 sg13g2_decap_8 FILLER_84_259 ();
 sg13g2_decap_8 FILLER_84_266 ();
 sg13g2_decap_8 FILLER_84_273 ();
 sg13g2_decap_8 FILLER_84_280 ();
 sg13g2_decap_8 FILLER_84_287 ();
 sg13g2_decap_8 FILLER_84_294 ();
 sg13g2_decap_8 FILLER_84_301 ();
 sg13g2_decap_8 FILLER_84_308 ();
 sg13g2_decap_8 FILLER_84_315 ();
 sg13g2_decap_8 FILLER_84_322 ();
 sg13g2_decap_8 FILLER_84_329 ();
 sg13g2_decap_8 FILLER_84_336 ();
 sg13g2_decap_8 FILLER_84_343 ();
 sg13g2_decap_8 FILLER_84_350 ();
 sg13g2_decap_8 FILLER_84_357 ();
 sg13g2_decap_8 FILLER_84_364 ();
 sg13g2_decap_8 FILLER_84_371 ();
 sg13g2_decap_8 FILLER_84_378 ();
 sg13g2_decap_8 FILLER_84_385 ();
 sg13g2_decap_8 FILLER_84_392 ();
 sg13g2_decap_8 FILLER_84_399 ();
 sg13g2_decap_8 FILLER_84_406 ();
 sg13g2_decap_8 FILLER_84_413 ();
 sg13g2_decap_8 FILLER_84_420 ();
 sg13g2_decap_8 FILLER_84_427 ();
 sg13g2_decap_8 FILLER_84_434 ();
 sg13g2_decap_8 FILLER_84_441 ();
 sg13g2_decap_8 FILLER_84_448 ();
 sg13g2_decap_8 FILLER_84_455 ();
 sg13g2_decap_8 FILLER_84_462 ();
 sg13g2_decap_8 FILLER_84_469 ();
 sg13g2_decap_8 FILLER_84_476 ();
 sg13g2_decap_8 FILLER_84_483 ();
 sg13g2_decap_8 FILLER_84_490 ();
 sg13g2_decap_8 FILLER_84_497 ();
 sg13g2_decap_8 FILLER_84_504 ();
 sg13g2_decap_8 FILLER_84_511 ();
 sg13g2_decap_8 FILLER_84_518 ();
 sg13g2_decap_8 FILLER_84_525 ();
 sg13g2_decap_8 FILLER_84_532 ();
 sg13g2_decap_8 FILLER_84_539 ();
 sg13g2_decap_8 FILLER_84_546 ();
 sg13g2_decap_8 FILLER_84_553 ();
 sg13g2_decap_8 FILLER_84_560 ();
 sg13g2_decap_8 FILLER_84_567 ();
 sg13g2_decap_8 FILLER_84_574 ();
 sg13g2_decap_8 FILLER_84_581 ();
 sg13g2_decap_8 FILLER_84_588 ();
 sg13g2_decap_8 FILLER_84_595 ();
 sg13g2_decap_8 FILLER_84_602 ();
 sg13g2_decap_8 FILLER_84_609 ();
 sg13g2_decap_8 FILLER_84_616 ();
 sg13g2_decap_8 FILLER_84_623 ();
 sg13g2_decap_8 FILLER_84_630 ();
 sg13g2_decap_8 FILLER_84_637 ();
 sg13g2_decap_8 FILLER_84_644 ();
 sg13g2_decap_8 FILLER_84_651 ();
 sg13g2_decap_8 FILLER_84_658 ();
 sg13g2_decap_8 FILLER_84_665 ();
 sg13g2_decap_8 FILLER_84_672 ();
 sg13g2_decap_8 FILLER_84_679 ();
 sg13g2_decap_8 FILLER_84_686 ();
 sg13g2_decap_8 FILLER_84_693 ();
 sg13g2_decap_8 FILLER_84_700 ();
 sg13g2_decap_8 FILLER_84_707 ();
 sg13g2_decap_8 FILLER_84_714 ();
 sg13g2_decap_8 FILLER_84_721 ();
 sg13g2_decap_8 FILLER_84_728 ();
 sg13g2_decap_8 FILLER_84_735 ();
 sg13g2_decap_8 FILLER_84_742 ();
 sg13g2_decap_8 FILLER_84_749 ();
 sg13g2_decap_8 FILLER_84_756 ();
 sg13g2_decap_8 FILLER_84_763 ();
 sg13g2_decap_8 FILLER_84_770 ();
 sg13g2_decap_8 FILLER_84_777 ();
 sg13g2_decap_8 FILLER_84_784 ();
 sg13g2_decap_8 FILLER_84_791 ();
 sg13g2_decap_8 FILLER_84_798 ();
 sg13g2_decap_8 FILLER_84_805 ();
 sg13g2_decap_8 FILLER_84_812 ();
 sg13g2_decap_8 FILLER_84_819 ();
 sg13g2_decap_8 FILLER_84_826 ();
 sg13g2_decap_8 FILLER_84_833 ();
 sg13g2_fill_1 FILLER_84_840 ();
 sg13g2_decap_8 FILLER_85_0 ();
 sg13g2_decap_8 FILLER_85_7 ();
 sg13g2_decap_8 FILLER_85_14 ();
 sg13g2_decap_8 FILLER_85_21 ();
 sg13g2_decap_8 FILLER_85_28 ();
 sg13g2_decap_8 FILLER_85_35 ();
 sg13g2_decap_8 FILLER_85_42 ();
 sg13g2_decap_8 FILLER_85_49 ();
 sg13g2_decap_8 FILLER_85_56 ();
 sg13g2_decap_8 FILLER_85_63 ();
 sg13g2_decap_8 FILLER_85_70 ();
 sg13g2_decap_8 FILLER_85_77 ();
 sg13g2_decap_8 FILLER_85_84 ();
 sg13g2_decap_8 FILLER_85_91 ();
 sg13g2_decap_8 FILLER_85_98 ();
 sg13g2_decap_8 FILLER_85_105 ();
 sg13g2_decap_8 FILLER_85_112 ();
 sg13g2_decap_8 FILLER_85_119 ();
 sg13g2_decap_8 FILLER_85_126 ();
 sg13g2_decap_8 FILLER_85_133 ();
 sg13g2_decap_8 FILLER_85_140 ();
 sg13g2_decap_8 FILLER_85_147 ();
 sg13g2_decap_8 FILLER_85_154 ();
 sg13g2_decap_8 FILLER_85_161 ();
 sg13g2_decap_8 FILLER_85_168 ();
 sg13g2_decap_8 FILLER_85_175 ();
 sg13g2_decap_8 FILLER_85_182 ();
 sg13g2_decap_8 FILLER_85_189 ();
 sg13g2_decap_8 FILLER_85_196 ();
 sg13g2_decap_8 FILLER_85_203 ();
 sg13g2_decap_8 FILLER_85_210 ();
 sg13g2_decap_8 FILLER_85_217 ();
 sg13g2_decap_8 FILLER_85_224 ();
 sg13g2_decap_8 FILLER_85_231 ();
 sg13g2_decap_8 FILLER_85_238 ();
 sg13g2_decap_8 FILLER_85_245 ();
 sg13g2_decap_8 FILLER_85_252 ();
 sg13g2_decap_8 FILLER_85_259 ();
 sg13g2_decap_8 FILLER_85_266 ();
 sg13g2_decap_8 FILLER_85_273 ();
 sg13g2_decap_8 FILLER_85_280 ();
 sg13g2_decap_8 FILLER_85_287 ();
 sg13g2_decap_8 FILLER_85_294 ();
 sg13g2_decap_8 FILLER_85_301 ();
 sg13g2_decap_8 FILLER_85_308 ();
 sg13g2_decap_8 FILLER_85_315 ();
 sg13g2_decap_8 FILLER_85_322 ();
 sg13g2_decap_8 FILLER_85_329 ();
 sg13g2_decap_8 FILLER_85_336 ();
 sg13g2_decap_8 FILLER_85_343 ();
 sg13g2_decap_8 FILLER_85_350 ();
 sg13g2_decap_8 FILLER_85_357 ();
 sg13g2_decap_8 FILLER_85_364 ();
 sg13g2_decap_8 FILLER_85_371 ();
 sg13g2_decap_8 FILLER_85_378 ();
 sg13g2_decap_8 FILLER_85_385 ();
 sg13g2_decap_8 FILLER_85_392 ();
 sg13g2_decap_8 FILLER_85_399 ();
 sg13g2_decap_8 FILLER_85_406 ();
 sg13g2_decap_8 FILLER_85_413 ();
 sg13g2_decap_8 FILLER_85_420 ();
 sg13g2_decap_8 FILLER_85_427 ();
 sg13g2_decap_8 FILLER_85_434 ();
 sg13g2_decap_8 FILLER_85_441 ();
 sg13g2_decap_8 FILLER_85_448 ();
 sg13g2_decap_8 FILLER_85_455 ();
 sg13g2_decap_8 FILLER_85_462 ();
 sg13g2_decap_8 FILLER_85_469 ();
 sg13g2_decap_8 FILLER_85_476 ();
 sg13g2_decap_8 FILLER_85_483 ();
 sg13g2_decap_8 FILLER_85_490 ();
 sg13g2_decap_8 FILLER_85_497 ();
 sg13g2_decap_8 FILLER_85_504 ();
 sg13g2_decap_8 FILLER_85_511 ();
 sg13g2_decap_8 FILLER_85_518 ();
 sg13g2_decap_8 FILLER_85_525 ();
 sg13g2_decap_8 FILLER_85_532 ();
 sg13g2_decap_8 FILLER_85_539 ();
 sg13g2_decap_8 FILLER_85_546 ();
 sg13g2_decap_8 FILLER_85_553 ();
 sg13g2_decap_8 FILLER_85_560 ();
 sg13g2_decap_8 FILLER_85_567 ();
 sg13g2_decap_8 FILLER_85_574 ();
 sg13g2_decap_8 FILLER_85_581 ();
 sg13g2_decap_8 FILLER_85_588 ();
 sg13g2_decap_8 FILLER_85_595 ();
 sg13g2_decap_8 FILLER_85_602 ();
 sg13g2_decap_8 FILLER_85_609 ();
 sg13g2_decap_8 FILLER_85_616 ();
 sg13g2_decap_8 FILLER_85_623 ();
 sg13g2_decap_8 FILLER_85_630 ();
 sg13g2_decap_8 FILLER_85_637 ();
 sg13g2_decap_8 FILLER_85_644 ();
 sg13g2_decap_8 FILLER_85_651 ();
 sg13g2_decap_8 FILLER_85_658 ();
 sg13g2_decap_8 FILLER_85_665 ();
 sg13g2_decap_8 FILLER_85_672 ();
 sg13g2_decap_8 FILLER_85_679 ();
 sg13g2_decap_8 FILLER_85_686 ();
 sg13g2_decap_8 FILLER_85_693 ();
 sg13g2_decap_8 FILLER_85_700 ();
 sg13g2_decap_8 FILLER_85_707 ();
 sg13g2_decap_8 FILLER_85_714 ();
 sg13g2_decap_8 FILLER_85_721 ();
 sg13g2_decap_8 FILLER_85_728 ();
 sg13g2_decap_8 FILLER_85_735 ();
 sg13g2_decap_8 FILLER_85_742 ();
 sg13g2_decap_8 FILLER_85_749 ();
 sg13g2_decap_8 FILLER_85_756 ();
 sg13g2_decap_8 FILLER_85_763 ();
 sg13g2_decap_8 FILLER_85_770 ();
 sg13g2_decap_8 FILLER_85_777 ();
 sg13g2_decap_8 FILLER_85_784 ();
 sg13g2_decap_8 FILLER_85_791 ();
 sg13g2_decap_8 FILLER_85_798 ();
 sg13g2_decap_8 FILLER_85_805 ();
 sg13g2_decap_8 FILLER_85_812 ();
 sg13g2_decap_8 FILLER_85_819 ();
 sg13g2_decap_8 FILLER_85_826 ();
 sg13g2_decap_8 FILLER_85_833 ();
 sg13g2_fill_1 FILLER_85_840 ();
 sg13g2_decap_8 FILLER_86_0 ();
 sg13g2_decap_8 FILLER_86_7 ();
 sg13g2_decap_8 FILLER_86_14 ();
 sg13g2_decap_8 FILLER_86_21 ();
 sg13g2_decap_8 FILLER_86_28 ();
 sg13g2_decap_8 FILLER_86_35 ();
 sg13g2_decap_8 FILLER_86_42 ();
 sg13g2_decap_8 FILLER_86_49 ();
 sg13g2_decap_8 FILLER_86_56 ();
 sg13g2_decap_8 FILLER_86_63 ();
 sg13g2_decap_8 FILLER_86_70 ();
 sg13g2_decap_8 FILLER_86_77 ();
 sg13g2_decap_8 FILLER_86_84 ();
 sg13g2_decap_8 FILLER_86_91 ();
 sg13g2_decap_8 FILLER_86_98 ();
 sg13g2_decap_8 FILLER_86_105 ();
 sg13g2_decap_8 FILLER_86_112 ();
 sg13g2_decap_8 FILLER_86_119 ();
 sg13g2_decap_8 FILLER_86_126 ();
 sg13g2_decap_8 FILLER_86_133 ();
 sg13g2_decap_8 FILLER_86_140 ();
 sg13g2_decap_8 FILLER_86_147 ();
 sg13g2_decap_8 FILLER_86_154 ();
 sg13g2_decap_8 FILLER_86_161 ();
 sg13g2_decap_8 FILLER_86_168 ();
 sg13g2_decap_8 FILLER_86_175 ();
 sg13g2_decap_8 FILLER_86_182 ();
 sg13g2_decap_8 FILLER_86_189 ();
 sg13g2_decap_8 FILLER_86_196 ();
 sg13g2_decap_8 FILLER_86_203 ();
 sg13g2_decap_8 FILLER_86_210 ();
 sg13g2_decap_8 FILLER_86_217 ();
 sg13g2_decap_8 FILLER_86_224 ();
 sg13g2_decap_8 FILLER_86_231 ();
 sg13g2_decap_8 FILLER_86_238 ();
 sg13g2_decap_8 FILLER_86_245 ();
 sg13g2_decap_8 FILLER_86_252 ();
 sg13g2_decap_8 FILLER_86_259 ();
 sg13g2_decap_8 FILLER_86_266 ();
 sg13g2_decap_8 FILLER_86_273 ();
 sg13g2_decap_8 FILLER_86_280 ();
 sg13g2_decap_8 FILLER_86_287 ();
 sg13g2_decap_8 FILLER_86_294 ();
 sg13g2_decap_8 FILLER_86_301 ();
 sg13g2_decap_8 FILLER_86_308 ();
 sg13g2_decap_8 FILLER_86_315 ();
 sg13g2_decap_8 FILLER_86_322 ();
 sg13g2_decap_8 FILLER_86_329 ();
 sg13g2_decap_8 FILLER_86_336 ();
 sg13g2_decap_8 FILLER_86_343 ();
 sg13g2_decap_8 FILLER_86_350 ();
 sg13g2_decap_8 FILLER_86_357 ();
 sg13g2_decap_8 FILLER_86_364 ();
 sg13g2_decap_8 FILLER_86_371 ();
 sg13g2_decap_8 FILLER_86_378 ();
 sg13g2_decap_8 FILLER_86_385 ();
 sg13g2_decap_8 FILLER_86_392 ();
 sg13g2_decap_8 FILLER_86_399 ();
 sg13g2_decap_8 FILLER_86_406 ();
 sg13g2_decap_8 FILLER_86_413 ();
 sg13g2_decap_8 FILLER_86_420 ();
 sg13g2_decap_8 FILLER_86_427 ();
 sg13g2_decap_8 FILLER_86_434 ();
 sg13g2_decap_8 FILLER_86_441 ();
 sg13g2_decap_8 FILLER_86_448 ();
 sg13g2_decap_8 FILLER_86_455 ();
 sg13g2_decap_8 FILLER_86_462 ();
 sg13g2_decap_8 FILLER_86_469 ();
 sg13g2_decap_8 FILLER_86_476 ();
 sg13g2_decap_8 FILLER_86_483 ();
 sg13g2_decap_8 FILLER_86_490 ();
 sg13g2_decap_8 FILLER_86_497 ();
 sg13g2_decap_8 FILLER_86_504 ();
 sg13g2_decap_8 FILLER_86_511 ();
 sg13g2_decap_8 FILLER_86_518 ();
 sg13g2_decap_8 FILLER_86_525 ();
 sg13g2_decap_8 FILLER_86_532 ();
 sg13g2_decap_8 FILLER_86_539 ();
 sg13g2_decap_8 FILLER_86_546 ();
 sg13g2_decap_8 FILLER_86_553 ();
 sg13g2_decap_8 FILLER_86_560 ();
 sg13g2_decap_8 FILLER_86_567 ();
 sg13g2_decap_8 FILLER_86_574 ();
 sg13g2_decap_8 FILLER_86_581 ();
 sg13g2_decap_8 FILLER_86_588 ();
 sg13g2_decap_8 FILLER_86_595 ();
 sg13g2_decap_8 FILLER_86_602 ();
 sg13g2_decap_8 FILLER_86_609 ();
 sg13g2_decap_8 FILLER_86_616 ();
 sg13g2_decap_8 FILLER_86_623 ();
 sg13g2_decap_8 FILLER_86_630 ();
 sg13g2_decap_8 FILLER_86_637 ();
 sg13g2_decap_8 FILLER_86_644 ();
 sg13g2_decap_8 FILLER_86_651 ();
 sg13g2_decap_8 FILLER_86_658 ();
 sg13g2_decap_8 FILLER_86_665 ();
 sg13g2_decap_8 FILLER_86_672 ();
 sg13g2_decap_8 FILLER_86_679 ();
 sg13g2_decap_8 FILLER_86_686 ();
 sg13g2_decap_8 FILLER_86_693 ();
 sg13g2_decap_8 FILLER_86_700 ();
 sg13g2_decap_8 FILLER_86_707 ();
 sg13g2_decap_8 FILLER_86_714 ();
 sg13g2_decap_8 FILLER_86_721 ();
 sg13g2_decap_8 FILLER_86_728 ();
 sg13g2_decap_8 FILLER_86_735 ();
 sg13g2_decap_8 FILLER_86_742 ();
 sg13g2_decap_8 FILLER_86_749 ();
 sg13g2_decap_8 FILLER_86_756 ();
 sg13g2_decap_8 FILLER_86_763 ();
 sg13g2_decap_8 FILLER_86_770 ();
 sg13g2_decap_8 FILLER_86_777 ();
 sg13g2_decap_8 FILLER_86_784 ();
 sg13g2_decap_8 FILLER_86_791 ();
 sg13g2_decap_8 FILLER_86_798 ();
 sg13g2_decap_8 FILLER_86_805 ();
 sg13g2_decap_8 FILLER_86_812 ();
 sg13g2_decap_8 FILLER_86_819 ();
 sg13g2_decap_8 FILLER_86_826 ();
 sg13g2_decap_8 FILLER_86_833 ();
 sg13g2_fill_1 FILLER_86_840 ();
 sg13g2_decap_8 FILLER_87_0 ();
 sg13g2_decap_8 FILLER_87_7 ();
 sg13g2_decap_8 FILLER_87_14 ();
 sg13g2_decap_8 FILLER_87_21 ();
 sg13g2_decap_8 FILLER_87_28 ();
 sg13g2_decap_8 FILLER_87_35 ();
 sg13g2_decap_8 FILLER_87_42 ();
 sg13g2_decap_8 FILLER_87_49 ();
 sg13g2_decap_8 FILLER_87_56 ();
 sg13g2_decap_8 FILLER_87_63 ();
 sg13g2_decap_8 FILLER_87_70 ();
 sg13g2_decap_8 FILLER_87_77 ();
 sg13g2_decap_8 FILLER_87_84 ();
 sg13g2_decap_8 FILLER_87_91 ();
 sg13g2_decap_8 FILLER_87_98 ();
 sg13g2_decap_8 FILLER_87_105 ();
 sg13g2_decap_8 FILLER_87_112 ();
 sg13g2_decap_8 FILLER_87_119 ();
 sg13g2_decap_8 FILLER_87_126 ();
 sg13g2_decap_8 FILLER_87_133 ();
 sg13g2_decap_8 FILLER_87_140 ();
 sg13g2_decap_8 FILLER_87_147 ();
 sg13g2_decap_8 FILLER_87_154 ();
 sg13g2_decap_8 FILLER_87_161 ();
 sg13g2_decap_8 FILLER_87_168 ();
 sg13g2_decap_8 FILLER_87_175 ();
 sg13g2_decap_8 FILLER_87_182 ();
 sg13g2_decap_8 FILLER_87_189 ();
 sg13g2_decap_8 FILLER_87_196 ();
 sg13g2_decap_8 FILLER_87_203 ();
 sg13g2_decap_8 FILLER_87_210 ();
 sg13g2_decap_8 FILLER_87_217 ();
 sg13g2_decap_8 FILLER_87_224 ();
 sg13g2_decap_8 FILLER_87_231 ();
 sg13g2_decap_8 FILLER_87_238 ();
 sg13g2_decap_8 FILLER_87_245 ();
 sg13g2_decap_8 FILLER_87_252 ();
 sg13g2_decap_8 FILLER_87_259 ();
 sg13g2_decap_8 FILLER_87_266 ();
 sg13g2_decap_8 FILLER_87_273 ();
 sg13g2_decap_8 FILLER_87_280 ();
 sg13g2_decap_8 FILLER_87_287 ();
 sg13g2_decap_8 FILLER_87_294 ();
 sg13g2_decap_8 FILLER_87_301 ();
 sg13g2_decap_8 FILLER_87_308 ();
 sg13g2_decap_8 FILLER_87_315 ();
 sg13g2_decap_8 FILLER_87_322 ();
 sg13g2_decap_8 FILLER_87_329 ();
 sg13g2_decap_8 FILLER_87_336 ();
 sg13g2_decap_8 FILLER_87_343 ();
 sg13g2_decap_8 FILLER_87_350 ();
 sg13g2_decap_8 FILLER_87_357 ();
 sg13g2_decap_8 FILLER_87_364 ();
 sg13g2_decap_8 FILLER_87_371 ();
 sg13g2_decap_8 FILLER_87_378 ();
 sg13g2_decap_8 FILLER_87_385 ();
 sg13g2_decap_8 FILLER_87_392 ();
 sg13g2_decap_8 FILLER_87_399 ();
 sg13g2_decap_8 FILLER_87_406 ();
 sg13g2_decap_8 FILLER_87_413 ();
 sg13g2_decap_8 FILLER_87_420 ();
 sg13g2_decap_8 FILLER_87_427 ();
 sg13g2_decap_8 FILLER_87_434 ();
 sg13g2_decap_8 FILLER_87_441 ();
 sg13g2_decap_8 FILLER_87_448 ();
 sg13g2_decap_8 FILLER_87_455 ();
 sg13g2_decap_8 FILLER_87_462 ();
 sg13g2_decap_8 FILLER_87_469 ();
 sg13g2_decap_8 FILLER_87_476 ();
 sg13g2_decap_8 FILLER_87_483 ();
 sg13g2_decap_8 FILLER_87_490 ();
 sg13g2_decap_8 FILLER_87_497 ();
 sg13g2_decap_8 FILLER_87_504 ();
 sg13g2_decap_8 FILLER_87_511 ();
 sg13g2_decap_8 FILLER_87_518 ();
 sg13g2_decap_8 FILLER_87_525 ();
 sg13g2_decap_8 FILLER_87_532 ();
 sg13g2_decap_8 FILLER_87_539 ();
 sg13g2_decap_8 FILLER_87_546 ();
 sg13g2_decap_8 FILLER_87_553 ();
 sg13g2_decap_8 FILLER_87_560 ();
 sg13g2_decap_8 FILLER_87_567 ();
 sg13g2_decap_8 FILLER_87_574 ();
 sg13g2_decap_8 FILLER_87_581 ();
 sg13g2_decap_8 FILLER_87_588 ();
 sg13g2_decap_8 FILLER_87_595 ();
 sg13g2_decap_8 FILLER_87_602 ();
 sg13g2_decap_8 FILLER_87_609 ();
 sg13g2_decap_8 FILLER_87_616 ();
 sg13g2_decap_8 FILLER_87_623 ();
 sg13g2_decap_8 FILLER_87_630 ();
 sg13g2_decap_8 FILLER_87_637 ();
 sg13g2_decap_8 FILLER_87_644 ();
 sg13g2_decap_8 FILLER_87_651 ();
 sg13g2_decap_8 FILLER_87_658 ();
 sg13g2_decap_8 FILLER_87_665 ();
 sg13g2_decap_8 FILLER_87_672 ();
 sg13g2_decap_8 FILLER_87_679 ();
 sg13g2_decap_8 FILLER_87_686 ();
 sg13g2_decap_8 FILLER_87_693 ();
 sg13g2_decap_8 FILLER_87_700 ();
 sg13g2_decap_8 FILLER_87_707 ();
 sg13g2_decap_8 FILLER_87_714 ();
 sg13g2_decap_8 FILLER_87_721 ();
 sg13g2_decap_8 FILLER_87_728 ();
 sg13g2_decap_8 FILLER_87_735 ();
 sg13g2_decap_8 FILLER_87_742 ();
 sg13g2_decap_8 FILLER_87_749 ();
 sg13g2_decap_8 FILLER_87_756 ();
 sg13g2_decap_8 FILLER_87_763 ();
 sg13g2_decap_8 FILLER_87_770 ();
 sg13g2_decap_8 FILLER_87_777 ();
 sg13g2_decap_8 FILLER_87_784 ();
 sg13g2_decap_8 FILLER_87_791 ();
 sg13g2_decap_8 FILLER_87_798 ();
 sg13g2_decap_8 FILLER_87_805 ();
 sg13g2_decap_8 FILLER_87_812 ();
 sg13g2_decap_8 FILLER_87_819 ();
 sg13g2_decap_8 FILLER_87_826 ();
 sg13g2_decap_8 FILLER_87_833 ();
 sg13g2_fill_1 FILLER_87_840 ();
 sg13g2_decap_8 FILLER_88_0 ();
 sg13g2_decap_8 FILLER_88_7 ();
 sg13g2_decap_8 FILLER_88_14 ();
 sg13g2_decap_8 FILLER_88_21 ();
 sg13g2_decap_8 FILLER_88_28 ();
 sg13g2_decap_8 FILLER_88_35 ();
 sg13g2_decap_8 FILLER_88_42 ();
 sg13g2_decap_8 FILLER_88_49 ();
 sg13g2_decap_8 FILLER_88_56 ();
 sg13g2_decap_8 FILLER_88_63 ();
 sg13g2_decap_8 FILLER_88_70 ();
 sg13g2_decap_8 FILLER_88_77 ();
 sg13g2_decap_8 FILLER_88_84 ();
 sg13g2_decap_8 FILLER_88_91 ();
 sg13g2_decap_8 FILLER_88_98 ();
 sg13g2_decap_8 FILLER_88_105 ();
 sg13g2_decap_8 FILLER_88_112 ();
 sg13g2_decap_8 FILLER_88_119 ();
 sg13g2_decap_8 FILLER_88_126 ();
 sg13g2_decap_8 FILLER_88_133 ();
 sg13g2_decap_8 FILLER_88_140 ();
 sg13g2_decap_8 FILLER_88_147 ();
 sg13g2_decap_8 FILLER_88_154 ();
 sg13g2_decap_8 FILLER_88_161 ();
 sg13g2_decap_8 FILLER_88_168 ();
 sg13g2_decap_8 FILLER_88_175 ();
 sg13g2_decap_8 FILLER_88_182 ();
 sg13g2_decap_8 FILLER_88_189 ();
 sg13g2_decap_8 FILLER_88_196 ();
 sg13g2_decap_8 FILLER_88_203 ();
 sg13g2_decap_8 FILLER_88_210 ();
 sg13g2_decap_8 FILLER_88_217 ();
 sg13g2_decap_8 FILLER_88_224 ();
 sg13g2_decap_8 FILLER_88_231 ();
 sg13g2_decap_8 FILLER_88_238 ();
 sg13g2_decap_8 FILLER_88_245 ();
 sg13g2_decap_8 FILLER_88_252 ();
 sg13g2_decap_8 FILLER_88_259 ();
 sg13g2_decap_8 FILLER_88_266 ();
 sg13g2_decap_8 FILLER_88_273 ();
 sg13g2_decap_8 FILLER_88_280 ();
 sg13g2_decap_8 FILLER_88_287 ();
 sg13g2_decap_8 FILLER_88_294 ();
 sg13g2_decap_8 FILLER_88_301 ();
 sg13g2_decap_8 FILLER_88_308 ();
 sg13g2_decap_8 FILLER_88_315 ();
 sg13g2_decap_8 FILLER_88_322 ();
 sg13g2_decap_8 FILLER_88_329 ();
 sg13g2_decap_8 FILLER_88_336 ();
 sg13g2_decap_8 FILLER_88_343 ();
 sg13g2_decap_8 FILLER_88_350 ();
 sg13g2_decap_8 FILLER_88_357 ();
 sg13g2_decap_8 FILLER_88_364 ();
 sg13g2_decap_8 FILLER_88_371 ();
 sg13g2_decap_8 FILLER_88_378 ();
 sg13g2_decap_8 FILLER_88_385 ();
 sg13g2_decap_8 FILLER_88_392 ();
 sg13g2_decap_8 FILLER_88_399 ();
 sg13g2_decap_8 FILLER_88_406 ();
 sg13g2_decap_8 FILLER_88_413 ();
 sg13g2_decap_8 FILLER_88_420 ();
 sg13g2_decap_8 FILLER_88_427 ();
 sg13g2_decap_8 FILLER_88_434 ();
 sg13g2_decap_8 FILLER_88_441 ();
 sg13g2_decap_8 FILLER_88_448 ();
 sg13g2_decap_8 FILLER_88_455 ();
 sg13g2_decap_8 FILLER_88_462 ();
 sg13g2_decap_8 FILLER_88_469 ();
 sg13g2_decap_8 FILLER_88_476 ();
 sg13g2_decap_8 FILLER_88_483 ();
 sg13g2_decap_8 FILLER_88_490 ();
 sg13g2_decap_8 FILLER_88_497 ();
 sg13g2_decap_8 FILLER_88_504 ();
 sg13g2_decap_8 FILLER_88_511 ();
 sg13g2_decap_8 FILLER_88_518 ();
 sg13g2_decap_8 FILLER_88_525 ();
 sg13g2_decap_8 FILLER_88_532 ();
 sg13g2_decap_8 FILLER_88_539 ();
 sg13g2_decap_8 FILLER_88_546 ();
 sg13g2_decap_8 FILLER_88_553 ();
 sg13g2_decap_8 FILLER_88_560 ();
 sg13g2_decap_8 FILLER_88_567 ();
 sg13g2_decap_8 FILLER_88_574 ();
 sg13g2_decap_8 FILLER_88_581 ();
 sg13g2_decap_8 FILLER_88_588 ();
 sg13g2_decap_8 FILLER_88_595 ();
 sg13g2_decap_8 FILLER_88_602 ();
 sg13g2_decap_8 FILLER_88_609 ();
 sg13g2_decap_8 FILLER_88_616 ();
 sg13g2_decap_8 FILLER_88_623 ();
 sg13g2_decap_8 FILLER_88_630 ();
 sg13g2_decap_8 FILLER_88_637 ();
 sg13g2_decap_8 FILLER_88_644 ();
 sg13g2_decap_8 FILLER_88_651 ();
 sg13g2_decap_8 FILLER_88_658 ();
 sg13g2_decap_8 FILLER_88_665 ();
 sg13g2_decap_8 FILLER_88_672 ();
 sg13g2_decap_8 FILLER_88_679 ();
 sg13g2_decap_8 FILLER_88_686 ();
 sg13g2_decap_8 FILLER_88_693 ();
 sg13g2_decap_8 FILLER_88_700 ();
 sg13g2_decap_8 FILLER_88_707 ();
 sg13g2_decap_8 FILLER_88_714 ();
 sg13g2_decap_8 FILLER_88_721 ();
 sg13g2_decap_8 FILLER_88_728 ();
 sg13g2_decap_8 FILLER_88_735 ();
 sg13g2_decap_8 FILLER_88_742 ();
 sg13g2_decap_8 FILLER_88_749 ();
 sg13g2_decap_8 FILLER_88_756 ();
 sg13g2_decap_8 FILLER_88_763 ();
 sg13g2_decap_8 FILLER_88_770 ();
 sg13g2_decap_8 FILLER_88_777 ();
 sg13g2_decap_8 FILLER_88_784 ();
 sg13g2_decap_8 FILLER_88_791 ();
 sg13g2_decap_8 FILLER_88_798 ();
 sg13g2_decap_8 FILLER_88_805 ();
 sg13g2_decap_8 FILLER_88_812 ();
 sg13g2_decap_8 FILLER_88_819 ();
 sg13g2_decap_8 FILLER_88_826 ();
 sg13g2_decap_8 FILLER_88_833 ();
 sg13g2_fill_1 FILLER_88_840 ();
 sg13g2_decap_8 FILLER_89_0 ();
 sg13g2_decap_8 FILLER_89_7 ();
 sg13g2_decap_8 FILLER_89_14 ();
 sg13g2_decap_8 FILLER_89_21 ();
 sg13g2_decap_8 FILLER_89_28 ();
 sg13g2_decap_8 FILLER_89_35 ();
 sg13g2_decap_8 FILLER_89_42 ();
 sg13g2_decap_8 FILLER_89_49 ();
 sg13g2_decap_8 FILLER_89_56 ();
 sg13g2_decap_8 FILLER_89_63 ();
 sg13g2_decap_8 FILLER_89_70 ();
 sg13g2_decap_8 FILLER_89_77 ();
 sg13g2_decap_8 FILLER_89_84 ();
 sg13g2_decap_8 FILLER_89_91 ();
 sg13g2_decap_8 FILLER_89_98 ();
 sg13g2_decap_8 FILLER_89_105 ();
 sg13g2_decap_8 FILLER_89_112 ();
 sg13g2_decap_8 FILLER_89_119 ();
 sg13g2_decap_8 FILLER_89_126 ();
 sg13g2_decap_8 FILLER_89_133 ();
 sg13g2_decap_8 FILLER_89_140 ();
 sg13g2_decap_8 FILLER_89_147 ();
 sg13g2_decap_8 FILLER_89_154 ();
 sg13g2_decap_8 FILLER_89_161 ();
 sg13g2_decap_8 FILLER_89_168 ();
 sg13g2_decap_8 FILLER_89_175 ();
 sg13g2_decap_8 FILLER_89_182 ();
 sg13g2_decap_8 FILLER_89_189 ();
 sg13g2_decap_8 FILLER_89_196 ();
 sg13g2_decap_8 FILLER_89_203 ();
 sg13g2_decap_8 FILLER_89_210 ();
 sg13g2_decap_8 FILLER_89_217 ();
 sg13g2_decap_8 FILLER_89_224 ();
 sg13g2_decap_8 FILLER_89_231 ();
 sg13g2_decap_8 FILLER_89_238 ();
 sg13g2_decap_8 FILLER_89_245 ();
 sg13g2_decap_8 FILLER_89_252 ();
 sg13g2_decap_8 FILLER_89_259 ();
 sg13g2_decap_8 FILLER_89_266 ();
 sg13g2_decap_8 FILLER_89_273 ();
 sg13g2_decap_8 FILLER_89_280 ();
 sg13g2_decap_8 FILLER_89_287 ();
 sg13g2_decap_8 FILLER_89_294 ();
 sg13g2_decap_8 FILLER_89_301 ();
 sg13g2_decap_8 FILLER_89_308 ();
 sg13g2_decap_8 FILLER_89_315 ();
 sg13g2_decap_8 FILLER_89_322 ();
 sg13g2_decap_8 FILLER_89_329 ();
 sg13g2_decap_8 FILLER_89_336 ();
 sg13g2_decap_8 FILLER_89_343 ();
 sg13g2_decap_8 FILLER_89_350 ();
 sg13g2_decap_8 FILLER_89_357 ();
 sg13g2_decap_8 FILLER_89_364 ();
 sg13g2_decap_8 FILLER_89_371 ();
 sg13g2_decap_8 FILLER_89_378 ();
 sg13g2_decap_8 FILLER_89_385 ();
 sg13g2_decap_8 FILLER_89_392 ();
 sg13g2_decap_8 FILLER_89_399 ();
 sg13g2_decap_8 FILLER_89_406 ();
 sg13g2_decap_8 FILLER_89_413 ();
 sg13g2_decap_8 FILLER_89_420 ();
 sg13g2_decap_8 FILLER_89_427 ();
 sg13g2_decap_8 FILLER_89_434 ();
 sg13g2_decap_8 FILLER_89_441 ();
 sg13g2_decap_8 FILLER_89_448 ();
 sg13g2_decap_8 FILLER_89_455 ();
 sg13g2_decap_8 FILLER_89_462 ();
 sg13g2_decap_8 FILLER_89_469 ();
 sg13g2_decap_8 FILLER_89_476 ();
 sg13g2_decap_8 FILLER_89_483 ();
 sg13g2_decap_8 FILLER_89_490 ();
 sg13g2_decap_8 FILLER_89_497 ();
 sg13g2_decap_8 FILLER_89_504 ();
 sg13g2_decap_8 FILLER_89_511 ();
 sg13g2_decap_8 FILLER_89_518 ();
 sg13g2_decap_8 FILLER_89_525 ();
 sg13g2_decap_8 FILLER_89_532 ();
 sg13g2_decap_8 FILLER_89_539 ();
 sg13g2_decap_8 FILLER_89_546 ();
 sg13g2_decap_8 FILLER_89_553 ();
 sg13g2_decap_8 FILLER_89_560 ();
 sg13g2_decap_8 FILLER_89_567 ();
 sg13g2_decap_8 FILLER_89_574 ();
 sg13g2_decap_8 FILLER_89_581 ();
 sg13g2_decap_8 FILLER_89_588 ();
 sg13g2_decap_8 FILLER_89_595 ();
 sg13g2_decap_8 FILLER_89_602 ();
 sg13g2_decap_8 FILLER_89_609 ();
 sg13g2_decap_8 FILLER_89_616 ();
 sg13g2_decap_8 FILLER_89_623 ();
 sg13g2_decap_8 FILLER_89_630 ();
 sg13g2_decap_8 FILLER_89_637 ();
 sg13g2_decap_8 FILLER_89_644 ();
 sg13g2_decap_8 FILLER_89_651 ();
 sg13g2_decap_8 FILLER_89_658 ();
 sg13g2_decap_8 FILLER_89_665 ();
 sg13g2_decap_8 FILLER_89_672 ();
 sg13g2_decap_8 FILLER_89_679 ();
 sg13g2_decap_8 FILLER_89_686 ();
 sg13g2_decap_8 FILLER_89_693 ();
 sg13g2_decap_8 FILLER_89_700 ();
 sg13g2_decap_8 FILLER_89_707 ();
 sg13g2_decap_8 FILLER_89_714 ();
 sg13g2_decap_8 FILLER_89_721 ();
 sg13g2_decap_8 FILLER_89_728 ();
 sg13g2_decap_8 FILLER_89_735 ();
 sg13g2_decap_8 FILLER_89_742 ();
 sg13g2_decap_8 FILLER_89_749 ();
 sg13g2_decap_8 FILLER_89_756 ();
 sg13g2_decap_8 FILLER_89_763 ();
 sg13g2_decap_8 FILLER_89_770 ();
 sg13g2_decap_8 FILLER_89_777 ();
 sg13g2_decap_8 FILLER_89_784 ();
 sg13g2_decap_8 FILLER_89_791 ();
 sg13g2_decap_8 FILLER_89_798 ();
 sg13g2_decap_8 FILLER_89_805 ();
 sg13g2_decap_8 FILLER_89_812 ();
 sg13g2_decap_8 FILLER_89_819 ();
 sg13g2_decap_8 FILLER_89_826 ();
 sg13g2_decap_8 FILLER_89_833 ();
 sg13g2_fill_1 FILLER_89_840 ();
 sg13g2_decap_8 FILLER_90_0 ();
 sg13g2_decap_8 FILLER_90_7 ();
 sg13g2_decap_8 FILLER_90_14 ();
 sg13g2_decap_8 FILLER_90_21 ();
 sg13g2_decap_8 FILLER_90_28 ();
 sg13g2_decap_8 FILLER_90_35 ();
 sg13g2_decap_8 FILLER_90_42 ();
 sg13g2_decap_8 FILLER_90_49 ();
 sg13g2_decap_8 FILLER_90_56 ();
 sg13g2_decap_8 FILLER_90_63 ();
 sg13g2_decap_8 FILLER_90_70 ();
 sg13g2_decap_8 FILLER_90_77 ();
 sg13g2_decap_8 FILLER_90_84 ();
 sg13g2_decap_8 FILLER_90_91 ();
 sg13g2_decap_8 FILLER_90_98 ();
 sg13g2_decap_8 FILLER_90_105 ();
 sg13g2_decap_8 FILLER_90_112 ();
 sg13g2_decap_8 FILLER_90_119 ();
 sg13g2_decap_8 FILLER_90_126 ();
 sg13g2_decap_8 FILLER_90_133 ();
 sg13g2_decap_8 FILLER_90_140 ();
 sg13g2_decap_8 FILLER_90_147 ();
 sg13g2_decap_8 FILLER_90_154 ();
 sg13g2_decap_8 FILLER_90_161 ();
 sg13g2_decap_8 FILLER_90_168 ();
 sg13g2_decap_8 FILLER_90_175 ();
 sg13g2_decap_8 FILLER_90_182 ();
 sg13g2_decap_8 FILLER_90_189 ();
 sg13g2_decap_8 FILLER_90_196 ();
 sg13g2_decap_8 FILLER_90_203 ();
 sg13g2_decap_8 FILLER_90_210 ();
 sg13g2_decap_8 FILLER_90_217 ();
 sg13g2_decap_8 FILLER_90_224 ();
 sg13g2_decap_8 FILLER_90_231 ();
 sg13g2_decap_8 FILLER_90_238 ();
 sg13g2_decap_8 FILLER_90_245 ();
 sg13g2_decap_8 FILLER_90_252 ();
 sg13g2_decap_8 FILLER_90_259 ();
 sg13g2_decap_8 FILLER_90_266 ();
 sg13g2_decap_8 FILLER_90_273 ();
 sg13g2_decap_8 FILLER_90_280 ();
 sg13g2_decap_8 FILLER_90_287 ();
 sg13g2_decap_8 FILLER_90_294 ();
 sg13g2_decap_8 FILLER_90_301 ();
 sg13g2_decap_8 FILLER_90_308 ();
 sg13g2_decap_8 FILLER_90_315 ();
 sg13g2_decap_8 FILLER_90_322 ();
 sg13g2_decap_8 FILLER_90_329 ();
 sg13g2_decap_8 FILLER_90_336 ();
 sg13g2_decap_8 FILLER_90_343 ();
 sg13g2_decap_8 FILLER_90_350 ();
 sg13g2_decap_8 FILLER_90_357 ();
 sg13g2_decap_8 FILLER_90_364 ();
 sg13g2_decap_8 FILLER_90_371 ();
 sg13g2_decap_8 FILLER_90_378 ();
 sg13g2_decap_8 FILLER_90_385 ();
 sg13g2_decap_8 FILLER_90_392 ();
 sg13g2_decap_8 FILLER_90_399 ();
 sg13g2_decap_8 FILLER_90_406 ();
 sg13g2_decap_8 FILLER_90_413 ();
 sg13g2_decap_8 FILLER_90_420 ();
 sg13g2_decap_8 FILLER_90_427 ();
 sg13g2_decap_8 FILLER_90_434 ();
 sg13g2_decap_8 FILLER_90_441 ();
 sg13g2_decap_8 FILLER_90_448 ();
 sg13g2_decap_8 FILLER_90_455 ();
 sg13g2_decap_8 FILLER_90_462 ();
 sg13g2_decap_8 FILLER_90_469 ();
 sg13g2_decap_8 FILLER_90_476 ();
 sg13g2_decap_8 FILLER_90_483 ();
 sg13g2_decap_8 FILLER_90_490 ();
 sg13g2_decap_8 FILLER_90_497 ();
 sg13g2_decap_8 FILLER_90_504 ();
 sg13g2_decap_8 FILLER_90_511 ();
 sg13g2_decap_8 FILLER_90_518 ();
 sg13g2_decap_8 FILLER_90_525 ();
 sg13g2_decap_8 FILLER_90_532 ();
 sg13g2_decap_8 FILLER_90_539 ();
 sg13g2_decap_8 FILLER_90_546 ();
 sg13g2_decap_8 FILLER_90_553 ();
 sg13g2_decap_8 FILLER_90_560 ();
 sg13g2_decap_8 FILLER_90_567 ();
 sg13g2_decap_8 FILLER_90_574 ();
 sg13g2_decap_8 FILLER_90_581 ();
 sg13g2_decap_8 FILLER_90_588 ();
 sg13g2_decap_8 FILLER_90_595 ();
 sg13g2_decap_8 FILLER_90_602 ();
 sg13g2_decap_8 FILLER_90_609 ();
 sg13g2_decap_8 FILLER_90_616 ();
 sg13g2_decap_8 FILLER_90_623 ();
 sg13g2_decap_8 FILLER_90_630 ();
 sg13g2_decap_8 FILLER_90_637 ();
 sg13g2_decap_8 FILLER_90_644 ();
 sg13g2_decap_8 FILLER_90_651 ();
 sg13g2_decap_8 FILLER_90_658 ();
 sg13g2_decap_8 FILLER_90_665 ();
 sg13g2_decap_8 FILLER_90_672 ();
 sg13g2_decap_8 FILLER_90_679 ();
 sg13g2_decap_8 FILLER_90_686 ();
 sg13g2_decap_8 FILLER_90_693 ();
 sg13g2_decap_8 FILLER_90_700 ();
 sg13g2_decap_8 FILLER_90_707 ();
 sg13g2_decap_8 FILLER_90_714 ();
 sg13g2_decap_8 FILLER_90_721 ();
 sg13g2_decap_8 FILLER_90_728 ();
 sg13g2_decap_8 FILLER_90_735 ();
 sg13g2_decap_8 FILLER_90_742 ();
 sg13g2_decap_8 FILLER_90_749 ();
 sg13g2_decap_8 FILLER_90_756 ();
 sg13g2_decap_8 FILLER_90_763 ();
 sg13g2_decap_8 FILLER_90_770 ();
 sg13g2_decap_8 FILLER_90_777 ();
 sg13g2_decap_8 FILLER_90_784 ();
 sg13g2_decap_8 FILLER_90_791 ();
 sg13g2_decap_8 FILLER_90_798 ();
 sg13g2_decap_8 FILLER_90_805 ();
 sg13g2_decap_8 FILLER_90_812 ();
 sg13g2_decap_8 FILLER_90_819 ();
 sg13g2_decap_8 FILLER_90_826 ();
 sg13g2_decap_8 FILLER_90_833 ();
 sg13g2_fill_1 FILLER_90_840 ();
 sg13g2_decap_8 FILLER_91_0 ();
 sg13g2_decap_8 FILLER_91_7 ();
 sg13g2_decap_8 FILLER_91_14 ();
 sg13g2_decap_8 FILLER_91_21 ();
 sg13g2_decap_8 FILLER_91_28 ();
 sg13g2_decap_8 FILLER_91_35 ();
 sg13g2_decap_8 FILLER_91_42 ();
 sg13g2_decap_8 FILLER_91_49 ();
 sg13g2_decap_8 FILLER_91_56 ();
 sg13g2_decap_8 FILLER_91_63 ();
 sg13g2_decap_8 FILLER_91_70 ();
 sg13g2_decap_8 FILLER_91_77 ();
 sg13g2_decap_8 FILLER_91_84 ();
 sg13g2_decap_8 FILLER_91_91 ();
 sg13g2_decap_8 FILLER_91_98 ();
 sg13g2_decap_8 FILLER_91_105 ();
 sg13g2_decap_8 FILLER_91_112 ();
 sg13g2_decap_8 FILLER_91_119 ();
 sg13g2_decap_8 FILLER_91_126 ();
 sg13g2_decap_8 FILLER_91_133 ();
 sg13g2_decap_8 FILLER_91_140 ();
 sg13g2_decap_8 FILLER_91_147 ();
 sg13g2_decap_8 FILLER_91_154 ();
 sg13g2_decap_8 FILLER_91_161 ();
 sg13g2_decap_8 FILLER_91_168 ();
 sg13g2_decap_8 FILLER_91_175 ();
 sg13g2_decap_8 FILLER_91_182 ();
 sg13g2_decap_8 FILLER_91_189 ();
 sg13g2_decap_8 FILLER_91_196 ();
 sg13g2_decap_8 FILLER_91_203 ();
 sg13g2_decap_8 FILLER_91_210 ();
 sg13g2_decap_8 FILLER_91_217 ();
 sg13g2_decap_8 FILLER_91_224 ();
 sg13g2_decap_8 FILLER_91_231 ();
 sg13g2_decap_8 FILLER_91_238 ();
 sg13g2_decap_8 FILLER_91_245 ();
 sg13g2_decap_8 FILLER_91_252 ();
 sg13g2_decap_8 FILLER_91_259 ();
 sg13g2_decap_8 FILLER_91_266 ();
 sg13g2_decap_8 FILLER_91_273 ();
 sg13g2_decap_8 FILLER_91_280 ();
 sg13g2_decap_8 FILLER_91_287 ();
 sg13g2_decap_8 FILLER_91_294 ();
 sg13g2_decap_8 FILLER_91_301 ();
 sg13g2_decap_8 FILLER_91_308 ();
 sg13g2_decap_8 FILLER_91_315 ();
 sg13g2_decap_8 FILLER_91_322 ();
 sg13g2_decap_8 FILLER_91_329 ();
 sg13g2_decap_8 FILLER_91_336 ();
 sg13g2_decap_8 FILLER_91_343 ();
 sg13g2_decap_8 FILLER_91_350 ();
 sg13g2_decap_8 FILLER_91_357 ();
 sg13g2_decap_8 FILLER_91_364 ();
 sg13g2_decap_8 FILLER_91_371 ();
 sg13g2_decap_8 FILLER_91_378 ();
 sg13g2_decap_8 FILLER_91_385 ();
 sg13g2_decap_8 FILLER_91_392 ();
 sg13g2_decap_8 FILLER_91_399 ();
 sg13g2_decap_8 FILLER_91_406 ();
 sg13g2_decap_8 FILLER_91_413 ();
 sg13g2_decap_8 FILLER_91_420 ();
 sg13g2_decap_8 FILLER_91_427 ();
 sg13g2_decap_8 FILLER_91_434 ();
 sg13g2_decap_8 FILLER_91_441 ();
 sg13g2_decap_8 FILLER_91_448 ();
 sg13g2_decap_8 FILLER_91_455 ();
 sg13g2_decap_8 FILLER_91_462 ();
 sg13g2_decap_8 FILLER_91_469 ();
 sg13g2_decap_8 FILLER_91_476 ();
 sg13g2_decap_8 FILLER_91_483 ();
 sg13g2_decap_8 FILLER_91_490 ();
 sg13g2_decap_8 FILLER_91_497 ();
 sg13g2_decap_8 FILLER_91_504 ();
 sg13g2_decap_8 FILLER_91_511 ();
 sg13g2_decap_8 FILLER_91_518 ();
 sg13g2_decap_8 FILLER_91_525 ();
 sg13g2_decap_8 FILLER_91_532 ();
 sg13g2_decap_8 FILLER_91_539 ();
 sg13g2_decap_8 FILLER_91_546 ();
 sg13g2_decap_8 FILLER_91_553 ();
 sg13g2_decap_8 FILLER_91_560 ();
 sg13g2_decap_8 FILLER_91_567 ();
 sg13g2_decap_8 FILLER_91_574 ();
 sg13g2_decap_8 FILLER_91_581 ();
 sg13g2_decap_8 FILLER_91_588 ();
 sg13g2_decap_8 FILLER_91_595 ();
 sg13g2_decap_8 FILLER_91_602 ();
 sg13g2_decap_8 FILLER_91_609 ();
 sg13g2_decap_8 FILLER_91_616 ();
 sg13g2_decap_8 FILLER_91_623 ();
 sg13g2_decap_8 FILLER_91_630 ();
 sg13g2_decap_8 FILLER_91_637 ();
 sg13g2_decap_8 FILLER_91_644 ();
 sg13g2_decap_8 FILLER_91_651 ();
 sg13g2_decap_8 FILLER_91_658 ();
 sg13g2_decap_8 FILLER_91_665 ();
 sg13g2_decap_8 FILLER_91_672 ();
 sg13g2_decap_8 FILLER_91_679 ();
 sg13g2_decap_8 FILLER_91_686 ();
 sg13g2_decap_8 FILLER_91_693 ();
 sg13g2_decap_8 FILLER_91_700 ();
 sg13g2_decap_8 FILLER_91_707 ();
 sg13g2_decap_8 FILLER_91_714 ();
 sg13g2_decap_8 FILLER_91_721 ();
 sg13g2_decap_8 FILLER_91_728 ();
 sg13g2_decap_8 FILLER_91_735 ();
 sg13g2_decap_8 FILLER_91_742 ();
 sg13g2_decap_8 FILLER_91_749 ();
 sg13g2_decap_8 FILLER_91_756 ();
 sg13g2_decap_8 FILLER_91_763 ();
 sg13g2_decap_8 FILLER_91_770 ();
 sg13g2_decap_8 FILLER_91_777 ();
 sg13g2_decap_8 FILLER_91_784 ();
 sg13g2_decap_8 FILLER_91_791 ();
 sg13g2_decap_8 FILLER_91_798 ();
 sg13g2_decap_8 FILLER_91_805 ();
 sg13g2_decap_8 FILLER_91_812 ();
 sg13g2_decap_8 FILLER_91_819 ();
 sg13g2_decap_8 FILLER_91_826 ();
 sg13g2_decap_8 FILLER_91_833 ();
 sg13g2_fill_1 FILLER_91_840 ();
 sg13g2_decap_8 FILLER_92_0 ();
 sg13g2_decap_8 FILLER_92_7 ();
 sg13g2_decap_8 FILLER_92_14 ();
 sg13g2_decap_8 FILLER_92_21 ();
 sg13g2_decap_8 FILLER_92_28 ();
 sg13g2_decap_8 FILLER_92_35 ();
 sg13g2_decap_8 FILLER_92_42 ();
 sg13g2_decap_8 FILLER_92_49 ();
 sg13g2_decap_8 FILLER_92_56 ();
 sg13g2_decap_8 FILLER_92_63 ();
 sg13g2_decap_8 FILLER_92_70 ();
 sg13g2_decap_8 FILLER_92_77 ();
 sg13g2_decap_8 FILLER_92_84 ();
 sg13g2_decap_8 FILLER_92_91 ();
 sg13g2_decap_8 FILLER_92_98 ();
 sg13g2_decap_8 FILLER_92_105 ();
 sg13g2_decap_8 FILLER_92_112 ();
 sg13g2_decap_8 FILLER_92_119 ();
 sg13g2_decap_8 FILLER_92_126 ();
 sg13g2_decap_8 FILLER_92_133 ();
 sg13g2_decap_8 FILLER_92_140 ();
 sg13g2_decap_8 FILLER_92_147 ();
 sg13g2_decap_8 FILLER_92_154 ();
 sg13g2_decap_8 FILLER_92_161 ();
 sg13g2_decap_8 FILLER_92_168 ();
 sg13g2_decap_8 FILLER_92_175 ();
 sg13g2_decap_8 FILLER_92_182 ();
 sg13g2_decap_8 FILLER_92_189 ();
 sg13g2_decap_8 FILLER_92_196 ();
 sg13g2_decap_8 FILLER_92_203 ();
 sg13g2_decap_8 FILLER_92_210 ();
 sg13g2_decap_8 FILLER_92_217 ();
 sg13g2_decap_8 FILLER_92_224 ();
 sg13g2_decap_8 FILLER_92_231 ();
 sg13g2_decap_8 FILLER_92_238 ();
 sg13g2_decap_8 FILLER_92_245 ();
 sg13g2_decap_8 FILLER_92_252 ();
 sg13g2_decap_8 FILLER_92_259 ();
 sg13g2_decap_8 FILLER_92_266 ();
 sg13g2_decap_8 FILLER_92_273 ();
 sg13g2_decap_8 FILLER_92_280 ();
 sg13g2_decap_8 FILLER_92_287 ();
 sg13g2_decap_8 FILLER_92_294 ();
 sg13g2_decap_8 FILLER_92_301 ();
 sg13g2_decap_8 FILLER_92_308 ();
 sg13g2_decap_8 FILLER_92_315 ();
 sg13g2_decap_8 FILLER_92_322 ();
 sg13g2_decap_8 FILLER_92_329 ();
 sg13g2_decap_8 FILLER_92_336 ();
 sg13g2_decap_8 FILLER_92_343 ();
 sg13g2_decap_8 FILLER_92_350 ();
 sg13g2_decap_8 FILLER_92_357 ();
 sg13g2_decap_8 FILLER_92_364 ();
 sg13g2_decap_8 FILLER_92_371 ();
 sg13g2_decap_8 FILLER_92_378 ();
 sg13g2_decap_8 FILLER_92_385 ();
 sg13g2_decap_8 FILLER_92_392 ();
 sg13g2_decap_8 FILLER_92_399 ();
 sg13g2_decap_8 FILLER_92_406 ();
 sg13g2_decap_8 FILLER_92_413 ();
 sg13g2_decap_8 FILLER_92_420 ();
 sg13g2_decap_8 FILLER_92_427 ();
 sg13g2_decap_8 FILLER_92_434 ();
 sg13g2_decap_8 FILLER_92_441 ();
 sg13g2_decap_8 FILLER_92_448 ();
 sg13g2_decap_8 FILLER_92_455 ();
 sg13g2_decap_8 FILLER_92_462 ();
 sg13g2_decap_8 FILLER_92_469 ();
 sg13g2_decap_8 FILLER_92_476 ();
 sg13g2_decap_8 FILLER_92_483 ();
 sg13g2_decap_8 FILLER_92_490 ();
 sg13g2_decap_8 FILLER_92_497 ();
 sg13g2_decap_8 FILLER_92_504 ();
 sg13g2_decap_8 FILLER_92_511 ();
 sg13g2_decap_8 FILLER_92_518 ();
 sg13g2_decap_8 FILLER_92_525 ();
 sg13g2_decap_8 FILLER_92_532 ();
 sg13g2_decap_8 FILLER_92_539 ();
 sg13g2_decap_8 FILLER_92_546 ();
 sg13g2_decap_8 FILLER_92_553 ();
 sg13g2_decap_8 FILLER_92_560 ();
 sg13g2_decap_8 FILLER_92_567 ();
 sg13g2_decap_8 FILLER_92_574 ();
 sg13g2_decap_8 FILLER_92_581 ();
 sg13g2_decap_8 FILLER_92_588 ();
 sg13g2_decap_8 FILLER_92_595 ();
 sg13g2_decap_8 FILLER_92_602 ();
 sg13g2_decap_8 FILLER_92_609 ();
 sg13g2_decap_8 FILLER_92_616 ();
 sg13g2_decap_8 FILLER_92_623 ();
 sg13g2_decap_8 FILLER_92_630 ();
 sg13g2_decap_8 FILLER_92_637 ();
 sg13g2_decap_8 FILLER_92_644 ();
 sg13g2_decap_8 FILLER_92_651 ();
 sg13g2_decap_8 FILLER_92_658 ();
 sg13g2_decap_8 FILLER_92_665 ();
 sg13g2_decap_8 FILLER_92_672 ();
 sg13g2_decap_8 FILLER_92_679 ();
 sg13g2_decap_8 FILLER_92_686 ();
 sg13g2_decap_8 FILLER_92_693 ();
 sg13g2_decap_8 FILLER_92_700 ();
 sg13g2_decap_8 FILLER_92_707 ();
 sg13g2_decap_8 FILLER_92_714 ();
 sg13g2_decap_8 FILLER_92_721 ();
 sg13g2_decap_8 FILLER_92_728 ();
 sg13g2_decap_8 FILLER_92_735 ();
 sg13g2_decap_8 FILLER_92_742 ();
 sg13g2_decap_8 FILLER_92_749 ();
 sg13g2_decap_8 FILLER_92_756 ();
 sg13g2_decap_8 FILLER_92_763 ();
 sg13g2_decap_8 FILLER_92_770 ();
 sg13g2_decap_8 FILLER_92_777 ();
 sg13g2_decap_8 FILLER_92_784 ();
 sg13g2_decap_8 FILLER_92_791 ();
 sg13g2_decap_8 FILLER_92_798 ();
 sg13g2_decap_8 FILLER_92_805 ();
 sg13g2_decap_8 FILLER_92_812 ();
 sg13g2_decap_8 FILLER_92_819 ();
 sg13g2_decap_8 FILLER_92_826 ();
 sg13g2_decap_8 FILLER_92_833 ();
 sg13g2_fill_1 FILLER_92_840 ();
 sg13g2_decap_8 FILLER_93_0 ();
 sg13g2_decap_8 FILLER_93_7 ();
 sg13g2_decap_8 FILLER_93_14 ();
 sg13g2_decap_8 FILLER_93_21 ();
 sg13g2_decap_8 FILLER_93_28 ();
 sg13g2_decap_8 FILLER_93_35 ();
 sg13g2_decap_8 FILLER_93_42 ();
 sg13g2_decap_8 FILLER_93_49 ();
 sg13g2_decap_8 FILLER_93_56 ();
 sg13g2_decap_8 FILLER_93_63 ();
 sg13g2_decap_8 FILLER_93_70 ();
 sg13g2_decap_8 FILLER_93_77 ();
 sg13g2_decap_8 FILLER_93_84 ();
 sg13g2_decap_8 FILLER_93_91 ();
 sg13g2_decap_8 FILLER_93_98 ();
 sg13g2_decap_8 FILLER_93_105 ();
 sg13g2_decap_8 FILLER_93_112 ();
 sg13g2_decap_8 FILLER_93_119 ();
 sg13g2_decap_8 FILLER_93_126 ();
 sg13g2_decap_8 FILLER_93_133 ();
 sg13g2_decap_8 FILLER_93_140 ();
 sg13g2_decap_8 FILLER_93_147 ();
 sg13g2_decap_8 FILLER_93_154 ();
 sg13g2_decap_8 FILLER_93_161 ();
 sg13g2_decap_8 FILLER_93_168 ();
 sg13g2_decap_8 FILLER_93_175 ();
 sg13g2_decap_8 FILLER_93_182 ();
 sg13g2_decap_8 FILLER_93_189 ();
 sg13g2_decap_8 FILLER_93_196 ();
 sg13g2_decap_8 FILLER_93_203 ();
 sg13g2_decap_8 FILLER_93_210 ();
 sg13g2_decap_8 FILLER_93_217 ();
 sg13g2_decap_8 FILLER_93_224 ();
 sg13g2_decap_8 FILLER_93_231 ();
 sg13g2_decap_8 FILLER_93_238 ();
 sg13g2_decap_8 FILLER_93_245 ();
 sg13g2_decap_8 FILLER_93_252 ();
 sg13g2_decap_8 FILLER_93_259 ();
 sg13g2_decap_8 FILLER_93_266 ();
 sg13g2_decap_8 FILLER_93_273 ();
 sg13g2_decap_8 FILLER_93_280 ();
 sg13g2_decap_8 FILLER_93_287 ();
 sg13g2_decap_8 FILLER_93_294 ();
 sg13g2_decap_8 FILLER_93_301 ();
 sg13g2_decap_8 FILLER_93_308 ();
 sg13g2_decap_8 FILLER_93_315 ();
 sg13g2_decap_8 FILLER_93_322 ();
 sg13g2_decap_8 FILLER_93_329 ();
 sg13g2_decap_8 FILLER_93_336 ();
 sg13g2_decap_8 FILLER_93_343 ();
 sg13g2_decap_8 FILLER_93_350 ();
 sg13g2_decap_8 FILLER_93_357 ();
 sg13g2_decap_8 FILLER_93_364 ();
 sg13g2_decap_8 FILLER_93_371 ();
 sg13g2_decap_8 FILLER_93_378 ();
 sg13g2_decap_8 FILLER_93_385 ();
 sg13g2_decap_8 FILLER_93_392 ();
 sg13g2_decap_8 FILLER_93_399 ();
 sg13g2_decap_8 FILLER_93_406 ();
 sg13g2_decap_8 FILLER_93_413 ();
 sg13g2_decap_8 FILLER_93_420 ();
 sg13g2_decap_8 FILLER_93_427 ();
 sg13g2_decap_8 FILLER_93_434 ();
 sg13g2_decap_8 FILLER_93_441 ();
 sg13g2_decap_8 FILLER_93_448 ();
 sg13g2_decap_8 FILLER_93_455 ();
 sg13g2_decap_8 FILLER_93_462 ();
 sg13g2_decap_8 FILLER_93_469 ();
 sg13g2_decap_8 FILLER_93_476 ();
 sg13g2_decap_8 FILLER_93_483 ();
 sg13g2_decap_8 FILLER_93_490 ();
 sg13g2_decap_8 FILLER_93_497 ();
 sg13g2_decap_8 FILLER_93_504 ();
 sg13g2_decap_8 FILLER_93_511 ();
 sg13g2_decap_8 FILLER_93_518 ();
 sg13g2_decap_8 FILLER_93_525 ();
 sg13g2_decap_8 FILLER_93_532 ();
 sg13g2_decap_8 FILLER_93_539 ();
 sg13g2_decap_8 FILLER_93_546 ();
 sg13g2_decap_8 FILLER_93_553 ();
 sg13g2_decap_8 FILLER_93_560 ();
 sg13g2_decap_8 FILLER_93_567 ();
 sg13g2_decap_8 FILLER_93_574 ();
 sg13g2_decap_8 FILLER_93_581 ();
 sg13g2_decap_8 FILLER_93_588 ();
 sg13g2_decap_8 FILLER_93_595 ();
 sg13g2_decap_8 FILLER_93_602 ();
 sg13g2_decap_8 FILLER_93_609 ();
 sg13g2_decap_8 FILLER_93_616 ();
 sg13g2_decap_8 FILLER_93_623 ();
 sg13g2_decap_8 FILLER_93_630 ();
 sg13g2_decap_8 FILLER_93_637 ();
 sg13g2_decap_8 FILLER_93_644 ();
 sg13g2_decap_8 FILLER_93_651 ();
 sg13g2_decap_8 FILLER_93_658 ();
 sg13g2_decap_8 FILLER_93_665 ();
 sg13g2_decap_8 FILLER_93_672 ();
 sg13g2_decap_8 FILLER_93_679 ();
 sg13g2_decap_8 FILLER_93_686 ();
 sg13g2_decap_8 FILLER_93_693 ();
 sg13g2_decap_8 FILLER_93_700 ();
 sg13g2_decap_8 FILLER_93_707 ();
 sg13g2_decap_8 FILLER_93_714 ();
 sg13g2_decap_8 FILLER_93_721 ();
 sg13g2_decap_8 FILLER_93_728 ();
 sg13g2_decap_8 FILLER_93_735 ();
 sg13g2_decap_8 FILLER_93_742 ();
 sg13g2_decap_8 FILLER_93_749 ();
 sg13g2_decap_8 FILLER_93_756 ();
 sg13g2_decap_8 FILLER_93_763 ();
 sg13g2_decap_8 FILLER_93_770 ();
 sg13g2_decap_8 FILLER_93_777 ();
 sg13g2_decap_8 FILLER_93_784 ();
 sg13g2_decap_8 FILLER_93_791 ();
 sg13g2_decap_8 FILLER_93_798 ();
 sg13g2_decap_8 FILLER_93_805 ();
 sg13g2_decap_8 FILLER_93_812 ();
 sg13g2_decap_8 FILLER_93_819 ();
 sg13g2_decap_8 FILLER_93_826 ();
 sg13g2_decap_8 FILLER_93_833 ();
 sg13g2_fill_1 FILLER_93_840 ();
 sg13g2_decap_8 FILLER_94_0 ();
 sg13g2_decap_8 FILLER_94_7 ();
 sg13g2_decap_8 FILLER_94_14 ();
 sg13g2_decap_8 FILLER_94_21 ();
 sg13g2_decap_8 FILLER_94_28 ();
 sg13g2_decap_8 FILLER_94_35 ();
 sg13g2_decap_8 FILLER_94_42 ();
 sg13g2_decap_8 FILLER_94_49 ();
 sg13g2_decap_8 FILLER_94_56 ();
 sg13g2_decap_8 FILLER_94_63 ();
 sg13g2_decap_8 FILLER_94_70 ();
 sg13g2_decap_8 FILLER_94_77 ();
 sg13g2_decap_8 FILLER_94_84 ();
 sg13g2_decap_8 FILLER_94_91 ();
 sg13g2_decap_8 FILLER_94_98 ();
 sg13g2_decap_8 FILLER_94_105 ();
 sg13g2_decap_8 FILLER_94_112 ();
 sg13g2_decap_8 FILLER_94_119 ();
 sg13g2_decap_8 FILLER_94_126 ();
 sg13g2_decap_8 FILLER_94_133 ();
 sg13g2_decap_8 FILLER_94_140 ();
 sg13g2_decap_8 FILLER_94_147 ();
 sg13g2_decap_8 FILLER_94_154 ();
 sg13g2_decap_8 FILLER_94_161 ();
 sg13g2_decap_8 FILLER_94_168 ();
 sg13g2_decap_8 FILLER_94_175 ();
 sg13g2_decap_8 FILLER_94_182 ();
 sg13g2_decap_8 FILLER_94_189 ();
 sg13g2_decap_8 FILLER_94_196 ();
 sg13g2_decap_8 FILLER_94_203 ();
 sg13g2_decap_8 FILLER_94_210 ();
 sg13g2_decap_8 FILLER_94_217 ();
 sg13g2_decap_8 FILLER_94_224 ();
 sg13g2_decap_8 FILLER_94_231 ();
 sg13g2_decap_8 FILLER_94_238 ();
 sg13g2_decap_8 FILLER_94_245 ();
 sg13g2_decap_8 FILLER_94_252 ();
 sg13g2_decap_8 FILLER_94_259 ();
 sg13g2_decap_8 FILLER_94_266 ();
 sg13g2_decap_8 FILLER_94_273 ();
 sg13g2_decap_8 FILLER_94_280 ();
 sg13g2_decap_8 FILLER_94_287 ();
 sg13g2_decap_8 FILLER_94_294 ();
 sg13g2_decap_8 FILLER_94_301 ();
 sg13g2_decap_8 FILLER_94_308 ();
 sg13g2_decap_8 FILLER_94_315 ();
 sg13g2_decap_8 FILLER_94_322 ();
 sg13g2_decap_8 FILLER_94_329 ();
 sg13g2_decap_8 FILLER_94_336 ();
 sg13g2_decap_8 FILLER_94_343 ();
 sg13g2_decap_8 FILLER_94_350 ();
 sg13g2_decap_8 FILLER_94_357 ();
 sg13g2_decap_8 FILLER_94_364 ();
 sg13g2_decap_8 FILLER_94_371 ();
 sg13g2_decap_8 FILLER_94_378 ();
 sg13g2_decap_8 FILLER_94_385 ();
 sg13g2_decap_8 FILLER_94_392 ();
 sg13g2_decap_8 FILLER_94_399 ();
 sg13g2_decap_8 FILLER_94_406 ();
 sg13g2_decap_8 FILLER_94_413 ();
 sg13g2_decap_8 FILLER_94_420 ();
 sg13g2_decap_8 FILLER_94_427 ();
 sg13g2_decap_8 FILLER_94_434 ();
 sg13g2_decap_8 FILLER_94_441 ();
 sg13g2_decap_8 FILLER_94_448 ();
 sg13g2_decap_8 FILLER_94_455 ();
 sg13g2_decap_8 FILLER_94_462 ();
 sg13g2_decap_8 FILLER_94_469 ();
 sg13g2_decap_8 FILLER_94_476 ();
 sg13g2_decap_8 FILLER_94_483 ();
 sg13g2_decap_8 FILLER_94_490 ();
 sg13g2_decap_8 FILLER_94_497 ();
 sg13g2_decap_8 FILLER_94_504 ();
 sg13g2_decap_8 FILLER_94_511 ();
 sg13g2_decap_8 FILLER_94_518 ();
 sg13g2_decap_8 FILLER_94_525 ();
 sg13g2_decap_8 FILLER_94_532 ();
 sg13g2_decap_8 FILLER_94_539 ();
 sg13g2_decap_8 FILLER_94_546 ();
 sg13g2_decap_8 FILLER_94_553 ();
 sg13g2_decap_8 FILLER_94_560 ();
 sg13g2_decap_8 FILLER_94_567 ();
 sg13g2_decap_8 FILLER_94_574 ();
 sg13g2_decap_8 FILLER_94_581 ();
 sg13g2_decap_8 FILLER_94_588 ();
 sg13g2_decap_8 FILLER_94_595 ();
 sg13g2_decap_8 FILLER_94_602 ();
 sg13g2_decap_8 FILLER_94_609 ();
 sg13g2_decap_8 FILLER_94_616 ();
 sg13g2_decap_8 FILLER_94_623 ();
 sg13g2_decap_8 FILLER_94_630 ();
 sg13g2_decap_8 FILLER_94_637 ();
 sg13g2_decap_8 FILLER_94_644 ();
 sg13g2_decap_8 FILLER_94_651 ();
 sg13g2_decap_8 FILLER_94_658 ();
 sg13g2_decap_8 FILLER_94_665 ();
 sg13g2_decap_8 FILLER_94_672 ();
 sg13g2_decap_8 FILLER_94_679 ();
 sg13g2_decap_8 FILLER_94_686 ();
 sg13g2_decap_8 FILLER_94_693 ();
 sg13g2_decap_8 FILLER_94_700 ();
 sg13g2_decap_8 FILLER_94_707 ();
 sg13g2_decap_8 FILLER_94_714 ();
 sg13g2_decap_8 FILLER_94_721 ();
 sg13g2_decap_8 FILLER_94_728 ();
 sg13g2_decap_8 FILLER_94_735 ();
 sg13g2_decap_8 FILLER_94_742 ();
 sg13g2_decap_8 FILLER_94_749 ();
 sg13g2_decap_8 FILLER_94_756 ();
 sg13g2_decap_8 FILLER_94_763 ();
 sg13g2_decap_8 FILLER_94_770 ();
 sg13g2_decap_8 FILLER_94_777 ();
 sg13g2_decap_8 FILLER_94_784 ();
 sg13g2_decap_8 FILLER_94_791 ();
 sg13g2_decap_8 FILLER_94_798 ();
 sg13g2_decap_8 FILLER_94_805 ();
 sg13g2_decap_8 FILLER_94_812 ();
 sg13g2_decap_8 FILLER_94_819 ();
 sg13g2_decap_8 FILLER_94_826 ();
 sg13g2_decap_8 FILLER_94_833 ();
 sg13g2_fill_1 FILLER_94_840 ();
 sg13g2_decap_8 FILLER_95_0 ();
 sg13g2_decap_8 FILLER_95_7 ();
 sg13g2_decap_8 FILLER_95_14 ();
 sg13g2_decap_8 FILLER_95_21 ();
 sg13g2_decap_8 FILLER_95_28 ();
 sg13g2_decap_8 FILLER_95_35 ();
 sg13g2_decap_8 FILLER_95_42 ();
 sg13g2_decap_8 FILLER_95_49 ();
 sg13g2_decap_8 FILLER_95_56 ();
 sg13g2_decap_8 FILLER_95_63 ();
 sg13g2_decap_8 FILLER_95_70 ();
 sg13g2_decap_8 FILLER_95_77 ();
 sg13g2_decap_8 FILLER_95_84 ();
 sg13g2_decap_8 FILLER_95_91 ();
 sg13g2_decap_8 FILLER_95_98 ();
 sg13g2_decap_8 FILLER_95_105 ();
 sg13g2_decap_8 FILLER_95_112 ();
 sg13g2_decap_8 FILLER_95_119 ();
 sg13g2_decap_8 FILLER_95_126 ();
 sg13g2_decap_8 FILLER_95_133 ();
 sg13g2_decap_8 FILLER_95_140 ();
 sg13g2_decap_8 FILLER_95_147 ();
 sg13g2_decap_8 FILLER_95_154 ();
 sg13g2_decap_8 FILLER_95_161 ();
 sg13g2_decap_8 FILLER_95_168 ();
 sg13g2_decap_8 FILLER_95_175 ();
 sg13g2_decap_8 FILLER_95_182 ();
 sg13g2_decap_8 FILLER_95_189 ();
 sg13g2_decap_8 FILLER_95_196 ();
 sg13g2_decap_8 FILLER_95_203 ();
 sg13g2_decap_8 FILLER_95_210 ();
 sg13g2_decap_8 FILLER_95_217 ();
 sg13g2_decap_8 FILLER_95_224 ();
 sg13g2_decap_8 FILLER_95_231 ();
 sg13g2_decap_8 FILLER_95_238 ();
 sg13g2_decap_8 FILLER_95_245 ();
 sg13g2_decap_8 FILLER_95_252 ();
 sg13g2_decap_8 FILLER_95_259 ();
 sg13g2_decap_8 FILLER_95_266 ();
 sg13g2_decap_8 FILLER_95_273 ();
 sg13g2_decap_8 FILLER_95_280 ();
 sg13g2_decap_8 FILLER_95_287 ();
 sg13g2_decap_8 FILLER_95_294 ();
 sg13g2_decap_8 FILLER_95_301 ();
 sg13g2_decap_8 FILLER_95_308 ();
 sg13g2_decap_8 FILLER_95_315 ();
 sg13g2_decap_8 FILLER_95_322 ();
 sg13g2_decap_8 FILLER_95_329 ();
 sg13g2_decap_8 FILLER_95_336 ();
 sg13g2_decap_8 FILLER_95_343 ();
 sg13g2_decap_8 FILLER_95_350 ();
 sg13g2_decap_8 FILLER_95_357 ();
 sg13g2_decap_8 FILLER_95_364 ();
 sg13g2_decap_8 FILLER_95_371 ();
 sg13g2_decap_8 FILLER_95_378 ();
 sg13g2_decap_8 FILLER_95_385 ();
 sg13g2_decap_8 FILLER_95_392 ();
 sg13g2_decap_8 FILLER_95_399 ();
 sg13g2_decap_8 FILLER_95_406 ();
 sg13g2_decap_8 FILLER_95_413 ();
 sg13g2_decap_8 FILLER_95_420 ();
 sg13g2_decap_8 FILLER_95_427 ();
 sg13g2_decap_8 FILLER_95_434 ();
 sg13g2_decap_8 FILLER_95_441 ();
 sg13g2_decap_8 FILLER_95_448 ();
 sg13g2_decap_8 FILLER_95_455 ();
 sg13g2_decap_8 FILLER_95_462 ();
 sg13g2_decap_8 FILLER_95_469 ();
 sg13g2_decap_8 FILLER_95_476 ();
 sg13g2_decap_8 FILLER_95_483 ();
 sg13g2_decap_8 FILLER_95_490 ();
 sg13g2_decap_8 FILLER_95_497 ();
 sg13g2_decap_8 FILLER_95_504 ();
 sg13g2_decap_8 FILLER_95_511 ();
 sg13g2_decap_8 FILLER_95_518 ();
 sg13g2_decap_8 FILLER_95_525 ();
 sg13g2_decap_8 FILLER_95_532 ();
 sg13g2_decap_8 FILLER_95_539 ();
 sg13g2_decap_8 FILLER_95_546 ();
 sg13g2_decap_8 FILLER_95_553 ();
 sg13g2_decap_8 FILLER_95_560 ();
 sg13g2_decap_8 FILLER_95_567 ();
 sg13g2_decap_8 FILLER_95_574 ();
 sg13g2_decap_8 FILLER_95_581 ();
 sg13g2_decap_8 FILLER_95_588 ();
 sg13g2_decap_8 FILLER_95_595 ();
 sg13g2_decap_8 FILLER_95_602 ();
 sg13g2_decap_8 FILLER_95_609 ();
 sg13g2_decap_8 FILLER_95_616 ();
 sg13g2_decap_8 FILLER_95_623 ();
 sg13g2_decap_8 FILLER_95_630 ();
 sg13g2_decap_8 FILLER_95_637 ();
 sg13g2_decap_8 FILLER_95_644 ();
 sg13g2_decap_8 FILLER_95_651 ();
 sg13g2_decap_8 FILLER_95_658 ();
 sg13g2_decap_8 FILLER_95_665 ();
 sg13g2_decap_8 FILLER_95_672 ();
 sg13g2_decap_8 FILLER_95_679 ();
 sg13g2_decap_8 FILLER_95_686 ();
 sg13g2_decap_8 FILLER_95_693 ();
 sg13g2_decap_8 FILLER_95_700 ();
 sg13g2_decap_8 FILLER_95_707 ();
 sg13g2_decap_8 FILLER_95_714 ();
 sg13g2_decap_8 FILLER_95_721 ();
 sg13g2_decap_8 FILLER_95_728 ();
 sg13g2_decap_8 FILLER_95_735 ();
 sg13g2_decap_8 FILLER_95_742 ();
 sg13g2_decap_8 FILLER_95_749 ();
 sg13g2_decap_8 FILLER_95_756 ();
 sg13g2_decap_8 FILLER_95_763 ();
 sg13g2_decap_8 FILLER_95_770 ();
 sg13g2_decap_8 FILLER_95_777 ();
 sg13g2_decap_8 FILLER_95_784 ();
 sg13g2_decap_8 FILLER_95_791 ();
 sg13g2_decap_8 FILLER_95_798 ();
 sg13g2_decap_8 FILLER_95_805 ();
 sg13g2_decap_8 FILLER_95_812 ();
 sg13g2_decap_8 FILLER_95_819 ();
 sg13g2_decap_8 FILLER_95_826 ();
 sg13g2_decap_8 FILLER_95_833 ();
 sg13g2_fill_1 FILLER_95_840 ();
 sg13g2_decap_8 FILLER_96_0 ();
 sg13g2_decap_8 FILLER_96_7 ();
 sg13g2_decap_8 FILLER_96_14 ();
 sg13g2_decap_8 FILLER_96_21 ();
 sg13g2_decap_8 FILLER_96_28 ();
 sg13g2_decap_8 FILLER_96_35 ();
 sg13g2_decap_8 FILLER_96_42 ();
 sg13g2_decap_8 FILLER_96_49 ();
 sg13g2_decap_8 FILLER_96_56 ();
 sg13g2_decap_8 FILLER_96_63 ();
 sg13g2_decap_8 FILLER_96_70 ();
 sg13g2_decap_8 FILLER_96_77 ();
 sg13g2_decap_8 FILLER_96_84 ();
 sg13g2_decap_8 FILLER_96_91 ();
 sg13g2_decap_8 FILLER_96_98 ();
 sg13g2_decap_8 FILLER_96_105 ();
 sg13g2_decap_8 FILLER_96_112 ();
 sg13g2_decap_8 FILLER_96_119 ();
 sg13g2_decap_8 FILLER_96_126 ();
 sg13g2_decap_8 FILLER_96_133 ();
 sg13g2_decap_8 FILLER_96_140 ();
 sg13g2_decap_8 FILLER_96_147 ();
 sg13g2_decap_8 FILLER_96_154 ();
 sg13g2_decap_8 FILLER_96_161 ();
 sg13g2_decap_8 FILLER_96_168 ();
 sg13g2_decap_8 FILLER_96_175 ();
 sg13g2_decap_8 FILLER_96_182 ();
 sg13g2_decap_8 FILLER_96_189 ();
 sg13g2_decap_8 FILLER_96_196 ();
 sg13g2_decap_8 FILLER_96_203 ();
 sg13g2_decap_8 FILLER_96_210 ();
 sg13g2_decap_8 FILLER_96_217 ();
 sg13g2_decap_8 FILLER_96_224 ();
 sg13g2_decap_8 FILLER_96_231 ();
 sg13g2_decap_8 FILLER_96_238 ();
 sg13g2_decap_8 FILLER_96_245 ();
 sg13g2_decap_8 FILLER_96_252 ();
 sg13g2_decap_8 FILLER_96_259 ();
 sg13g2_decap_8 FILLER_96_266 ();
 sg13g2_decap_8 FILLER_96_273 ();
 sg13g2_decap_8 FILLER_96_280 ();
 sg13g2_decap_8 FILLER_96_287 ();
 sg13g2_decap_8 FILLER_96_294 ();
 sg13g2_decap_8 FILLER_96_301 ();
 sg13g2_decap_8 FILLER_96_308 ();
 sg13g2_decap_8 FILLER_96_315 ();
 sg13g2_decap_8 FILLER_96_322 ();
 sg13g2_decap_8 FILLER_96_329 ();
 sg13g2_decap_8 FILLER_96_336 ();
 sg13g2_decap_8 FILLER_96_343 ();
 sg13g2_decap_8 FILLER_96_350 ();
 sg13g2_decap_8 FILLER_96_357 ();
 sg13g2_decap_8 FILLER_96_364 ();
 sg13g2_decap_8 FILLER_96_371 ();
 sg13g2_decap_8 FILLER_96_378 ();
 sg13g2_decap_8 FILLER_96_385 ();
 sg13g2_decap_8 FILLER_96_392 ();
 sg13g2_decap_8 FILLER_96_399 ();
 sg13g2_decap_8 FILLER_96_406 ();
 sg13g2_decap_8 FILLER_96_413 ();
 sg13g2_decap_8 FILLER_96_420 ();
 sg13g2_decap_8 FILLER_96_427 ();
 sg13g2_decap_8 FILLER_96_434 ();
 sg13g2_decap_8 FILLER_96_441 ();
 sg13g2_decap_8 FILLER_96_448 ();
 sg13g2_decap_8 FILLER_96_455 ();
 sg13g2_decap_8 FILLER_96_462 ();
 sg13g2_decap_8 FILLER_96_469 ();
 sg13g2_decap_8 FILLER_96_476 ();
 sg13g2_decap_8 FILLER_96_483 ();
 sg13g2_decap_8 FILLER_96_490 ();
 sg13g2_decap_8 FILLER_96_497 ();
 sg13g2_decap_8 FILLER_96_504 ();
 sg13g2_decap_8 FILLER_96_511 ();
 sg13g2_decap_8 FILLER_96_518 ();
 sg13g2_decap_8 FILLER_96_525 ();
 sg13g2_decap_8 FILLER_96_532 ();
 sg13g2_decap_8 FILLER_96_539 ();
 sg13g2_decap_8 FILLER_96_546 ();
 sg13g2_decap_8 FILLER_96_553 ();
 sg13g2_decap_8 FILLER_96_560 ();
 sg13g2_decap_8 FILLER_96_567 ();
 sg13g2_decap_8 FILLER_96_574 ();
 sg13g2_decap_8 FILLER_96_581 ();
 sg13g2_decap_8 FILLER_96_588 ();
 sg13g2_decap_8 FILLER_96_595 ();
 sg13g2_decap_8 FILLER_96_602 ();
 sg13g2_decap_8 FILLER_96_609 ();
 sg13g2_decap_8 FILLER_96_616 ();
 sg13g2_decap_8 FILLER_96_623 ();
 sg13g2_decap_8 FILLER_96_630 ();
 sg13g2_decap_8 FILLER_96_637 ();
 sg13g2_decap_8 FILLER_96_644 ();
 sg13g2_decap_8 FILLER_96_651 ();
 sg13g2_decap_8 FILLER_96_658 ();
 sg13g2_decap_8 FILLER_96_665 ();
 sg13g2_decap_8 FILLER_96_672 ();
 sg13g2_decap_8 FILLER_96_679 ();
 sg13g2_decap_8 FILLER_96_686 ();
 sg13g2_decap_8 FILLER_96_693 ();
 sg13g2_decap_8 FILLER_96_700 ();
 sg13g2_decap_8 FILLER_96_707 ();
 sg13g2_decap_8 FILLER_96_714 ();
 sg13g2_decap_8 FILLER_96_721 ();
 sg13g2_decap_8 FILLER_96_728 ();
 sg13g2_decap_8 FILLER_96_735 ();
 sg13g2_decap_8 FILLER_96_742 ();
 sg13g2_decap_8 FILLER_96_749 ();
 sg13g2_decap_8 FILLER_96_756 ();
 sg13g2_decap_8 FILLER_96_763 ();
 sg13g2_decap_8 FILLER_96_770 ();
 sg13g2_decap_8 FILLER_96_777 ();
 sg13g2_decap_8 FILLER_96_784 ();
 sg13g2_decap_8 FILLER_96_791 ();
 sg13g2_decap_8 FILLER_96_798 ();
 sg13g2_decap_8 FILLER_96_805 ();
 sg13g2_decap_8 FILLER_96_812 ();
 sg13g2_decap_8 FILLER_96_819 ();
 sg13g2_decap_8 FILLER_96_826 ();
 sg13g2_decap_8 FILLER_96_833 ();
 sg13g2_fill_1 FILLER_96_840 ();
 sg13g2_decap_8 FILLER_97_0 ();
 sg13g2_decap_8 FILLER_97_7 ();
 sg13g2_decap_8 FILLER_97_14 ();
 sg13g2_decap_8 FILLER_97_21 ();
 sg13g2_decap_8 FILLER_97_28 ();
 sg13g2_decap_8 FILLER_97_35 ();
 sg13g2_decap_8 FILLER_97_42 ();
 sg13g2_decap_8 FILLER_97_49 ();
 sg13g2_decap_8 FILLER_97_56 ();
 sg13g2_decap_8 FILLER_97_63 ();
 sg13g2_decap_8 FILLER_97_70 ();
 sg13g2_decap_8 FILLER_97_77 ();
 sg13g2_decap_8 FILLER_97_84 ();
 sg13g2_decap_8 FILLER_97_91 ();
 sg13g2_decap_8 FILLER_97_98 ();
 sg13g2_decap_8 FILLER_97_105 ();
 sg13g2_decap_8 FILLER_97_112 ();
 sg13g2_decap_8 FILLER_97_119 ();
 sg13g2_decap_8 FILLER_97_126 ();
 sg13g2_decap_8 FILLER_97_133 ();
 sg13g2_decap_8 FILLER_97_140 ();
 sg13g2_decap_8 FILLER_97_147 ();
 sg13g2_decap_8 FILLER_97_154 ();
 sg13g2_decap_8 FILLER_97_161 ();
 sg13g2_decap_8 FILLER_97_168 ();
 sg13g2_decap_8 FILLER_97_175 ();
 sg13g2_decap_8 FILLER_97_182 ();
 sg13g2_decap_8 FILLER_97_189 ();
 sg13g2_decap_8 FILLER_97_196 ();
 sg13g2_decap_8 FILLER_97_203 ();
 sg13g2_decap_8 FILLER_97_210 ();
 sg13g2_decap_8 FILLER_97_217 ();
 sg13g2_decap_8 FILLER_97_224 ();
 sg13g2_decap_8 FILLER_97_231 ();
 sg13g2_decap_8 FILLER_97_238 ();
 sg13g2_decap_8 FILLER_97_245 ();
 sg13g2_decap_8 FILLER_97_252 ();
 sg13g2_decap_8 FILLER_97_259 ();
 sg13g2_decap_8 FILLER_97_266 ();
 sg13g2_decap_8 FILLER_97_273 ();
 sg13g2_decap_8 FILLER_97_280 ();
 sg13g2_decap_8 FILLER_97_287 ();
 sg13g2_decap_8 FILLER_97_294 ();
 sg13g2_decap_8 FILLER_97_301 ();
 sg13g2_decap_8 FILLER_97_308 ();
 sg13g2_decap_8 FILLER_97_315 ();
 sg13g2_decap_8 FILLER_97_322 ();
 sg13g2_decap_8 FILLER_97_329 ();
 sg13g2_decap_8 FILLER_97_336 ();
 sg13g2_decap_8 FILLER_97_343 ();
 sg13g2_decap_8 FILLER_97_350 ();
 sg13g2_decap_8 FILLER_97_357 ();
 sg13g2_decap_8 FILLER_97_364 ();
 sg13g2_decap_8 FILLER_97_371 ();
 sg13g2_decap_8 FILLER_97_378 ();
 sg13g2_decap_8 FILLER_97_385 ();
 sg13g2_decap_8 FILLER_97_392 ();
 sg13g2_decap_8 FILLER_97_399 ();
 sg13g2_decap_8 FILLER_97_406 ();
 sg13g2_decap_8 FILLER_97_413 ();
 sg13g2_decap_8 FILLER_97_420 ();
 sg13g2_decap_8 FILLER_97_427 ();
 sg13g2_decap_8 FILLER_97_434 ();
 sg13g2_decap_8 FILLER_97_441 ();
 sg13g2_decap_8 FILLER_97_448 ();
 sg13g2_decap_8 FILLER_97_455 ();
 sg13g2_decap_8 FILLER_97_462 ();
 sg13g2_decap_8 FILLER_97_469 ();
 sg13g2_decap_8 FILLER_97_476 ();
 sg13g2_decap_8 FILLER_97_483 ();
 sg13g2_decap_8 FILLER_97_490 ();
 sg13g2_decap_8 FILLER_97_497 ();
 sg13g2_decap_8 FILLER_97_504 ();
 sg13g2_decap_8 FILLER_97_511 ();
 sg13g2_decap_8 FILLER_97_518 ();
 sg13g2_decap_8 FILLER_97_525 ();
 sg13g2_decap_8 FILLER_97_532 ();
 sg13g2_decap_8 FILLER_97_539 ();
 sg13g2_decap_8 FILLER_97_546 ();
 sg13g2_decap_8 FILLER_97_553 ();
 sg13g2_decap_8 FILLER_97_560 ();
 sg13g2_decap_8 FILLER_97_567 ();
 sg13g2_decap_8 FILLER_97_574 ();
 sg13g2_decap_8 FILLER_97_581 ();
 sg13g2_decap_8 FILLER_97_588 ();
 sg13g2_decap_8 FILLER_97_595 ();
 sg13g2_decap_8 FILLER_97_602 ();
 sg13g2_decap_8 FILLER_97_609 ();
 sg13g2_decap_8 FILLER_97_616 ();
 sg13g2_decap_8 FILLER_97_623 ();
 sg13g2_decap_8 FILLER_97_630 ();
 sg13g2_decap_8 FILLER_97_637 ();
 sg13g2_decap_8 FILLER_97_644 ();
 sg13g2_decap_8 FILLER_97_651 ();
 sg13g2_decap_8 FILLER_97_658 ();
 sg13g2_decap_8 FILLER_97_665 ();
 sg13g2_decap_8 FILLER_97_672 ();
 sg13g2_decap_8 FILLER_97_679 ();
 sg13g2_decap_8 FILLER_97_686 ();
 sg13g2_decap_8 FILLER_97_693 ();
 sg13g2_decap_8 FILLER_97_700 ();
 sg13g2_decap_8 FILLER_97_707 ();
 sg13g2_decap_8 FILLER_97_714 ();
 sg13g2_decap_8 FILLER_97_721 ();
 sg13g2_decap_8 FILLER_97_728 ();
 sg13g2_decap_8 FILLER_97_735 ();
 sg13g2_decap_8 FILLER_97_742 ();
 sg13g2_decap_8 FILLER_97_749 ();
 sg13g2_decap_8 FILLER_97_756 ();
 sg13g2_decap_8 FILLER_97_763 ();
 sg13g2_decap_8 FILLER_97_770 ();
 sg13g2_decap_8 FILLER_97_777 ();
 sg13g2_decap_8 FILLER_97_784 ();
 sg13g2_decap_8 FILLER_97_791 ();
 sg13g2_decap_8 FILLER_97_798 ();
 sg13g2_decap_8 FILLER_97_805 ();
 sg13g2_decap_8 FILLER_97_812 ();
 sg13g2_decap_8 FILLER_97_819 ();
 sg13g2_decap_8 FILLER_97_826 ();
 sg13g2_decap_8 FILLER_97_833 ();
 sg13g2_fill_1 FILLER_97_840 ();
 sg13g2_decap_8 FILLER_98_0 ();
 sg13g2_decap_8 FILLER_98_7 ();
 sg13g2_decap_8 FILLER_98_14 ();
 sg13g2_decap_8 FILLER_98_21 ();
 sg13g2_decap_8 FILLER_98_28 ();
 sg13g2_decap_8 FILLER_98_35 ();
 sg13g2_decap_8 FILLER_98_42 ();
 sg13g2_decap_8 FILLER_98_49 ();
 sg13g2_decap_8 FILLER_98_56 ();
 sg13g2_decap_8 FILLER_98_63 ();
 sg13g2_decap_8 FILLER_98_70 ();
 sg13g2_decap_8 FILLER_98_77 ();
 sg13g2_decap_8 FILLER_98_84 ();
 sg13g2_decap_8 FILLER_98_91 ();
 sg13g2_decap_8 FILLER_98_98 ();
 sg13g2_decap_8 FILLER_98_105 ();
 sg13g2_decap_8 FILLER_98_112 ();
 sg13g2_decap_8 FILLER_98_119 ();
 sg13g2_decap_8 FILLER_98_126 ();
 sg13g2_decap_8 FILLER_98_133 ();
 sg13g2_decap_8 FILLER_98_140 ();
 sg13g2_decap_8 FILLER_98_147 ();
 sg13g2_decap_8 FILLER_98_154 ();
 sg13g2_decap_8 FILLER_98_161 ();
 sg13g2_decap_8 FILLER_98_168 ();
 sg13g2_decap_8 FILLER_98_175 ();
 sg13g2_decap_8 FILLER_98_182 ();
 sg13g2_decap_8 FILLER_98_189 ();
 sg13g2_decap_8 FILLER_98_196 ();
 sg13g2_decap_8 FILLER_98_203 ();
 sg13g2_decap_8 FILLER_98_210 ();
 sg13g2_decap_8 FILLER_98_217 ();
 sg13g2_decap_8 FILLER_98_224 ();
 sg13g2_decap_8 FILLER_98_231 ();
 sg13g2_decap_8 FILLER_98_238 ();
 sg13g2_decap_8 FILLER_98_245 ();
 sg13g2_decap_8 FILLER_98_252 ();
 sg13g2_decap_8 FILLER_98_259 ();
 sg13g2_decap_8 FILLER_98_266 ();
 sg13g2_decap_8 FILLER_98_273 ();
 sg13g2_decap_8 FILLER_98_280 ();
 sg13g2_decap_8 FILLER_98_287 ();
 sg13g2_decap_8 FILLER_98_294 ();
 sg13g2_decap_8 FILLER_98_301 ();
 sg13g2_decap_8 FILLER_98_308 ();
 sg13g2_decap_8 FILLER_98_315 ();
 sg13g2_decap_8 FILLER_98_322 ();
 sg13g2_decap_8 FILLER_98_329 ();
 sg13g2_decap_8 FILLER_98_336 ();
 sg13g2_decap_8 FILLER_98_343 ();
 sg13g2_decap_8 FILLER_98_350 ();
 sg13g2_decap_8 FILLER_98_357 ();
 sg13g2_decap_8 FILLER_98_364 ();
 sg13g2_decap_8 FILLER_98_371 ();
 sg13g2_decap_8 FILLER_98_378 ();
 sg13g2_decap_8 FILLER_98_385 ();
 sg13g2_decap_8 FILLER_98_392 ();
 sg13g2_decap_8 FILLER_98_399 ();
 sg13g2_decap_8 FILLER_98_406 ();
 sg13g2_decap_8 FILLER_98_413 ();
 sg13g2_decap_8 FILLER_98_420 ();
 sg13g2_decap_8 FILLER_98_427 ();
 sg13g2_decap_8 FILLER_98_434 ();
 sg13g2_decap_8 FILLER_98_441 ();
 sg13g2_decap_8 FILLER_98_448 ();
 sg13g2_decap_8 FILLER_98_455 ();
 sg13g2_decap_8 FILLER_98_462 ();
 sg13g2_decap_8 FILLER_98_469 ();
 sg13g2_decap_8 FILLER_98_476 ();
 sg13g2_decap_8 FILLER_98_483 ();
 sg13g2_decap_8 FILLER_98_490 ();
 sg13g2_decap_8 FILLER_98_497 ();
 sg13g2_decap_8 FILLER_98_504 ();
 sg13g2_decap_8 FILLER_98_511 ();
 sg13g2_decap_8 FILLER_98_518 ();
 sg13g2_decap_8 FILLER_98_525 ();
 sg13g2_decap_8 FILLER_98_532 ();
 sg13g2_decap_8 FILLER_98_539 ();
 sg13g2_decap_8 FILLER_98_546 ();
 sg13g2_decap_8 FILLER_98_553 ();
 sg13g2_decap_8 FILLER_98_560 ();
 sg13g2_decap_8 FILLER_98_567 ();
 sg13g2_decap_8 FILLER_98_574 ();
 sg13g2_decap_8 FILLER_98_581 ();
 sg13g2_decap_8 FILLER_98_588 ();
 sg13g2_decap_8 FILLER_98_595 ();
 sg13g2_decap_8 FILLER_98_602 ();
 sg13g2_decap_8 FILLER_98_609 ();
 sg13g2_decap_8 FILLER_98_616 ();
 sg13g2_decap_8 FILLER_98_623 ();
 sg13g2_decap_8 FILLER_98_630 ();
 sg13g2_decap_8 FILLER_98_637 ();
 sg13g2_decap_8 FILLER_98_644 ();
 sg13g2_decap_8 FILLER_98_651 ();
 sg13g2_decap_8 FILLER_98_658 ();
 sg13g2_decap_8 FILLER_98_665 ();
 sg13g2_decap_8 FILLER_98_672 ();
 sg13g2_decap_8 FILLER_98_679 ();
 sg13g2_decap_8 FILLER_98_686 ();
 sg13g2_decap_8 FILLER_98_693 ();
 sg13g2_decap_8 FILLER_98_700 ();
 sg13g2_decap_8 FILLER_98_707 ();
 sg13g2_decap_8 FILLER_98_714 ();
 sg13g2_decap_8 FILLER_98_721 ();
 sg13g2_decap_8 FILLER_98_728 ();
 sg13g2_decap_8 FILLER_98_735 ();
 sg13g2_decap_8 FILLER_98_742 ();
 sg13g2_decap_8 FILLER_98_749 ();
 sg13g2_decap_8 FILLER_98_756 ();
 sg13g2_decap_8 FILLER_98_763 ();
 sg13g2_decap_8 FILLER_98_770 ();
 sg13g2_decap_8 FILLER_98_777 ();
 sg13g2_decap_8 FILLER_98_784 ();
 sg13g2_decap_8 FILLER_98_791 ();
 sg13g2_decap_8 FILLER_98_798 ();
 sg13g2_decap_8 FILLER_98_805 ();
 sg13g2_decap_8 FILLER_98_812 ();
 sg13g2_decap_8 FILLER_98_819 ();
 sg13g2_decap_8 FILLER_98_826 ();
 sg13g2_decap_8 FILLER_98_833 ();
 sg13g2_fill_1 FILLER_98_840 ();
 sg13g2_decap_8 FILLER_99_0 ();
 sg13g2_decap_8 FILLER_99_7 ();
 sg13g2_decap_8 FILLER_99_14 ();
 sg13g2_decap_8 FILLER_99_21 ();
 sg13g2_decap_8 FILLER_99_28 ();
 sg13g2_decap_8 FILLER_99_35 ();
 sg13g2_decap_8 FILLER_99_42 ();
 sg13g2_decap_8 FILLER_99_49 ();
 sg13g2_decap_8 FILLER_99_56 ();
 sg13g2_decap_8 FILLER_99_63 ();
 sg13g2_decap_8 FILLER_99_70 ();
 sg13g2_decap_8 FILLER_99_77 ();
 sg13g2_decap_8 FILLER_99_84 ();
 sg13g2_decap_8 FILLER_99_91 ();
 sg13g2_decap_8 FILLER_99_98 ();
 sg13g2_decap_8 FILLER_99_105 ();
 sg13g2_decap_8 FILLER_99_112 ();
 sg13g2_decap_8 FILLER_99_119 ();
 sg13g2_decap_8 FILLER_99_126 ();
 sg13g2_decap_8 FILLER_99_133 ();
 sg13g2_decap_8 FILLER_99_140 ();
 sg13g2_decap_8 FILLER_99_147 ();
 sg13g2_decap_8 FILLER_99_154 ();
 sg13g2_decap_8 FILLER_99_161 ();
 sg13g2_decap_8 FILLER_99_168 ();
 sg13g2_decap_8 FILLER_99_175 ();
 sg13g2_decap_8 FILLER_99_182 ();
 sg13g2_decap_8 FILLER_99_189 ();
 sg13g2_decap_8 FILLER_99_196 ();
 sg13g2_decap_8 FILLER_99_203 ();
 sg13g2_decap_8 FILLER_99_210 ();
 sg13g2_decap_8 FILLER_99_217 ();
 sg13g2_decap_8 FILLER_99_224 ();
 sg13g2_decap_8 FILLER_99_231 ();
 sg13g2_decap_8 FILLER_99_238 ();
 sg13g2_decap_8 FILLER_99_245 ();
 sg13g2_decap_8 FILLER_99_252 ();
 sg13g2_decap_8 FILLER_99_259 ();
 sg13g2_decap_8 FILLER_99_266 ();
 sg13g2_decap_8 FILLER_99_273 ();
 sg13g2_decap_8 FILLER_99_280 ();
 sg13g2_decap_8 FILLER_99_287 ();
 sg13g2_decap_8 FILLER_99_294 ();
 sg13g2_decap_8 FILLER_99_301 ();
 sg13g2_decap_8 FILLER_99_308 ();
 sg13g2_decap_8 FILLER_99_315 ();
 sg13g2_decap_8 FILLER_99_322 ();
 sg13g2_decap_8 FILLER_99_329 ();
 sg13g2_decap_8 FILLER_99_336 ();
 sg13g2_decap_8 FILLER_99_343 ();
 sg13g2_decap_8 FILLER_99_350 ();
 sg13g2_decap_8 FILLER_99_357 ();
 sg13g2_decap_8 FILLER_99_364 ();
 sg13g2_decap_8 FILLER_99_371 ();
 sg13g2_decap_8 FILLER_99_378 ();
 sg13g2_decap_8 FILLER_99_385 ();
 sg13g2_decap_8 FILLER_99_392 ();
 sg13g2_decap_8 FILLER_99_399 ();
 sg13g2_decap_8 FILLER_99_406 ();
 sg13g2_decap_8 FILLER_99_413 ();
 sg13g2_decap_8 FILLER_99_420 ();
 sg13g2_decap_8 FILLER_99_427 ();
 sg13g2_decap_8 FILLER_99_434 ();
 sg13g2_decap_8 FILLER_99_441 ();
 sg13g2_decap_8 FILLER_99_448 ();
 sg13g2_decap_8 FILLER_99_455 ();
 sg13g2_decap_8 FILLER_99_462 ();
 sg13g2_decap_8 FILLER_99_469 ();
 sg13g2_decap_8 FILLER_99_476 ();
 sg13g2_decap_8 FILLER_99_483 ();
 sg13g2_decap_8 FILLER_99_490 ();
 sg13g2_decap_8 FILLER_99_497 ();
 sg13g2_decap_8 FILLER_99_504 ();
 sg13g2_decap_8 FILLER_99_511 ();
 sg13g2_decap_8 FILLER_99_518 ();
 sg13g2_decap_8 FILLER_99_525 ();
 sg13g2_decap_8 FILLER_99_532 ();
 sg13g2_decap_8 FILLER_99_539 ();
 sg13g2_decap_8 FILLER_99_546 ();
 sg13g2_decap_8 FILLER_99_553 ();
 sg13g2_decap_8 FILLER_99_560 ();
 sg13g2_decap_8 FILLER_99_567 ();
 sg13g2_decap_8 FILLER_99_574 ();
 sg13g2_decap_8 FILLER_99_581 ();
 sg13g2_decap_8 FILLER_99_588 ();
 sg13g2_decap_8 FILLER_99_595 ();
 sg13g2_decap_8 FILLER_99_602 ();
 sg13g2_decap_8 FILLER_99_609 ();
 sg13g2_decap_8 FILLER_99_616 ();
 sg13g2_decap_8 FILLER_99_623 ();
 sg13g2_decap_8 FILLER_99_630 ();
 sg13g2_decap_8 FILLER_99_637 ();
 sg13g2_decap_8 FILLER_99_644 ();
 sg13g2_decap_8 FILLER_99_651 ();
 sg13g2_decap_8 FILLER_99_658 ();
 sg13g2_decap_8 FILLER_99_665 ();
 sg13g2_decap_8 FILLER_99_672 ();
 sg13g2_decap_8 FILLER_99_679 ();
 sg13g2_decap_8 FILLER_99_686 ();
 sg13g2_decap_8 FILLER_99_693 ();
 sg13g2_decap_8 FILLER_99_700 ();
 sg13g2_decap_8 FILLER_99_707 ();
 sg13g2_decap_8 FILLER_99_714 ();
 sg13g2_decap_8 FILLER_99_721 ();
 sg13g2_decap_8 FILLER_99_728 ();
 sg13g2_decap_8 FILLER_99_735 ();
 sg13g2_decap_8 FILLER_99_742 ();
 sg13g2_decap_8 FILLER_99_749 ();
 sg13g2_decap_8 FILLER_99_756 ();
 sg13g2_decap_8 FILLER_99_763 ();
 sg13g2_decap_8 FILLER_99_770 ();
 sg13g2_decap_8 FILLER_99_777 ();
 sg13g2_decap_8 FILLER_99_784 ();
 sg13g2_decap_8 FILLER_99_791 ();
 sg13g2_decap_8 FILLER_99_798 ();
 sg13g2_decap_8 FILLER_99_805 ();
 sg13g2_decap_8 FILLER_99_812 ();
 sg13g2_decap_8 FILLER_99_819 ();
 sg13g2_decap_8 FILLER_99_826 ();
 sg13g2_decap_8 FILLER_99_833 ();
 sg13g2_fill_1 FILLER_99_840 ();
 sg13g2_decap_8 FILLER_100_0 ();
 sg13g2_decap_8 FILLER_100_7 ();
 sg13g2_decap_8 FILLER_100_14 ();
 sg13g2_decap_8 FILLER_100_21 ();
 sg13g2_decap_8 FILLER_100_28 ();
 sg13g2_decap_8 FILLER_100_35 ();
 sg13g2_decap_8 FILLER_100_42 ();
 sg13g2_decap_8 FILLER_100_49 ();
 sg13g2_decap_8 FILLER_100_56 ();
 sg13g2_decap_8 FILLER_100_63 ();
 sg13g2_decap_8 FILLER_100_70 ();
 sg13g2_decap_8 FILLER_100_77 ();
 sg13g2_decap_8 FILLER_100_84 ();
 sg13g2_decap_8 FILLER_100_91 ();
 sg13g2_decap_8 FILLER_100_98 ();
 sg13g2_decap_8 FILLER_100_105 ();
 sg13g2_decap_8 FILLER_100_112 ();
 sg13g2_decap_8 FILLER_100_119 ();
 sg13g2_decap_8 FILLER_100_126 ();
 sg13g2_decap_8 FILLER_100_133 ();
 sg13g2_decap_8 FILLER_100_140 ();
 sg13g2_decap_8 FILLER_100_147 ();
 sg13g2_decap_8 FILLER_100_154 ();
 sg13g2_decap_8 FILLER_100_161 ();
 sg13g2_decap_8 FILLER_100_168 ();
 sg13g2_decap_8 FILLER_100_175 ();
 sg13g2_decap_8 FILLER_100_182 ();
 sg13g2_decap_8 FILLER_100_189 ();
 sg13g2_decap_8 FILLER_100_196 ();
 sg13g2_decap_8 FILLER_100_203 ();
 sg13g2_decap_8 FILLER_100_210 ();
 sg13g2_decap_8 FILLER_100_217 ();
 sg13g2_decap_8 FILLER_100_224 ();
 sg13g2_decap_8 FILLER_100_231 ();
 sg13g2_decap_8 FILLER_100_238 ();
 sg13g2_decap_8 FILLER_100_245 ();
 sg13g2_decap_8 FILLER_100_252 ();
 sg13g2_decap_8 FILLER_100_259 ();
 sg13g2_decap_8 FILLER_100_266 ();
 sg13g2_decap_8 FILLER_100_273 ();
 sg13g2_decap_8 FILLER_100_280 ();
 sg13g2_decap_8 FILLER_100_287 ();
 sg13g2_decap_8 FILLER_100_294 ();
 sg13g2_decap_8 FILLER_100_301 ();
 sg13g2_decap_8 FILLER_100_308 ();
 sg13g2_decap_8 FILLER_100_315 ();
 sg13g2_decap_8 FILLER_100_322 ();
 sg13g2_decap_8 FILLER_100_329 ();
 sg13g2_decap_8 FILLER_100_336 ();
 sg13g2_decap_8 FILLER_100_343 ();
 sg13g2_decap_8 FILLER_100_350 ();
 sg13g2_decap_8 FILLER_100_357 ();
 sg13g2_decap_8 FILLER_100_364 ();
 sg13g2_decap_8 FILLER_100_371 ();
 sg13g2_decap_8 FILLER_100_378 ();
 sg13g2_decap_8 FILLER_100_385 ();
 sg13g2_decap_8 FILLER_100_392 ();
 sg13g2_decap_8 FILLER_100_399 ();
 sg13g2_decap_8 FILLER_100_406 ();
 sg13g2_decap_8 FILLER_100_413 ();
 sg13g2_decap_8 FILLER_100_420 ();
 sg13g2_decap_8 FILLER_100_427 ();
 sg13g2_decap_8 FILLER_100_434 ();
 sg13g2_decap_8 FILLER_100_441 ();
 sg13g2_decap_8 FILLER_100_448 ();
 sg13g2_decap_8 FILLER_100_455 ();
 sg13g2_decap_8 FILLER_100_462 ();
 sg13g2_decap_8 FILLER_100_469 ();
 sg13g2_decap_8 FILLER_100_476 ();
 sg13g2_decap_8 FILLER_100_483 ();
 sg13g2_decap_8 FILLER_100_490 ();
 sg13g2_decap_8 FILLER_100_497 ();
 sg13g2_decap_8 FILLER_100_504 ();
 sg13g2_decap_8 FILLER_100_511 ();
 sg13g2_decap_8 FILLER_100_518 ();
 sg13g2_decap_8 FILLER_100_525 ();
 sg13g2_decap_8 FILLER_100_532 ();
 sg13g2_decap_8 FILLER_100_539 ();
 sg13g2_decap_8 FILLER_100_546 ();
 sg13g2_decap_8 FILLER_100_553 ();
 sg13g2_decap_8 FILLER_100_560 ();
 sg13g2_decap_8 FILLER_100_567 ();
 sg13g2_decap_8 FILLER_100_574 ();
 sg13g2_decap_8 FILLER_100_581 ();
 sg13g2_decap_8 FILLER_100_588 ();
 sg13g2_decap_8 FILLER_100_595 ();
 sg13g2_decap_8 FILLER_100_602 ();
 sg13g2_decap_8 FILLER_100_609 ();
 sg13g2_decap_8 FILLER_100_616 ();
 sg13g2_decap_8 FILLER_100_623 ();
 sg13g2_decap_8 FILLER_100_630 ();
 sg13g2_decap_8 FILLER_100_637 ();
 sg13g2_decap_8 FILLER_100_644 ();
 sg13g2_decap_8 FILLER_100_651 ();
 sg13g2_decap_8 FILLER_100_658 ();
 sg13g2_decap_8 FILLER_100_665 ();
 sg13g2_decap_8 FILLER_100_672 ();
 sg13g2_decap_8 FILLER_100_679 ();
 sg13g2_decap_8 FILLER_100_686 ();
 sg13g2_decap_8 FILLER_100_693 ();
 sg13g2_decap_8 FILLER_100_700 ();
 sg13g2_decap_8 FILLER_100_707 ();
 sg13g2_decap_8 FILLER_100_714 ();
 sg13g2_decap_8 FILLER_100_721 ();
 sg13g2_decap_8 FILLER_100_728 ();
 sg13g2_decap_8 FILLER_100_735 ();
 sg13g2_decap_8 FILLER_100_742 ();
 sg13g2_decap_8 FILLER_100_749 ();
 sg13g2_decap_8 FILLER_100_756 ();
 sg13g2_decap_8 FILLER_100_763 ();
 sg13g2_decap_8 FILLER_100_770 ();
 sg13g2_decap_8 FILLER_100_777 ();
 sg13g2_decap_8 FILLER_100_784 ();
 sg13g2_decap_8 FILLER_100_791 ();
 sg13g2_decap_8 FILLER_100_798 ();
 sg13g2_decap_8 FILLER_100_805 ();
 sg13g2_decap_8 FILLER_100_812 ();
 sg13g2_decap_8 FILLER_100_819 ();
 sg13g2_decap_8 FILLER_100_826 ();
 sg13g2_decap_8 FILLER_100_833 ();
 sg13g2_fill_1 FILLER_100_840 ();
 sg13g2_decap_8 FILLER_101_0 ();
 sg13g2_decap_8 FILLER_101_7 ();
 sg13g2_decap_8 FILLER_101_14 ();
 sg13g2_decap_8 FILLER_101_21 ();
 sg13g2_decap_8 FILLER_101_28 ();
 sg13g2_decap_8 FILLER_101_35 ();
 sg13g2_decap_8 FILLER_101_42 ();
 sg13g2_decap_8 FILLER_101_49 ();
 sg13g2_decap_8 FILLER_101_56 ();
 sg13g2_decap_8 FILLER_101_63 ();
 sg13g2_decap_8 FILLER_101_70 ();
 sg13g2_decap_8 FILLER_101_77 ();
 sg13g2_decap_8 FILLER_101_84 ();
 sg13g2_decap_8 FILLER_101_91 ();
 sg13g2_decap_8 FILLER_101_98 ();
 sg13g2_decap_8 FILLER_101_105 ();
 sg13g2_decap_8 FILLER_101_112 ();
 sg13g2_decap_8 FILLER_101_119 ();
 sg13g2_decap_8 FILLER_101_126 ();
 sg13g2_decap_8 FILLER_101_133 ();
 sg13g2_decap_8 FILLER_101_140 ();
 sg13g2_decap_8 FILLER_101_147 ();
 sg13g2_decap_8 FILLER_101_154 ();
 sg13g2_decap_8 FILLER_101_161 ();
 sg13g2_decap_8 FILLER_101_168 ();
 sg13g2_decap_8 FILLER_101_175 ();
 sg13g2_decap_8 FILLER_101_182 ();
 sg13g2_decap_8 FILLER_101_189 ();
 sg13g2_decap_8 FILLER_101_196 ();
 sg13g2_decap_8 FILLER_101_203 ();
 sg13g2_decap_8 FILLER_101_210 ();
 sg13g2_decap_8 FILLER_101_217 ();
 sg13g2_decap_8 FILLER_101_224 ();
 sg13g2_decap_8 FILLER_101_231 ();
 sg13g2_decap_8 FILLER_101_238 ();
 sg13g2_decap_8 FILLER_101_245 ();
 sg13g2_decap_8 FILLER_101_252 ();
 sg13g2_decap_8 FILLER_101_259 ();
 sg13g2_decap_8 FILLER_101_266 ();
 sg13g2_decap_8 FILLER_101_273 ();
 sg13g2_decap_8 FILLER_101_280 ();
 sg13g2_decap_8 FILLER_101_287 ();
 sg13g2_decap_8 FILLER_101_294 ();
 sg13g2_decap_8 FILLER_101_301 ();
 sg13g2_decap_8 FILLER_101_308 ();
 sg13g2_decap_8 FILLER_101_315 ();
 sg13g2_decap_8 FILLER_101_322 ();
 sg13g2_decap_8 FILLER_101_329 ();
 sg13g2_decap_8 FILLER_101_336 ();
 sg13g2_decap_8 FILLER_101_343 ();
 sg13g2_decap_8 FILLER_101_350 ();
 sg13g2_decap_8 FILLER_101_357 ();
 sg13g2_decap_8 FILLER_101_364 ();
 sg13g2_decap_8 FILLER_101_371 ();
 sg13g2_decap_8 FILLER_101_378 ();
 sg13g2_decap_8 FILLER_101_385 ();
 sg13g2_decap_8 FILLER_101_392 ();
 sg13g2_decap_8 FILLER_101_399 ();
 sg13g2_decap_8 FILLER_101_406 ();
 sg13g2_decap_8 FILLER_101_413 ();
 sg13g2_decap_8 FILLER_101_420 ();
 sg13g2_decap_8 FILLER_101_427 ();
 sg13g2_decap_8 FILLER_101_434 ();
 sg13g2_decap_8 FILLER_101_441 ();
 sg13g2_decap_8 FILLER_101_448 ();
 sg13g2_decap_8 FILLER_101_455 ();
 sg13g2_decap_8 FILLER_101_462 ();
 sg13g2_decap_8 FILLER_101_469 ();
 sg13g2_decap_8 FILLER_101_476 ();
 sg13g2_decap_8 FILLER_101_483 ();
 sg13g2_decap_8 FILLER_101_490 ();
 sg13g2_decap_8 FILLER_101_497 ();
 sg13g2_decap_8 FILLER_101_504 ();
 sg13g2_decap_8 FILLER_101_511 ();
 sg13g2_decap_8 FILLER_101_518 ();
 sg13g2_decap_8 FILLER_101_525 ();
 sg13g2_decap_8 FILLER_101_532 ();
 sg13g2_decap_8 FILLER_101_539 ();
 sg13g2_decap_8 FILLER_101_546 ();
 sg13g2_decap_8 FILLER_101_553 ();
 sg13g2_decap_8 FILLER_101_560 ();
 sg13g2_decap_8 FILLER_101_567 ();
 sg13g2_decap_8 FILLER_101_574 ();
 sg13g2_decap_8 FILLER_101_581 ();
 sg13g2_decap_8 FILLER_101_588 ();
 sg13g2_decap_8 FILLER_101_595 ();
 sg13g2_decap_8 FILLER_101_602 ();
 sg13g2_decap_8 FILLER_101_609 ();
 sg13g2_decap_8 FILLER_101_616 ();
 sg13g2_decap_8 FILLER_101_623 ();
 sg13g2_decap_8 FILLER_101_630 ();
 sg13g2_decap_8 FILLER_101_637 ();
 sg13g2_decap_8 FILLER_101_644 ();
 sg13g2_decap_8 FILLER_101_651 ();
 sg13g2_decap_8 FILLER_101_658 ();
 sg13g2_decap_8 FILLER_101_665 ();
 sg13g2_decap_8 FILLER_101_672 ();
 sg13g2_decap_8 FILLER_101_679 ();
 sg13g2_decap_8 FILLER_101_686 ();
 sg13g2_decap_8 FILLER_101_693 ();
 sg13g2_decap_8 FILLER_101_700 ();
 sg13g2_decap_8 FILLER_101_707 ();
 sg13g2_decap_8 FILLER_101_714 ();
 sg13g2_decap_8 FILLER_101_721 ();
 sg13g2_decap_8 FILLER_101_728 ();
 sg13g2_decap_8 FILLER_101_735 ();
 sg13g2_decap_8 FILLER_101_742 ();
 sg13g2_decap_8 FILLER_101_749 ();
 sg13g2_decap_8 FILLER_101_756 ();
 sg13g2_decap_8 FILLER_101_763 ();
 sg13g2_decap_8 FILLER_101_770 ();
 sg13g2_decap_8 FILLER_101_777 ();
 sg13g2_decap_8 FILLER_101_784 ();
 sg13g2_decap_8 FILLER_101_791 ();
 sg13g2_decap_8 FILLER_101_798 ();
 sg13g2_decap_8 FILLER_101_805 ();
 sg13g2_decap_8 FILLER_101_812 ();
 sg13g2_decap_8 FILLER_101_819 ();
 sg13g2_decap_8 FILLER_101_826 ();
 sg13g2_decap_8 FILLER_101_833 ();
 sg13g2_fill_1 FILLER_101_840 ();
 sg13g2_decap_8 FILLER_102_0 ();
 sg13g2_decap_8 FILLER_102_7 ();
 sg13g2_decap_8 FILLER_102_14 ();
 sg13g2_decap_8 FILLER_102_21 ();
 sg13g2_decap_8 FILLER_102_28 ();
 sg13g2_decap_8 FILLER_102_35 ();
 sg13g2_decap_8 FILLER_102_42 ();
 sg13g2_decap_8 FILLER_102_49 ();
 sg13g2_decap_8 FILLER_102_56 ();
 sg13g2_decap_8 FILLER_102_63 ();
 sg13g2_decap_8 FILLER_102_70 ();
 sg13g2_decap_8 FILLER_102_77 ();
 sg13g2_decap_8 FILLER_102_84 ();
 sg13g2_decap_8 FILLER_102_91 ();
 sg13g2_decap_8 FILLER_102_98 ();
 sg13g2_decap_8 FILLER_102_105 ();
 sg13g2_decap_8 FILLER_102_112 ();
 sg13g2_decap_8 FILLER_102_119 ();
 sg13g2_decap_8 FILLER_102_126 ();
 sg13g2_decap_8 FILLER_102_133 ();
 sg13g2_decap_8 FILLER_102_140 ();
 sg13g2_decap_8 FILLER_102_147 ();
 sg13g2_decap_8 FILLER_102_154 ();
 sg13g2_decap_8 FILLER_102_161 ();
 sg13g2_decap_8 FILLER_102_168 ();
 sg13g2_decap_8 FILLER_102_175 ();
 sg13g2_decap_8 FILLER_102_182 ();
 sg13g2_decap_8 FILLER_102_189 ();
 sg13g2_decap_8 FILLER_102_196 ();
 sg13g2_decap_8 FILLER_102_203 ();
 sg13g2_decap_8 FILLER_102_210 ();
 sg13g2_decap_8 FILLER_102_217 ();
 sg13g2_decap_8 FILLER_102_224 ();
 sg13g2_decap_8 FILLER_102_231 ();
 sg13g2_decap_8 FILLER_102_238 ();
 sg13g2_decap_8 FILLER_102_245 ();
 sg13g2_decap_8 FILLER_102_252 ();
 sg13g2_decap_8 FILLER_102_259 ();
 sg13g2_decap_8 FILLER_102_266 ();
 sg13g2_decap_8 FILLER_102_273 ();
 sg13g2_decap_8 FILLER_102_280 ();
 sg13g2_decap_8 FILLER_102_287 ();
 sg13g2_decap_8 FILLER_102_294 ();
 sg13g2_decap_8 FILLER_102_301 ();
 sg13g2_decap_8 FILLER_102_308 ();
 sg13g2_decap_8 FILLER_102_315 ();
 sg13g2_decap_8 FILLER_102_322 ();
 sg13g2_decap_8 FILLER_102_329 ();
 sg13g2_decap_8 FILLER_102_336 ();
 sg13g2_decap_8 FILLER_102_343 ();
 sg13g2_decap_8 FILLER_102_350 ();
 sg13g2_decap_8 FILLER_102_357 ();
 sg13g2_decap_8 FILLER_102_364 ();
 sg13g2_decap_8 FILLER_102_371 ();
 sg13g2_decap_8 FILLER_102_378 ();
 sg13g2_decap_8 FILLER_102_385 ();
 sg13g2_decap_8 FILLER_102_392 ();
 sg13g2_decap_8 FILLER_102_399 ();
 sg13g2_decap_8 FILLER_102_406 ();
 sg13g2_decap_8 FILLER_102_413 ();
 sg13g2_decap_8 FILLER_102_420 ();
 sg13g2_decap_8 FILLER_102_427 ();
 sg13g2_decap_8 FILLER_102_434 ();
 sg13g2_decap_8 FILLER_102_441 ();
 sg13g2_decap_8 FILLER_102_448 ();
 sg13g2_decap_8 FILLER_102_455 ();
 sg13g2_decap_8 FILLER_102_462 ();
 sg13g2_decap_8 FILLER_102_469 ();
 sg13g2_decap_8 FILLER_102_476 ();
 sg13g2_decap_8 FILLER_102_483 ();
 sg13g2_decap_8 FILLER_102_490 ();
 sg13g2_decap_8 FILLER_102_497 ();
 sg13g2_decap_8 FILLER_102_504 ();
 sg13g2_decap_8 FILLER_102_511 ();
 sg13g2_decap_8 FILLER_102_518 ();
 sg13g2_decap_8 FILLER_102_525 ();
 sg13g2_decap_8 FILLER_102_532 ();
 sg13g2_decap_8 FILLER_102_539 ();
 sg13g2_decap_8 FILLER_102_546 ();
 sg13g2_decap_8 FILLER_102_553 ();
 sg13g2_decap_8 FILLER_102_560 ();
 sg13g2_decap_8 FILLER_102_567 ();
 sg13g2_decap_8 FILLER_102_574 ();
 sg13g2_decap_8 FILLER_102_581 ();
 sg13g2_decap_8 FILLER_102_588 ();
 sg13g2_decap_8 FILLER_102_595 ();
 sg13g2_decap_8 FILLER_102_602 ();
 sg13g2_decap_8 FILLER_102_609 ();
 sg13g2_decap_8 FILLER_102_616 ();
 sg13g2_decap_8 FILLER_102_623 ();
 sg13g2_decap_8 FILLER_102_630 ();
 sg13g2_decap_8 FILLER_102_637 ();
 sg13g2_decap_8 FILLER_102_644 ();
 sg13g2_decap_8 FILLER_102_651 ();
 sg13g2_decap_8 FILLER_102_658 ();
 sg13g2_decap_8 FILLER_102_665 ();
 sg13g2_decap_8 FILLER_102_672 ();
 sg13g2_decap_8 FILLER_102_679 ();
 sg13g2_decap_8 FILLER_102_686 ();
 sg13g2_decap_8 FILLER_102_693 ();
 sg13g2_decap_8 FILLER_102_700 ();
 sg13g2_decap_8 FILLER_102_707 ();
 sg13g2_decap_8 FILLER_102_714 ();
 sg13g2_decap_8 FILLER_102_721 ();
 sg13g2_decap_8 FILLER_102_728 ();
 sg13g2_decap_8 FILLER_102_735 ();
 sg13g2_decap_8 FILLER_102_742 ();
 sg13g2_decap_8 FILLER_102_749 ();
 sg13g2_decap_8 FILLER_102_756 ();
 sg13g2_decap_8 FILLER_102_763 ();
 sg13g2_decap_8 FILLER_102_770 ();
 sg13g2_decap_8 FILLER_102_777 ();
 sg13g2_decap_8 FILLER_102_784 ();
 sg13g2_decap_8 FILLER_102_791 ();
 sg13g2_decap_8 FILLER_102_798 ();
 sg13g2_decap_8 FILLER_102_805 ();
 sg13g2_decap_8 FILLER_102_812 ();
 sg13g2_decap_8 FILLER_102_819 ();
 sg13g2_decap_8 FILLER_102_826 ();
 sg13g2_decap_8 FILLER_102_833 ();
 sg13g2_fill_1 FILLER_102_840 ();
 sg13g2_decap_8 FILLER_103_0 ();
 sg13g2_decap_8 FILLER_103_7 ();
 sg13g2_decap_8 FILLER_103_14 ();
 sg13g2_decap_8 FILLER_103_21 ();
 sg13g2_decap_8 FILLER_103_28 ();
 sg13g2_decap_8 FILLER_103_35 ();
 sg13g2_decap_8 FILLER_103_42 ();
 sg13g2_decap_8 FILLER_103_49 ();
 sg13g2_decap_8 FILLER_103_56 ();
 sg13g2_decap_8 FILLER_103_63 ();
 sg13g2_decap_8 FILLER_103_70 ();
 sg13g2_decap_8 FILLER_103_77 ();
 sg13g2_decap_8 FILLER_103_84 ();
 sg13g2_decap_8 FILLER_103_91 ();
 sg13g2_decap_8 FILLER_103_98 ();
 sg13g2_decap_8 FILLER_103_105 ();
 sg13g2_decap_8 FILLER_103_112 ();
 sg13g2_decap_8 FILLER_103_119 ();
 sg13g2_decap_8 FILLER_103_126 ();
 sg13g2_decap_8 FILLER_103_133 ();
 sg13g2_decap_8 FILLER_103_140 ();
 sg13g2_decap_8 FILLER_103_147 ();
 sg13g2_decap_8 FILLER_103_154 ();
 sg13g2_decap_8 FILLER_103_161 ();
 sg13g2_decap_8 FILLER_103_168 ();
 sg13g2_decap_8 FILLER_103_175 ();
 sg13g2_decap_8 FILLER_103_182 ();
 sg13g2_decap_8 FILLER_103_189 ();
 sg13g2_decap_8 FILLER_103_196 ();
 sg13g2_decap_8 FILLER_103_203 ();
 sg13g2_decap_8 FILLER_103_210 ();
 sg13g2_decap_8 FILLER_103_217 ();
 sg13g2_decap_8 FILLER_103_224 ();
 sg13g2_decap_8 FILLER_103_231 ();
 sg13g2_decap_8 FILLER_103_238 ();
 sg13g2_decap_8 FILLER_103_245 ();
 sg13g2_decap_8 FILLER_103_252 ();
 sg13g2_decap_8 FILLER_103_259 ();
 sg13g2_decap_8 FILLER_103_266 ();
 sg13g2_decap_8 FILLER_103_273 ();
 sg13g2_decap_8 FILLER_103_280 ();
 sg13g2_decap_8 FILLER_103_287 ();
 sg13g2_decap_8 FILLER_103_294 ();
 sg13g2_decap_8 FILLER_103_301 ();
 sg13g2_decap_8 FILLER_103_308 ();
 sg13g2_decap_8 FILLER_103_315 ();
 sg13g2_decap_8 FILLER_103_322 ();
 sg13g2_decap_8 FILLER_103_329 ();
 sg13g2_decap_8 FILLER_103_336 ();
 sg13g2_decap_8 FILLER_103_343 ();
 sg13g2_decap_8 FILLER_103_350 ();
 sg13g2_decap_8 FILLER_103_357 ();
 sg13g2_decap_8 FILLER_103_364 ();
 sg13g2_decap_8 FILLER_103_371 ();
 sg13g2_decap_8 FILLER_103_378 ();
 sg13g2_decap_8 FILLER_103_385 ();
 sg13g2_decap_8 FILLER_103_392 ();
 sg13g2_decap_8 FILLER_103_399 ();
 sg13g2_decap_8 FILLER_103_406 ();
 sg13g2_decap_8 FILLER_103_413 ();
 sg13g2_decap_8 FILLER_103_420 ();
 sg13g2_decap_8 FILLER_103_427 ();
 sg13g2_decap_8 FILLER_103_434 ();
 sg13g2_decap_8 FILLER_103_441 ();
 sg13g2_decap_8 FILLER_103_448 ();
 sg13g2_decap_8 FILLER_103_455 ();
 sg13g2_decap_8 FILLER_103_462 ();
 sg13g2_decap_8 FILLER_103_469 ();
 sg13g2_decap_8 FILLER_103_476 ();
 sg13g2_decap_8 FILLER_103_483 ();
 sg13g2_decap_8 FILLER_103_490 ();
 sg13g2_decap_8 FILLER_103_497 ();
 sg13g2_decap_8 FILLER_103_504 ();
 sg13g2_decap_8 FILLER_103_511 ();
 sg13g2_decap_8 FILLER_103_518 ();
 sg13g2_decap_8 FILLER_103_525 ();
 sg13g2_decap_8 FILLER_103_532 ();
 sg13g2_decap_8 FILLER_103_539 ();
 sg13g2_decap_8 FILLER_103_546 ();
 sg13g2_decap_8 FILLER_103_553 ();
 sg13g2_decap_8 FILLER_103_560 ();
 sg13g2_decap_8 FILLER_103_567 ();
 sg13g2_decap_8 FILLER_103_574 ();
 sg13g2_decap_8 FILLER_103_581 ();
 sg13g2_decap_8 FILLER_103_588 ();
 sg13g2_decap_8 FILLER_103_595 ();
 sg13g2_decap_8 FILLER_103_602 ();
 sg13g2_decap_8 FILLER_103_609 ();
 sg13g2_decap_8 FILLER_103_616 ();
 sg13g2_decap_8 FILLER_103_623 ();
 sg13g2_decap_8 FILLER_103_630 ();
 sg13g2_decap_8 FILLER_103_637 ();
 sg13g2_decap_8 FILLER_103_644 ();
 sg13g2_decap_8 FILLER_103_651 ();
 sg13g2_decap_8 FILLER_103_658 ();
 sg13g2_decap_8 FILLER_103_665 ();
 sg13g2_decap_8 FILLER_103_672 ();
 sg13g2_decap_8 FILLER_103_679 ();
 sg13g2_decap_8 FILLER_103_686 ();
 sg13g2_decap_8 FILLER_103_693 ();
 sg13g2_decap_8 FILLER_103_700 ();
 sg13g2_decap_8 FILLER_103_707 ();
 sg13g2_decap_8 FILLER_103_714 ();
 sg13g2_decap_8 FILLER_103_721 ();
 sg13g2_decap_8 FILLER_103_728 ();
 sg13g2_decap_8 FILLER_103_735 ();
 sg13g2_decap_8 FILLER_103_742 ();
 sg13g2_decap_8 FILLER_103_749 ();
 sg13g2_decap_8 FILLER_103_756 ();
 sg13g2_decap_8 FILLER_103_763 ();
 sg13g2_decap_8 FILLER_103_770 ();
 sg13g2_decap_8 FILLER_103_777 ();
 sg13g2_decap_8 FILLER_103_784 ();
 sg13g2_decap_8 FILLER_103_791 ();
 sg13g2_decap_8 FILLER_103_798 ();
 sg13g2_decap_8 FILLER_103_805 ();
 sg13g2_decap_8 FILLER_103_812 ();
 sg13g2_decap_8 FILLER_103_819 ();
 sg13g2_decap_8 FILLER_103_826 ();
 sg13g2_decap_8 FILLER_103_833 ();
 sg13g2_fill_1 FILLER_103_840 ();
 sg13g2_decap_8 FILLER_104_0 ();
 sg13g2_decap_8 FILLER_104_7 ();
 sg13g2_decap_8 FILLER_104_14 ();
 sg13g2_decap_8 FILLER_104_21 ();
 sg13g2_decap_8 FILLER_104_28 ();
 sg13g2_decap_8 FILLER_104_35 ();
 sg13g2_decap_8 FILLER_104_42 ();
 sg13g2_decap_8 FILLER_104_49 ();
 sg13g2_decap_8 FILLER_104_56 ();
 sg13g2_decap_8 FILLER_104_63 ();
 sg13g2_decap_8 FILLER_104_70 ();
 sg13g2_decap_8 FILLER_104_77 ();
 sg13g2_decap_8 FILLER_104_84 ();
 sg13g2_decap_8 FILLER_104_91 ();
 sg13g2_decap_8 FILLER_104_98 ();
 sg13g2_decap_8 FILLER_104_105 ();
 sg13g2_decap_8 FILLER_104_112 ();
 sg13g2_decap_8 FILLER_104_119 ();
 sg13g2_decap_8 FILLER_104_126 ();
 sg13g2_decap_8 FILLER_104_133 ();
 sg13g2_decap_8 FILLER_104_140 ();
 sg13g2_decap_8 FILLER_104_147 ();
 sg13g2_decap_8 FILLER_104_154 ();
 sg13g2_decap_8 FILLER_104_161 ();
 sg13g2_decap_8 FILLER_104_168 ();
 sg13g2_decap_8 FILLER_104_175 ();
 sg13g2_decap_8 FILLER_104_182 ();
 sg13g2_decap_8 FILLER_104_189 ();
 sg13g2_decap_8 FILLER_104_196 ();
 sg13g2_decap_8 FILLER_104_203 ();
 sg13g2_decap_8 FILLER_104_210 ();
 sg13g2_decap_8 FILLER_104_217 ();
 sg13g2_decap_8 FILLER_104_224 ();
 sg13g2_decap_8 FILLER_104_231 ();
 sg13g2_decap_8 FILLER_104_238 ();
 sg13g2_decap_8 FILLER_104_245 ();
 sg13g2_decap_8 FILLER_104_252 ();
 sg13g2_decap_8 FILLER_104_259 ();
 sg13g2_decap_8 FILLER_104_266 ();
 sg13g2_decap_8 FILLER_104_273 ();
 sg13g2_decap_8 FILLER_104_280 ();
 sg13g2_decap_8 FILLER_104_287 ();
 sg13g2_decap_8 FILLER_104_294 ();
 sg13g2_decap_8 FILLER_104_301 ();
 sg13g2_decap_8 FILLER_104_308 ();
 sg13g2_decap_8 FILLER_104_315 ();
 sg13g2_decap_8 FILLER_104_322 ();
 sg13g2_decap_8 FILLER_104_329 ();
 sg13g2_decap_8 FILLER_104_336 ();
 sg13g2_decap_8 FILLER_104_343 ();
 sg13g2_decap_8 FILLER_104_350 ();
 sg13g2_decap_8 FILLER_104_357 ();
 sg13g2_decap_8 FILLER_104_364 ();
 sg13g2_decap_8 FILLER_104_371 ();
 sg13g2_decap_8 FILLER_104_378 ();
 sg13g2_decap_8 FILLER_104_385 ();
 sg13g2_decap_8 FILLER_104_392 ();
 sg13g2_decap_8 FILLER_104_399 ();
 sg13g2_decap_8 FILLER_104_406 ();
 sg13g2_decap_8 FILLER_104_413 ();
 sg13g2_decap_8 FILLER_104_420 ();
 sg13g2_decap_8 FILLER_104_427 ();
 sg13g2_decap_8 FILLER_104_434 ();
 sg13g2_decap_8 FILLER_104_441 ();
 sg13g2_decap_8 FILLER_104_448 ();
 sg13g2_decap_8 FILLER_104_455 ();
 sg13g2_decap_8 FILLER_104_462 ();
 sg13g2_decap_8 FILLER_104_469 ();
 sg13g2_decap_8 FILLER_104_476 ();
 sg13g2_decap_8 FILLER_104_483 ();
 sg13g2_decap_8 FILLER_104_490 ();
 sg13g2_decap_8 FILLER_104_497 ();
 sg13g2_decap_8 FILLER_104_504 ();
 sg13g2_decap_8 FILLER_104_511 ();
 sg13g2_decap_8 FILLER_104_518 ();
 sg13g2_decap_8 FILLER_104_525 ();
 sg13g2_decap_8 FILLER_104_532 ();
 sg13g2_decap_8 FILLER_104_539 ();
 sg13g2_decap_8 FILLER_104_546 ();
 sg13g2_decap_8 FILLER_104_553 ();
 sg13g2_decap_8 FILLER_104_560 ();
 sg13g2_decap_8 FILLER_104_567 ();
 sg13g2_decap_8 FILLER_104_574 ();
 sg13g2_decap_8 FILLER_104_581 ();
 sg13g2_decap_8 FILLER_104_588 ();
 sg13g2_decap_8 FILLER_104_595 ();
 sg13g2_decap_8 FILLER_104_602 ();
 sg13g2_decap_8 FILLER_104_609 ();
 sg13g2_decap_8 FILLER_104_616 ();
 sg13g2_decap_8 FILLER_104_623 ();
 sg13g2_decap_8 FILLER_104_630 ();
 sg13g2_decap_8 FILLER_104_637 ();
 sg13g2_decap_8 FILLER_104_644 ();
 sg13g2_decap_8 FILLER_104_651 ();
 sg13g2_decap_8 FILLER_104_658 ();
 sg13g2_decap_8 FILLER_104_665 ();
 sg13g2_decap_8 FILLER_104_672 ();
 sg13g2_decap_8 FILLER_104_679 ();
 sg13g2_decap_8 FILLER_104_686 ();
 sg13g2_decap_8 FILLER_104_693 ();
 sg13g2_decap_8 FILLER_104_700 ();
 sg13g2_decap_8 FILLER_104_707 ();
 sg13g2_decap_8 FILLER_104_714 ();
 sg13g2_decap_8 FILLER_104_721 ();
 sg13g2_decap_8 FILLER_104_728 ();
 sg13g2_decap_8 FILLER_104_735 ();
 sg13g2_decap_8 FILLER_104_742 ();
 sg13g2_decap_8 FILLER_104_749 ();
 sg13g2_decap_8 FILLER_104_756 ();
 sg13g2_decap_8 FILLER_104_763 ();
 sg13g2_decap_8 FILLER_104_770 ();
 sg13g2_decap_8 FILLER_104_777 ();
 sg13g2_decap_8 FILLER_104_784 ();
 sg13g2_decap_8 FILLER_104_791 ();
 sg13g2_decap_8 FILLER_104_798 ();
 sg13g2_decap_8 FILLER_104_805 ();
 sg13g2_decap_8 FILLER_104_812 ();
 sg13g2_decap_8 FILLER_104_819 ();
 sg13g2_decap_8 FILLER_104_826 ();
 sg13g2_decap_8 FILLER_104_833 ();
 sg13g2_fill_1 FILLER_104_840 ();
 sg13g2_decap_8 FILLER_105_0 ();
 sg13g2_decap_8 FILLER_105_7 ();
 sg13g2_decap_8 FILLER_105_14 ();
 sg13g2_decap_8 FILLER_105_21 ();
 sg13g2_decap_8 FILLER_105_28 ();
 sg13g2_decap_8 FILLER_105_35 ();
 sg13g2_decap_8 FILLER_105_42 ();
 sg13g2_decap_8 FILLER_105_49 ();
 sg13g2_decap_8 FILLER_105_56 ();
 sg13g2_decap_8 FILLER_105_63 ();
 sg13g2_decap_8 FILLER_105_70 ();
 sg13g2_decap_8 FILLER_105_77 ();
 sg13g2_decap_8 FILLER_105_84 ();
 sg13g2_decap_8 FILLER_105_91 ();
 sg13g2_decap_8 FILLER_105_98 ();
 sg13g2_decap_8 FILLER_105_105 ();
 sg13g2_decap_8 FILLER_105_112 ();
 sg13g2_decap_8 FILLER_105_119 ();
 sg13g2_decap_8 FILLER_105_126 ();
 sg13g2_decap_8 FILLER_105_133 ();
 sg13g2_decap_8 FILLER_105_140 ();
 sg13g2_decap_8 FILLER_105_147 ();
 sg13g2_decap_8 FILLER_105_154 ();
 sg13g2_decap_8 FILLER_105_161 ();
 sg13g2_decap_8 FILLER_105_168 ();
 sg13g2_decap_8 FILLER_105_175 ();
 sg13g2_decap_8 FILLER_105_182 ();
 sg13g2_decap_8 FILLER_105_189 ();
 sg13g2_decap_8 FILLER_105_196 ();
 sg13g2_decap_8 FILLER_105_203 ();
 sg13g2_decap_8 FILLER_105_210 ();
 sg13g2_decap_8 FILLER_105_217 ();
 sg13g2_decap_8 FILLER_105_224 ();
 sg13g2_decap_8 FILLER_105_231 ();
 sg13g2_decap_8 FILLER_105_238 ();
 sg13g2_decap_8 FILLER_105_245 ();
 sg13g2_decap_8 FILLER_105_252 ();
 sg13g2_decap_8 FILLER_105_259 ();
 sg13g2_decap_8 FILLER_105_266 ();
 sg13g2_decap_8 FILLER_105_273 ();
 sg13g2_decap_8 FILLER_105_280 ();
 sg13g2_decap_8 FILLER_105_287 ();
 sg13g2_decap_8 FILLER_105_294 ();
 sg13g2_decap_8 FILLER_105_301 ();
 sg13g2_decap_8 FILLER_105_308 ();
 sg13g2_decap_8 FILLER_105_315 ();
 sg13g2_decap_8 FILLER_105_322 ();
 sg13g2_decap_8 FILLER_105_329 ();
 sg13g2_decap_8 FILLER_105_336 ();
 sg13g2_decap_8 FILLER_105_343 ();
 sg13g2_decap_8 FILLER_105_350 ();
 sg13g2_decap_8 FILLER_105_357 ();
 sg13g2_decap_8 FILLER_105_364 ();
 sg13g2_decap_8 FILLER_105_371 ();
 sg13g2_decap_8 FILLER_105_378 ();
 sg13g2_decap_8 FILLER_105_385 ();
 sg13g2_decap_8 FILLER_105_392 ();
 sg13g2_decap_8 FILLER_105_399 ();
 sg13g2_decap_8 FILLER_105_406 ();
 sg13g2_decap_8 FILLER_105_413 ();
 sg13g2_decap_8 FILLER_105_420 ();
 sg13g2_decap_8 FILLER_105_427 ();
 sg13g2_decap_8 FILLER_105_434 ();
 sg13g2_decap_8 FILLER_105_441 ();
 sg13g2_decap_8 FILLER_105_448 ();
 sg13g2_decap_8 FILLER_105_455 ();
 sg13g2_decap_8 FILLER_105_462 ();
 sg13g2_decap_8 FILLER_105_469 ();
 sg13g2_decap_8 FILLER_105_476 ();
 sg13g2_decap_8 FILLER_105_483 ();
 sg13g2_decap_8 FILLER_105_490 ();
 sg13g2_decap_8 FILLER_105_497 ();
 sg13g2_decap_8 FILLER_105_504 ();
 sg13g2_decap_8 FILLER_105_511 ();
 sg13g2_decap_8 FILLER_105_518 ();
 sg13g2_decap_8 FILLER_105_525 ();
 sg13g2_decap_8 FILLER_105_532 ();
 sg13g2_decap_8 FILLER_105_539 ();
 sg13g2_decap_8 FILLER_105_546 ();
 sg13g2_decap_8 FILLER_105_553 ();
 sg13g2_decap_8 FILLER_105_560 ();
 sg13g2_decap_8 FILLER_105_567 ();
 sg13g2_decap_8 FILLER_105_574 ();
 sg13g2_decap_8 FILLER_105_581 ();
 sg13g2_decap_8 FILLER_105_588 ();
 sg13g2_decap_8 FILLER_105_595 ();
 sg13g2_decap_8 FILLER_105_602 ();
 sg13g2_decap_8 FILLER_105_609 ();
 sg13g2_decap_8 FILLER_105_616 ();
 sg13g2_decap_8 FILLER_105_623 ();
 sg13g2_decap_8 FILLER_105_630 ();
 sg13g2_decap_8 FILLER_105_637 ();
 sg13g2_decap_8 FILLER_105_644 ();
 sg13g2_decap_8 FILLER_105_651 ();
 sg13g2_decap_8 FILLER_105_658 ();
 sg13g2_decap_8 FILLER_105_665 ();
 sg13g2_decap_8 FILLER_105_672 ();
 sg13g2_decap_8 FILLER_105_679 ();
 sg13g2_decap_8 FILLER_105_686 ();
 sg13g2_decap_8 FILLER_105_693 ();
 sg13g2_decap_8 FILLER_105_700 ();
 sg13g2_decap_8 FILLER_105_707 ();
 sg13g2_decap_8 FILLER_105_714 ();
 sg13g2_decap_8 FILLER_105_721 ();
 sg13g2_decap_8 FILLER_105_728 ();
 sg13g2_decap_8 FILLER_105_735 ();
 sg13g2_decap_8 FILLER_105_742 ();
 sg13g2_decap_8 FILLER_105_749 ();
 sg13g2_decap_8 FILLER_105_756 ();
 sg13g2_decap_8 FILLER_105_763 ();
 sg13g2_decap_8 FILLER_105_770 ();
 sg13g2_decap_8 FILLER_105_777 ();
 sg13g2_decap_8 FILLER_105_784 ();
 sg13g2_decap_8 FILLER_105_791 ();
 sg13g2_decap_8 FILLER_105_798 ();
 sg13g2_decap_8 FILLER_105_805 ();
 sg13g2_decap_8 FILLER_105_812 ();
 sg13g2_decap_8 FILLER_105_819 ();
 sg13g2_decap_8 FILLER_105_826 ();
 sg13g2_decap_8 FILLER_105_833 ();
 sg13g2_fill_1 FILLER_105_840 ();
endmodule
