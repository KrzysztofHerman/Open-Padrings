* NGSPICE file created from FMD_QNC_Padframe24.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for bondpad_70x70_novias abstract view
.subckt bondpad_70x70_novias pad
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_IOPadOut30mA abstract view
.subckt sg13g2_IOPadOut30mA c2p iovdd iovss pad vdd vss
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_Corner abstract view
.subckt sg13g2_Corner iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadVss abstract view
.subckt sg13g2_IOPadVss iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_IOPadIn abstract view
.subckt sg13g2_IOPadIn iovdd iovss p2c pad vdd vss
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_IOPadIOVss abstract view
.subckt sg13g2_IOPadIOVss iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadIOVdd abstract view
.subckt sg13g2_IOPadIOVdd iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadVdd abstract view
.subckt sg13g2_IOPadVdd iovdd iovss vdd vss
.ends

.subckt FMD_QNC_Padframe24 IOVDD IOVSS VDD VSS clk_PAD input_PAD[0] input_PAD[1] input_PAD[2]
+ input_PAD[3] input_PAD[4] input_PAD[5] input_PAD[6] input_PAD[7] output_PAD[0] output_PAD[1]
+ output_PAD[2] output_PAD[3] output_PAD[4] output_PAD[5] output_PAD[6] output_PAD[7]
+ output_PAD[8] output_PAD[9] rst_n_PAD
XFILLER_67_520 VDD VSS sg13g2_decap_8
XFILLER_94_350 VDD VSS sg13g2_decap_8
XFILLER_27_406 VDD VSS sg13g2_decap_8
XFILLER_39_266 VDD VSS sg13g2_decap_8
XFILLER_54_203 VDD VSS sg13g2_decap_8
XFILLER_67_597 VDD VSS sg13g2_decap_8
XFILLER_82_567 VDD VSS sg13g2_decap_8
XFILLER_70_729 VDD VSS sg13g2_decap_8
XFILLER_23_623 VDD VSS sg13g2_decap_8
XFILLER_35_483 VDD VSS sg13g2_decap_8
XFILLER_62_280 VDD VSS sg13g2_decap_8
XFILLER_22_133 VDD VSS sg13g2_decap_8
XFILLER_50_420 VDD VSS sg13g2_decap_8
XFILLER_50_497 VDD VSS sg13g2_decap_8
XFILLER_7_7 VDD VSS sg13g2_decap_8
XFILLER_89_133 VDD VSS sg13g2_decap_8
XFILLER_85_350 VDD VSS sg13g2_decap_8
XFILLER_93_14 VDD VSS sg13g2_decap_8
XFILLER_58_553 VDD VSS sg13g2_decap_8
XFILLER_18_406 VDD VSS sg13g2_decap_8
XFILLER_73_534 VDD VSS sg13g2_decap_8
XFILLER_45_203 VDD VSS sg13g2_decap_8
XFILLER_61_707 VDD VSS sg13g2_decap_8
XFILLER_26_63 VDD VSS sg13g2_decap_8
XFILLER_26_461 VDD VSS sg13g2_decap_8
XFILLER_60_217 VDD VSS sg13g2_decap_8
XFILLER_14_623 VDD VSS sg13g2_decap_8
XFILLER_13_133 VDD VSS sg13g2_decap_8
XFILLER_41_420 VDD VSS sg13g2_decap_8
XFILLER_53_280 VDD VSS sg13g2_decap_8
XFILLER_9_126 VDD VSS sg13g2_decap_8
XFILLER_41_497 VDD VSS sg13g2_decap_8
XFILLER_42_84 VDD VSS sg13g2_decap_8
XFILLER_5_343 VDD VSS sg13g2_decap_8
XFILLER_68_328 VDD VSS sg13g2_decap_8
XFILLER_1_560 VDD VSS sg13g2_decap_8
XFILLER_3_56 VDD VSS sg13g2_decap_8
XFILLER_95_147 VDD VSS sg13g2_decap_8
X_83_ _83__7/L_HI VSS VDD _83_/D _83_/Q _83_/CLK sg13g2_dfrbpq_1
XFILLER_67_70 VDD VSS sg13g2_decap_8
XFILLER_49_553 VDD VSS sg13g2_decap_8
XFILLER_76_383 VDD VSS sg13g2_decap_8
XFILLER_36_203 VDD VSS sg13g2_decap_8
XFILLER_64_567 VDD VSS sg13g2_decap_8
XFILLER_52_707 VDD VSS sg13g2_decap_8
XFILLER_91_364 VDD VSS sg13g2_decap_8
XFILLER_51_217 VDD VSS sg13g2_decap_8
XFILLER_17_483 VDD VSS sg13g2_decap_8
XFILLER_83_91 VDD VSS sg13g2_decap_8
XFILLER_32_420 VDD VSS sg13g2_decap_8
XFILLER_44_280 VDD VSS sg13g2_decap_8
XFILLER_20_637 VDD VSS sg13g2_decap_8
XFILLER_32_497 VDD VSS sg13g2_decap_8
XFILLER_66_0 VDD VSS sg13g2_decap_8
XFILLER_9_693 VDD VSS sg13g2_decap_8
XFILLER_87_637 VDD VSS sg13g2_decap_8
XFILLER_86_147 VDD VSS sg13g2_decap_8
XFILLER_74_309 VDD VSS sg13g2_decap_8
XFILLER_67_394 VDD VSS sg13g2_decap_8
XFILLER_27_203 VDD VSS sg13g2_decap_8
XFILLER_55_567 VDD VSS sg13g2_decap_8
XFILLER_43_707 VDD VSS sg13g2_decap_8
XFILLER_70_526 VDD VSS sg13g2_decap_8
XFILLER_82_364 VDD VSS sg13g2_decap_8
XFILLER_63_28 VDD VSS sg13g2_decap_8
XFILLER_42_217 VDD VSS sg13g2_decap_8
XFILLER_23_420 VDD VSS sg13g2_decap_8
XFILLER_35_280 VDD VSS sg13g2_decap_8
XFILLER_11_637 VDD VSS sg13g2_decap_8
XFILLER_50_294 VDD VSS sg13g2_decap_8
XFILLER_23_497 VDD VSS sg13g2_decap_8
XFILLER_10_147 VDD VSS sg13g2_decap_8
XFILLER_12_21 VDD VSS sg13g2_decap_8
XFILLER_88_14 VDD VSS sg13g2_decap_8
XFILLER_12_98 VDD VSS sg13g2_decap_8
XFILLER_2_357 VDD VSS sg13g2_decap_8
XFILLER_78_637 VDD VSS sg13g2_decap_8
XFILLER_77_147 VDD VSS sg13g2_decap_8
XFILLER_58_350 VDD VSS sg13g2_decap_8
XFILLER_18_203 VDD VSS sg13g2_decap_8
XFILLER_46_567 VDD VSS sg13g2_decap_8
XFILLER_37_84 VDD VSS sg13g2_decap_8
XFILLER_34_707 VDD VSS sg13g2_decap_8
XFILLER_73_386 VDD VSS sg13g2_fill_1
XFILLER_73_364 VDD VSS sg13g2_fill_1
XFILLER_61_504 VDD VSS sg13g2_decap_8
XFILLER_33_217 VDD VSS sg13g2_decap_8
XFILLER_14_420 VDD VSS sg13g2_decap_8
XFILLER_26_280 VDD VSS sg13g2_decap_8
XFILLER_14_497 VDD VSS sg13g2_decap_8
XFILLER_41_294 VDD VSS sg13g2_decap_8
XFILLER_6_630 VDD VSS sg13g2_decap_8
XFILLER_5_140 VDD VSS sg13g2_decap_8
XFILLER_69_615 VDD VSS sg13g2_decap_8
XFILLER_78_91 VDD VSS sg13g2_decap_8
XFILLER_68_147 VDD VSS sg13g2_decap_8
XFILLER_49_350 VDD VSS sg13g2_decap_8
XFILLER_77_681 VDD VSS sg13g2_decap_8
XFILLER_92_651 VDD VSS sg13g2_decap_8
X_66_ _66_/B _78_/Q _80_/Q _74_/D VDD VSS _66_/D sg13g2_nand4_1
XFILLER_25_707 VDD VSS sg13g2_decap_8
XFILLER_37_567 VDD VSS sg13g2_decap_8
XFILLER_91_161 VDD VSS sg13g2_decap_8
XFILLER_64_364 VDD VSS sg13g2_decap_8
XFILLER_52_504 VDD VSS sg13g2_decap_8
XFILLER_24_217 VDD VSS sg13g2_decap_8
XFILLER_17_280 VDD VSS sg13g2_decap_8
XFILLER_60_581 VDD VSS sg13g2_decap_8
XFILLER_20_434 VDD VSS sg13g2_decap_8
XFILLER_32_294 VDD VSS sg13g2_decap_8
XFILLER_9_490 VDD VSS sg13g2_decap_8
XFILLER_58_28 VDD VSS sg13g2_decap_8
XFILLER_87_434 VDD VSS sg13g2_decap_8
XFILLER_59_147 VDD VSS sg13g2_decap_8
XFILLER_68_692 VDD VSS sg13g2_decap_8
XFILLER_83_651 VDD VSS sg13g2_decap_8
XFILLER_74_49 VDD VSS sg13g2_decap_8
XFILLER_16_707 VDD VSS sg13g2_decap_8
XFILLER_28_567 VDD VSS sg13g2_decap_8
XFILLER_82_161 VDD VSS sg13g2_decap_8
XFILLER_15_217 VDD VSS sg13g2_decap_8
XFILLER_55_364 VDD VSS sg13g2_decap_8
XFILLER_43_504 VDD VSS sg13g2_decap_8
XFILLER_70_334 VDD VSS sg13g2_decap_8
XFILLER_51_581 VDD VSS sg13g2_decap_8
XFILLER_11_434 VDD VSS sg13g2_decap_8
XFILLER_23_42 VDD VSS sg13g2_decap_8
XFILLER_23_294 VDD VSS sg13g2_decap_8
XFILLER_7_427 VDD VSS sg13g2_decap_8
XFILLER_3_644 VDD VSS sg13g2_decap_8
XFILLER_2_154 VDD VSS sg13g2_decap_8
XFILLER_78_434 VDD VSS sg13g2_decap_8
XFILLER_66_618 VDD VSS sg13g2_decap_8
XFILLER_74_651 VDD VSS sg13g2_decap_8
XFILLER_93_448 VDD VSS sg13g2_decap_8
XFILLER_0_35 VDD VSS sg13g2_decap_8
XFILLER_73_161 VDD VSS sg13g2_decap_8
XFILLER_46_364 VDD VSS sg13g2_decap_8
XFILLER_61_301 VDD VSS sg13g2_decap_8
XFILLER_19_567 VDD VSS sg13g2_decap_8
XFILLER_34_504 VDD VSS sg13g2_decap_8
XFILLER_61_378 VDD VSS sg13g2_decap_8
XFILLER_30_721 VDD VSS sg13g2_decap_8
XFILLER_42_581 VDD VSS sg13g2_decap_8
XFILLER_9_77 VDD VSS sg13g2_decap_8
XFILLER_14_294 VDD VSS sg13g2_decap_8
XFILLER_80_70 VDD VSS sg13g2_decap_8
XFILLER_69_401 VDD VSS sg13g2_decap_8
XFILLER_69_456 VDD VSS sg13g2_fill_1
XFILLER_29_0 VDD VSS sg13g2_decap_8
XFILLER_65_640 VDD VSS sg13g2_decap_8
XFILLER_84_448 VDD VSS sg13g2_decap_8
X_49_ _51_/A _51_/B _52_/A _49_/Y VDD VSS _49_/D sg13g2_nand4_1
XFILLER_64_161 VDD VSS sg13g2_decap_8
XFILLER_37_364 VDD VSS sg13g2_decap_8
XFILLER_52_301 VDD VSS sg13g2_decap_8
XFILLER_25_504 VDD VSS sg13g2_decap_8
XFILLER_80_665 VDD VSS sg13g2_decap_8
XFILLER_52_378 VDD VSS sg13g2_decap_8
XFILLER_40_518 VDD VSS sg13g2_decap_8
XFILLER_21_721 VDD VSS sg13g2_decap_8
XFILLER_33_581 VDD VSS sg13g2_decap_8
XFILLER_20_231 VDD VSS sg13g2_decap_8
XFILLER_69_49 VDD VSS sg13g2_decap_8
XFILLER_88_721 VDD VSS sg13g2_decap_8
XFILLER_87_231 VDD VSS sg13g2_decap_8
XFILLER_0_658 VDD VSS sg13g2_decap_8
XFILLER_75_437 VDD VSS sg13g2_decap_8
XFILLER_56_651 VDD VSS sg13g2_decap_8
XFILLER_18_42 VDD VSS sg13g2_decap_8
XFILLER_28_364 VDD VSS sg13g2_decap_8
XFILLER_43_301 VDD VSS sg13g2_decap_8
XFILLER_55_161 VDD VSS sg13g2_decap_8
XFILLER_16_504 VDD VSS sg13g2_decap_8
XFILLER_71_632 VDD VSS sg13g2_decap_8
XFILLER_31_518 VDD VSS sg13g2_decap_8
XFILLER_70_175 VDD VSS sg13g2_decap_8
XFILLER_12_721 VDD VSS sg13g2_decap_8
XFILLER_34_63 VDD VSS sg13g2_decap_8
XFILLER_43_378 VDD VSS sg13g2_decap_8
XFILLER_24_581 VDD VSS sg13g2_decap_8
XFILLER_11_231 VDD VSS sg13g2_decap_8
XFILLER_8_714 VDD VSS sg13g2_decap_8
X_83__7 VDD VSS _83__7/L_HI sg13g2_tiehi
XFILLER_7_224 VDD VSS sg13g2_decap_8
XFILLER_50_84 VDD VSS sg13g2_decap_8
XFILLER_3_441 VDD VSS sg13g2_decap_8
XFILLER_79_721 VDD VSS sg13g2_decap_8
XFILLER_78_231 VDD VSS sg13g2_decap_8
XFILLER_22_7 VDD VSS sg13g2_decap_8
XFILLER_94_735 VDD VSS sg13g2_decap_8
XFILLER_93_245 VDD VSS sg13g2_decap_8
XFILLER_66_448 VDD VSS sg13g2_fill_2
XFILLER_75_81 VDD VSS sg13g2_decap_8
XFILLER_47_651 VDD VSS sg13g2_decap_8
XFILLER_19_364 VDD VSS sg13g2_decap_8
XFILLER_34_301 VDD VSS sg13g2_decap_8
XFILLER_46_161 VDD VSS sg13g2_decap_8
XFILLER_62_665 VDD VSS sg13g2_decap_8
XFILLER_34_378 VDD VSS sg13g2_decap_8
XFILLER_61_175 VDD VSS sg13g2_decap_8
XFILLER_15_581 VDD VSS sg13g2_decap_8
XFILLER_22_518 VDD VSS sg13g2_decap_8
XFILLER_91_91 VDD VSS sg13g2_decap_8
XFILLER_30_595 VDD VSS sg13g2_decap_8
XFILLER_89_518 VDD VSS sg13g2_decap_8
XFILLER_69_231 VDD VSS sg13g2_decap_8
XFILLER_85_735 VDD VSS sg13g2_decap_8
XFILLER_69_275 VDD VSS sg13g2_decap_8
XFILLER_84_245 VDD VSS sg13g2_decap_8
XFILLER_57_448 VDD VSS sg13g2_decap_8
XFILLER_38_651 VDD VSS sg13g2_decap_8
XFILLER_25_301 VDD VSS sg13g2_decap_8
XFILLER_37_161 VDD VSS sg13g2_decap_8
XFILLER_80_462 VDD VSS sg13g2_decap_8
XFILLER_53_665 VDD VSS sg13g2_decap_8
XFILLER_71_28 VDD VSS sg13g2_decap_8
XFILLER_13_518 VDD VSS sg13g2_decap_8
XFILLER_25_378 VDD VSS sg13g2_decap_8
XFILLER_40_315 VDD VSS sg13g2_decap_8
XFILLER_52_175 VDD VSS sg13g2_decap_8
XFILLER_21_595 VDD VSS sg13g2_decap_8
XFILLER_5_728 VDD VSS sg13g2_decap_8
XFILLER_4_238 VDD VSS sg13g2_decap_8
XFILLER_20_21 VDD VSS sg13g2_decap_8
XFILLER_20_98 VDD VSS sg13g2_decap_8
XFILLER_0_455 VDD VSS sg13g2_decap_8
XFILLER_88_595 VDD VSS sg13g2_decap_8
XFILLER_76_713 VDD VSS sg13g2_decap_8
Xhold30 _66_/D VDD VSS _58_/C sg13g2_dlygate4sd3_1
XFILLER_29_63 VDD VSS sg13g2_decap_8
XFILLER_48_448 VDD VSS sg13g2_decap_8
XFILLER_75_278 VDD VSS sg13g2_decap_4
XFILLER_29_651 VDD VSS sg13g2_decap_8
XFILLER_91_749 VDD VSS sg13g2_decap_8
XFILLER_16_301 VDD VSS sg13g2_decap_8
XFILLER_28_161 VDD VSS sg13g2_decap_8
XFILLER_90_259 VDD VSS sg13g2_decap_8
XFILLER_44_665 VDD VSS sg13g2_decap_8
XFILLER_45_84 VDD VSS sg13g2_decap_8
XFILLER_16_378 VDD VSS sg13g2_decap_8
XFILLER_31_315 VDD VSS sg13g2_decap_8
XFILLER_43_175 VDD VSS sg13g2_decap_8
XFILLER_8_511 VDD VSS sg13g2_decap_8
XFILLER_12_595 VDD VSS sg13g2_decap_8
XFILLER_8_588 VDD VSS sg13g2_decap_8
XFILLER_6_56 VDD VSS sg13g2_decap_8
XFILLER_79_595 VDD VSS sg13g2_decap_8
XFILLER_67_702 VDD VSS sg13g2_decap_8
XFILLER_94_532 VDD VSS sg13g2_decap_8
XFILLER_66_245 VDD VSS sg13g2_decap_8
XFILLER_86_91 VDD VSS sg13g2_decap_8
XFILLER_39_448 VDD VSS sg13g2_decap_8
XFILLER_82_749 VDD VSS sg13g2_decap_8
XFILLER_19_161 VDD VSS sg13g2_decap_8
XFILLER_81_259 VDD VSS sg13g2_decap_8
XFILLER_35_665 VDD VSS sg13g2_decap_8
XFILLER_62_462 VDD VSS sg13g2_decap_8
XFILLER_50_602 VDD VSS sg13g2_decap_8
XFILLER_22_315 VDD VSS sg13g2_decap_8
XFILLER_34_175 VDD VSS sg13g2_decap_8
XFILLER_50_679 VDD VSS sg13g2_decap_8
XFILLER_30_392 VDD VSS sg13g2_decap_8
XFILLER_89_315 VDD VSS sg13g2_decap_8
XFILLER_58_735 VDD VSS sg13g2_decap_8
XFILLER_85_532 VDD VSS sg13g2_decap_8
XFILLER_66_28 VDD VSS sg13g2_decap_8
XFILLER_57_245 VDD VSS sg13g2_decap_8
XFILLER_73_716 VDD VSS sg13g2_decap_8
XFILLER_26_643 VDD VSS sg13g2_decap_8
XFILLER_82_49 VDD VSS sg13g2_decap_8
XFILLER_13_315 VDD VSS sg13g2_decap_8
XFILLER_15_21 VDD VSS sg13g2_decap_8
XFILLER_25_175 VDD VSS sg13g2_decap_8
XFILLER_53_462 VDD VSS sg13g2_decap_8
XFILLER_41_602 VDD VSS sg13g2_decap_8
XFILLER_40_112 VDD VSS sg13g2_decap_8
XFILLER_9_308 VDD VSS sg13g2_decap_8
XFILLER_15_98 VDD VSS sg13g2_decap_8
XFILLER_41_679 VDD VSS sg13g2_decap_8
XFILLER_40_189 VDD VSS sg13g2_decap_8
XFILLER_31_42 VDD VSS sg13g2_decap_8
XFILLER_21_392 VDD VSS sg13g2_decap_8
XFILLER_5_525 VDD VSS sg13g2_decap_8
XFILLER_1_742 VDD VSS sg13g2_decap_8
XFILLER_76_510 VDD VSS sg13g2_decap_8
XFILLER_95_329 VDD VSS sg13g2_decap_8
XFILLER_0_252 VDD VSS sg13g2_decap_8
XFILLER_88_392 VDD VSS sg13g2_decap_8
XFILLER_49_735 VDD VSS sg13g2_decap_8
XFILLER_76_587 VDD VSS sg13g2_decap_8
XFILLER_48_245 VDD VSS sg13g2_decap_8
XFILLER_91_546 VDD VSS sg13g2_decap_8
XFILLER_64_749 VDD VSS sg13g2_decap_8
XFILLER_63_259 VDD VSS sg13g2_decap_8
XFILLER_17_665 VDD VSS sg13g2_decap_8
XFILLER_16_175 VDD VSS sg13g2_decap_8
XFILLER_44_462 VDD VSS sg13g2_decap_8
XFILLER_32_602 VDD VSS sg13g2_decap_8
XFILLER_71_270 VDD VSS sg13g2_decap_8
XFILLER_31_112 VDD VSS sg13g2_decap_8
XFILLER_32_679 VDD VSS sg13g2_decap_8
XFILLER_31_189 VDD VSS sg13g2_decap_8
XFILLER_12_392 VDD VSS sg13g2_decap_8
XFILLER_8_385 VDD VSS sg13g2_decap_8
XFILLER_86_329 VDD VSS sg13g2_decap_8
XFILLER_79_392 VDD VSS sg13g2_decap_8
XFILLER_67_576 VDD VSS sg13g2_decap_8
XFILLER_11_0 VDD VSS sg13g2_decap_8
XFILLER_39_245 VDD VSS sg13g2_decap_8
XFILLER_55_749 VDD VSS sg13g2_decap_8
XFILLER_82_546 VDD VSS sg13g2_decap_8
XFILLER_70_708 VDD VSS sg13g2_decap_8
XFILLER_54_259 VDD VSS sg13g2_decap_8
XFILLER_35_462 VDD VSS sg13g2_decap_8
XFILLER_23_602 VDD VSS sg13g2_decap_8
XFILLER_22_112 VDD VSS sg13g2_decap_8
XFILLER_50_476 VDD VSS sg13g2_decap_8
XFILLER_23_679 VDD VSS sg13g2_decap_8
XFILLER_10_329 VDD VSS sg13g2_decap_8
XFILLER_22_189 VDD VSS sg13g2_decap_8
XFILLER_89_112 VDD VSS sg13g2_decap_8
XFILLER_2_539 VDD VSS sg13g2_decap_8
XFILLER_89_189 VDD VSS sg13g2_decap_8
XFILLER_77_49 VDD VSS sg13g2_decap_8
XFILLER_58_532 VDD VSS sg13g2_decap_8
XFILLER_73_513 VDD VSS sg13g2_decap_8
XFILLER_46_749 VDD VSS sg13g2_decap_8
XFILLER_26_42 VDD VSS sg13g2_decap_8
XFILLER_26_440 VDD VSS sg13g2_decap_8
XFILLER_45_259 VDD VSS sg13g2_decap_8
XFILLER_14_602 VDD VSS sg13g2_decap_8
XFILLER_13_112 VDD VSS sg13g2_decap_8
XFILLER_9_105 VDD VSS sg13g2_decap_8
XFILLER_41_476 VDD VSS sg13g2_decap_8
XFILLER_14_679 VDD VSS sg13g2_decap_8
XFILLER_13_189 VDD VSS sg13g2_decap_8
XFILLER_42_63 VDD VSS sg13g2_decap_8
XFILLER_5_322 VDD VSS sg13g2_decap_8
XFILLER_5_399 VDD VSS sg13g2_decap_8
XFILLER_68_307 VDD VSS sg13g2_decap_8
XFILLER_3_35 VDD VSS sg13g2_decap_8
XFILLER_95_126 VDD VSS sg13g2_decap_8
XFILLER_49_532 VDD VSS sg13g2_decap_8
X_82_ _82__5/L_HI VSS VDD _82_/D _82_/Q _83_/CLK sg13g2_dfrbpq_1
XFILLER_76_362 VDD VSS sg13g2_decap_8
XFILLER_37_749 VDD VSS sg13g2_decap_8
XFILLER_64_546 VDD VSS sg13g2_decap_8
XFILLER_91_343 VDD VSS sg13g2_decap_8
XFILLER_36_259 VDD VSS sg13g2_decap_8
XFILLER_83_70 VDD VSS sg13g2_decap_8
XFILLER_17_462 VDD VSS sg13g2_decap_8
XFILLER_20_616 VDD VSS sg13g2_decap_8
XFILLER_32_476 VDD VSS sg13g2_decap_8
XFILLER_9_672 VDD VSS sg13g2_decap_8
XFILLER_8_182 VDD VSS sg13g2_decap_8
XFILLER_59_0 VDD VSS sg13g2_decap_8
XFILLER_87_616 VDD VSS sg13g2_decap_8
XFILLER_86_126 VDD VSS sg13g2_decap_8
XFILLER_59_329 VDD VSS sg13g2_decap_8
XFILLER_95_693 VDD VSS sg13g2_decap_8
XFILLER_67_373 VDD VSS sg13g2_decap_8
XFILLER_28_749 VDD VSS sg13g2_decap_8
XFILLER_82_343 VDD VSS sg13g2_decap_8
XFILLER_55_546 VDD VSS sg13g2_decap_8
XFILLER_27_259 VDD VSS sg13g2_decap_8
XFILLER_70_505 VDD VSS sg13g2_decap_8
XFILLER_11_616 VDD VSS sg13g2_decap_8
XFILLER_23_476 VDD VSS sg13g2_decap_8
XFILLER_50_273 VDD VSS sg13g2_decap_8
XFILLER_7_609 VDD VSS sg13g2_decap_8
XFILLER_10_126 VDD VSS sg13g2_decap_8
XFILLER_6_119 VDD VSS sg13g2_decap_8
XFILLER_12_77 VDD VSS sg13g2_decap_8
XFILLER_2_336 VDD VSS sg13g2_decap_8
XFILLER_78_616 VDD VSS sg13g2_decap_8
XFILLER_77_126 VDD VSS sg13g2_decap_8
XFILLER_86_693 VDD VSS sg13g2_decap_8
XFILLER_19_749 VDD VSS sg13g2_decap_8
XFILLER_73_332 VDD VSS sg13g2_decap_8
XFILLER_73_343 VDD VSS sg13g2_fill_2
XFILLER_46_546 VDD VSS sg13g2_decap_8
XFILLER_37_63 VDD VSS sg13g2_decap_8
XFILLER_18_259 VDD VSS sg13g2_decap_8
XFILLER_53_84 VDD VSS sg13g2_decap_8
XFILLER_14_476 VDD VSS sg13g2_decap_8
XFILLER_41_273 VDD VSS sg13g2_decap_8
XFILLER_10_693 VDD VSS sg13g2_decap_8
XFILLER_6_686 VDD VSS sg13g2_decap_8
XFILLER_52_7 VDD VSS sg13g2_decap_8
XFILLER_5_196 VDD VSS sg13g2_decap_8
XFILLER_68_126 VDD VSS sg13g2_decap_8
XFILLER_78_70 VDD VSS sg13g2_decap_8
XFILLER_77_660 VDD VSS sg13g2_decap_8
XFILLER_92_630 VDD VSS sg13g2_decap_8
X_65_ _65_/Y _65_/B hold23/X VDD VSS sg13g2_nand2b_1
XFILLER_64_343 VDD VSS sg13g2_decap_8
XFILLER_37_546 VDD VSS sg13g2_decap_8
XFILLER_91_140 VDD VSS sg13g2_decap_8
XFILLER_94_91 VDD VSS sg13g2_decap_8
XFILLER_60_560 VDD VSS sg13g2_decap_8
XFILLER_20_413 VDD VSS sg13g2_decap_8
XFILLER_32_273 VDD VSS sg13g2_decap_8
XFILLER_87_413 VDD VSS sg13g2_decap_8
XFILLER_59_126 VDD VSS sg13g2_decap_8
XFILLER_68_671 VDD VSS sg13g2_decap_8
XFILLER_95_490 VDD VSS sg13g2_decap_8
XFILLER_83_630 VDD VSS sg13g2_decap_8
XFILLER_74_28 VDD VSS sg13g2_decap_8
XFILLER_55_343 VDD VSS sg13g2_decap_8
XFILLER_28_546 VDD VSS sg13g2_decap_8
XFILLER_82_140 VDD VSS sg13g2_decap_8
XFILLER_70_313 VDD VSS sg13g2_decap_8
XFILLER_90_49 VDD VSS sg13g2_decap_8
XFILLER_51_560 VDD VSS sg13g2_decap_8
XFILLER_11_413 VDD VSS sg13g2_decap_8
XFILLER_23_21 VDD VSS sg13g2_decap_8
XFILLER_23_273 VDD VSS sg13g2_decap_8
XFILLER_7_406 VDD VSS sg13g2_decap_8
XFILLER_23_98 VDD VSS sg13g2_decap_8
XFILLER_3_623 VDD VSS sg13g2_decap_8
XFILLER_2_133 VDD VSS sg13g2_decap_8
XFILLER_78_413 VDD VSS sg13g2_decap_8
XFILLER_93_427 VDD VSS sg13g2_decap_8
XFILLER_48_84 VDD VSS sg13g2_decap_8
XFILLER_86_490 VDD VSS sg13g2_decap_8
XFILLER_74_630 VDD VSS sg13g2_decap_8
XFILLER_59_693 VDD VSS sg13g2_decap_8
XFILLER_0_14 VDD VSS sg13g2_decap_8
XFILLER_46_343 VDD VSS sg13g2_decap_8
XFILLER_19_546 VDD VSS sg13g2_decap_8
XFILLER_73_140 VDD VSS sg13g2_decap_8
XFILLER_61_357 VDD VSS sg13g2_decap_8
XFILLER_14_273 VDD VSS sg13g2_decap_8
XFILLER_30_700 VDD VSS sg13g2_decap_8
XFILLER_42_560 VDD VSS sg13g2_decap_8
XFILLER_9_56 VDD VSS sg13g2_decap_8
XFILLER_10_490 VDD VSS sg13g2_decap_8
XFILLER_6_483 VDD VSS sg13g2_decap_8
XFILLER_89_91 VDD VSS sg13g2_decap_8
XFILLER_84_427 VDD VSS sg13g2_decap_8
X_48_ _52_/C _52_/D _51_/C _60_/B VDD VSS _51_/D sg13g2_nand4_1
XFILLER_64_140 VDD VSS sg13g2_decap_8
XFILLER_37_343 VDD VSS sg13g2_decap_8
XFILLER_80_644 VDD VSS sg13g2_decap_8
XFILLER_65_696 VDD VSS sg13g2_decap_8
XFILLER_52_357 VDD VSS sg13g2_decap_8
XFILLER_21_700 VDD VSS sg13g2_decap_8
XFILLER_33_560 VDD VSS sg13g2_decap_8
XFILLER_20_210 VDD VSS sg13g2_decap_8
XFILLER_20_287 VDD VSS sg13g2_decap_8
XFILLER_69_28 VDD VSS sg13g2_decap_8
XFILLER_88_700 VDD VSS sg13g2_decap_8
XFILLER_87_210 VDD VSS sg13g2_decap_8
XFILLER_0_637 VDD VSS sg13g2_decap_8
XFILLER_87_287 VDD VSS sg13g2_decap_8
XFILLER_75_416 VDD VSS sg13g2_decap_8
XFILLER_85_49 VDD VSS sg13g2_decap_8
XFILLER_56_630 VDD VSS sg13g2_decap_8
XFILLER_18_21 VDD VSS sg13g2_decap_8
XFILLER_28_343 VDD VSS sg13g2_decap_8
XFILLER_55_140 VDD VSS sg13g2_decap_8
XFILLER_71_611 VDD VSS sg13g2_decap_8
XFILLER_18_98 VDD VSS sg13g2_decap_8
XFILLER_70_154 VDD VSS sg13g2_decap_8
XFILLER_43_357 VDD VSS sg13g2_decap_8
XFILLER_71_688 VDD VSS sg13g2_decap_8
XFILLER_12_700 VDD VSS sg13g2_decap_8
XFILLER_34_42 VDD VSS sg13g2_decap_8
XFILLER_24_560 VDD VSS sg13g2_decap_8
XFILLER_11_210 VDD VSS sg13g2_decap_8
XFILLER_7_203 VDD VSS sg13g2_decap_8
XFILLER_11_287 VDD VSS sg13g2_decap_8
XFILLER_50_63 VDD VSS sg13g2_decap_8
XFILLER_3_420 VDD VSS sg13g2_decap_8
XFILLER_79_700 VDD VSS sg13g2_decap_8
XFILLER_78_210 VDD VSS sg13g2_decap_8
XFILLER_3_497 VDD VSS sg13g2_decap_8
XFILLER_94_714 VDD VSS sg13g2_decap_8
XFILLER_78_287 VDD VSS sg13g2_decap_8
XFILLER_66_427 VDD VSS sg13g2_decap_8
XFILLER_93_224 VDD VSS sg13g2_decap_8
XFILLER_59_490 VDD VSS sg13g2_decap_8
XFILLER_47_630 VDD VSS sg13g2_decap_8
XFILLER_15_7 VDD VSS sg13g2_decap_8
XFILLER_75_60 VDD VSS sg13g2_decap_8
XFILLER_19_343 VDD VSS sg13g2_decap_8
XFILLER_46_140 VDD VSS sg13g2_decap_8
XFILLER_62_644 VDD VSS sg13g2_decap_8
XFILLER_34_357 VDD VSS sg13g2_decap_8
XFILLER_61_154 VDD VSS sg13g2_decap_8
XFILLER_15_560 VDD VSS sg13g2_decap_8
XFILLER_91_70 VDD VSS sg13g2_decap_8
XFILLER_30_574 VDD VSS sg13g2_decap_8
XFILLER_6_280 VDD VSS sg13g2_decap_8
XFILLER_69_210 VDD VSS sg13g2_decap_8
XFILLER_41_0 VDD VSS sg13g2_decap_8
XFILLER_85_714 VDD VSS sg13g2_decap_8
XFILLER_69_254 VDD VSS sg13g2_decap_8
XFILLER_57_427 VDD VSS sg13g2_decap_8
XFILLER_84_224 VDD VSS sg13g2_decap_8
XFILLER_38_630 VDD VSS sg13g2_decap_8
XFILLER_37_140 VDD VSS sg13g2_decap_8
XFILLER_65_493 VDD VSS sg13g2_decap_8
XFILLER_65_471 VDD VSS sg13g2_fill_1
XFILLER_80_441 VDD VSS sg13g2_decap_8
XFILLER_53_644 VDD VSS sg13g2_decap_8
XFILLER_25_357 VDD VSS sg13g2_decap_8
XFILLER_52_154 VDD VSS sg13g2_decap_8
XFILLER_21_574 VDD VSS sg13g2_decap_8
XFILLER_5_707 VDD VSS sg13g2_decap_8
XFILLER_4_217 VDD VSS sg13g2_decap_8
XFILLER_20_77 VDD VSS sg13g2_decap_8
XFILLER_0_434 VDD VSS sg13g2_decap_8
XFILLER_88_574 VDD VSS sg13g2_decap_8
Xhold20 _81_/Q VDD VSS _45_/A sg13g2_dlygate4sd3_1
Xhold31 _58_/Y VDD VSS _77_/D sg13g2_dlygate4sd3_1
XFILLER_29_42 VDD VSS sg13g2_decap_8
XFILLER_48_427 VDD VSS sg13g2_decap_8
XFILLER_75_235 VDD VSS sg13g2_fill_2
XFILLER_29_630 VDD VSS sg13g2_decap_8
XFILLER_91_728 VDD VSS sg13g2_decap_8
XFILLER_75_257 VDD VSS sg13g2_decap_8
XFILLER_28_140 VDD VSS sg13g2_decap_8
XFILLER_90_238 VDD VSS sg13g2_decap_8
X_78__8 VDD VSS _78__8/L_HI sg13g2_tiehi
XFILLER_45_63 VDD VSS sg13g2_decap_8
XFILLER_16_357 VDD VSS sg13g2_decap_8
XFILLER_44_644 VDD VSS sg13g2_decap_8
XFILLER_71_485 VDD VSS sg13g2_decap_8
XFILLER_43_154 VDD VSS sg13g2_decap_8
XFILLER_12_574 VDD VSS sg13g2_decap_8
XFILLER_61_84 VDD VSS sg13g2_decap_8
XFILLER_8_567 VDD VSS sg13g2_decap_8
XFILLER_6_35 VDD VSS sg13g2_decap_8
XFILLER_3_294 VDD VSS sg13g2_decap_8
XFILLER_94_511 VDD VSS sg13g2_decap_8
XFILLER_79_574 VDD VSS sg13g2_decap_8
XFILLER_66_224 VDD VSS sg13g2_decap_8
XFILLER_86_70 VDD VSS sg13g2_decap_8
XFILLER_39_427 VDD VSS sg13g2_decap_8
XFILLER_94_588 VDD VSS sg13g2_decap_8
XFILLER_82_728 VDD VSS sg13g2_decap_8
XFILLER_19_140 VDD VSS sg13g2_decap_8
XFILLER_81_238 VDD VSS sg13g2_decap_8
XFILLER_62_441 VDD VSS sg13g2_decap_8
XFILLER_35_644 VDD VSS sg13g2_decap_8
XFILLER_34_154 VDD VSS sg13g2_decap_8
XFILLER_50_658 VDD VSS sg13g2_decap_8
XFILLER_89_0 VDD VSS sg13g2_decap_8
XFILLER_30_371 VDD VSS sg13g2_decap_8
XFILLER_85_511 VDD VSS sg13g2_decap_8
XFILLER_58_714 VDD VSS sg13g2_decap_8
XFILLER_57_224 VDD VSS sg13g2_decap_8
XFILLER_85_588 VDD VSS sg13g2_decap_8
XFILLER_26_622 VDD VSS sg13g2_decap_8
XFILLER_72_249 VDD VSS sg13g2_decap_8
XFILLER_82_28 VDD VSS sg13g2_decap_8
XFILLER_53_441 VDD VSS sg13g2_decap_8
XFILLER_25_154 VDD VSS sg13g2_decap_8
XFILLER_26_699 VDD VSS sg13g2_decap_8
XFILLER_41_658 VDD VSS sg13g2_decap_8
XFILLER_15_77 VDD VSS sg13g2_decap_8
XFILLER_40_168 VDD VSS sg13g2_decap_8
XFILLER_21_371 VDD VSS sg13g2_decap_8
XFILLER_5_504 VDD VSS sg13g2_decap_8
XFILLER_31_21 VDD VSS sg13g2_decap_8
XFILLER_31_98 VDD VSS sg13g2_decap_8
XFILLER_1_721 VDD VSS sg13g2_decap_8
XFILLER_95_308 VDD VSS sg13g2_decap_8
XFILLER_49_714 VDD VSS sg13g2_decap_8
XFILLER_0_231 VDD VSS sg13g2_decap_8
XFILLER_88_371 VDD VSS sg13g2_decap_8
XFILLER_48_224 VDD VSS sg13g2_decap_8
XFILLER_76_566 VDD VSS sg13g2_decap_8
XFILLER_91_525 VDD VSS sg13g2_decap_8
XFILLER_64_728 VDD VSS sg13g2_decap_8
XFILLER_56_84 VDD VSS sg13g2_decap_8
XFILLER_63_238 VDD VSS sg13g2_decap_8
XFILLER_44_441 VDD VSS sg13g2_decap_8
XFILLER_17_644 VDD VSS sg13g2_decap_8
XFILLER_16_154 VDD VSS sg13g2_decap_8
XFILLER_32_658 VDD VSS sg13g2_decap_8
XFILLER_31_168 VDD VSS sg13g2_decap_8
XFILLER_82_7 VDD VSS sg13g2_decap_8
XFILLER_12_371 VDD VSS sg13g2_decap_8
XFILLER_8_364 VDD VSS sg13g2_decap_8
XFILLER_4_581 VDD VSS sg13g2_decap_8
XFILLER_86_308 VDD VSS sg13g2_decap_8
XFILLER_79_371 VDD VSS sg13g2_decap_8
XFILLER_39_224 VDD VSS sg13g2_decap_8
XFILLER_67_555 VDD VSS sg13g2_decap_8
XFILLER_82_525 VDD VSS sg13g2_decap_8
XFILLER_94_385 VDD VSS sg13g2_decap_8
XFILLER_55_728 VDD VSS sg13g2_decap_8
XFILLER_35_441 VDD VSS sg13g2_decap_8
XFILLER_54_238 VDD VSS sg13g2_decap_8
XFILLER_10_308 VDD VSS sg13g2_decap_8
XFILLER_50_455 VDD VSS sg13g2_decap_8
XFILLER_23_658 VDD VSS sg13g2_decap_8
XFILLER_22_168 VDD VSS sg13g2_decap_8
XFILLER_2_518 VDD VSS sg13g2_decap_8
XFILLER_77_28 VDD VSS sg13g2_decap_8
XFILLER_89_168 VDD VSS sg13g2_decap_8
XFILLER_58_511 VDD VSS sg13g2_decap_8
XFILLER_85_385 VDD VSS sg13g2_decap_8
XFILLER_58_588 VDD VSS sg13g2_decap_8
XFILLER_46_728 VDD VSS sg13g2_decap_8
XFILLER_73_569 VDD VSS sg13g2_decap_8
XFILLER_93_49 VDD VSS sg13g2_decap_8
XFILLER_26_21 VDD VSS sg13g2_decap_8
XFILLER_45_238 VDD VSS sg13g2_decap_8
XFILLER_26_98 VDD VSS sg13g2_decap_8
XFILLER_26_496 VDD VSS sg13g2_decap_8
XFILLER_41_455 VDD VSS sg13g2_decap_8
XFILLER_14_658 VDD VSS sg13g2_decap_8
XFILLER_13_168 VDD VSS sg13g2_decap_8
XFILLER_42_42 VDD VSS sg13g2_decap_8
XFILLER_5_301 VDD VSS sg13g2_decap_8
XFILLER_5_378 VDD VSS sg13g2_decap_8
XFILLER_95_105 VDD VSS sg13g2_decap_8
XFILLER_3_14 VDD VSS sg13g2_decap_8
XFILLER_49_511 VDD VSS sg13g2_decap_8
XFILLER_1_595 VDD VSS sg13g2_decap_8
X_81_ _81__9/L_HI VSS VDD _81_/D _81_/Q _83_/CLK sg13g2_dfrbpq_1
XFILLER_76_341 VDD VSS sg13g2_decap_8
XFILLER_64_525 VDD VSS sg13g2_decap_8
XFILLER_49_588 VDD VSS sg13g2_decap_8
XFILLER_37_728 VDD VSS sg13g2_decap_8
XFILLER_91_322 VDD VSS sg13g2_decap_8
XFILLER_36_238 VDD VSS sg13g2_decap_8
XFILLER_17_441 VDD VSS sg13g2_decap_8
XFILLER_91_399 VDD VSS sg13g2_decap_8
XFILLER_60_742 VDD VSS sg13g2_decap_8
XFILLER_32_455 VDD VSS sg13g2_decap_8
XFILLER_9_651 VDD VSS sg13g2_decap_8
XFILLER_8_161 VDD VSS sg13g2_decap_8
XFILLER_86_105 VDD VSS sg13g2_decap_8
XFILLER_59_308 VDD VSS sg13g2_decap_8
XFILLER_67_352 VDD VSS sg13g2_decap_8
XFILLER_95_672 VDD VSS sg13g2_decap_8
XFILLER_55_525 VDD VSS sg13g2_decap_8
XFILLER_28_728 VDD VSS sg13g2_decap_8
XFILLER_94_182 VDD VSS sg13g2_decap_8
XFILLER_82_322 VDD VSS sg13g2_decap_8
XFILLER_27_238 VDD VSS sg13g2_decap_8
XFILLER_82_399 VDD VSS sg13g2_decap_8
XFILLER_51_742 VDD VSS sg13g2_decap_8
XFILLER_23_455 VDD VSS sg13g2_decap_8
XIO_BOND_outputs\[4\].output_pad output_PAD[4] bondpad_70x70_novias
XFILLER_10_105 VDD VSS sg13g2_decap_8
XFILLER_50_252 VDD VSS sg13g2_decap_8
XFILLER_12_56 VDD VSS sg13g2_decap_8
XFILLER_88_49 VDD VSS sg13g2_decap_8
XFILLER_2_315 VDD VSS sg13g2_decap_8
XFILLER_77_105 VDD VSS sg13g2_decap_8
XFILLER_93_609 VDD VSS sg13g2_decap_8
XFILLER_86_672 VDD VSS sg13g2_decap_8
XFILLER_92_119 VDD VSS sg13g2_decap_8
XFILLER_73_311 VDD VSS sg13g2_decap_8
XFILLER_46_525 VDD VSS sg13g2_decap_8
XFILLER_37_42 VDD VSS sg13g2_decap_8
XFILLER_58_385 VDD VSS sg13g2_decap_8
XFILLER_19_728 VDD VSS sg13g2_decap_8
XFILLER_85_182 VDD VSS sg13g2_decap_8
XFILLER_18_238 VDD VSS sg13g2_decap_8
XFILLER_61_539 VDD VSS sg13g2_decap_8
XFILLER_53_63 VDD VSS sg13g2_decap_8
XFILLER_14_455 VDD VSS sg13g2_decap_8
XFILLER_42_742 VDD VSS sg13g2_decap_8
XFILLER_41_252 VDD VSS sg13g2_decap_8
XFILLER_10_672 VDD VSS sg13g2_decap_8
XFILLER_6_665 VDD VSS sg13g2_decap_8
XFILLER_5_175 VDD VSS sg13g2_decap_8
XFILLER_45_7 VDD VSS sg13g2_decap_8
XFILLER_68_105 VDD VSS sg13g2_decap_8
XFILLER_84_609 VDD VSS sg13g2_decap_8
XFILLER_1_392 VDD VSS sg13g2_decap_8
XFILLER_83_119 VDD VSS sg13g2_decap_8
X_64_ _64_/A _65_/B _64_/Y VDD VSS sg13g2_nor2b_1
XFILLER_37_525 VDD VSS sg13g2_decap_8
XFILLER_76_182 VDD VSS sg13g2_decap_8
XFILLER_64_322 VDD VSS sg13g2_decap_8
XFILLER_94_70 VDD VSS sg13g2_decap_8
XFILLER_49_385 VDD VSS sg13g2_decap_8
XFILLER_92_686 VDD VSS sg13g2_decap_8
XFILLER_91_196 VDD VSS sg13g2_decap_8
XFILLER_64_399 VDD VSS sg13g2_decap_8
XFILLER_52_539 VDD VSS sg13g2_decap_8
XFILLER_33_742 VDD VSS sg13g2_decap_8
XFILLER_32_252 VDD VSS sg13g2_decap_8
XFILLER_71_0 VDD VSS sg13g2_decap_8
XFILLER_20_469 VDD VSS sg13g2_decap_8
XFILLER_59_105 VDD VSS sg13g2_decap_8
XFILLER_68_650 VDD VSS sg13g2_decap_8
XFILLER_87_469 VDD VSS sg13g2_decap_8
XFILLER_74_119 VDD VSS sg13g2_decap_8
XFILLER_67_182 VDD VSS sg13g2_decap_8
XFILLER_55_322 VDD VSS sg13g2_decap_8
XFILLER_28_525 VDD VSS sg13g2_decap_8
XFILLER_83_686 VDD VSS sg13g2_decap_8
XFILLER_82_196 VDD VSS sg13g2_decap_8
XFILLER_55_399 VDD VSS sg13g2_decap_8
XFILLER_43_539 VDD VSS sg13g2_decap_8
XFILLER_70_369 VDD VSS sg13g2_decap_8
XFILLER_90_28 VDD VSS sg13g2_decap_8
XFILLER_24_742 VDD VSS sg13g2_decap_8
XFILLER_23_252 VDD VSS sg13g2_decap_8
XFILLER_11_469 VDD VSS sg13g2_decap_8
XFILLER_23_77 VDD VSS sg13g2_decap_8
XFILLER_3_602 VDD VSS sg13g2_decap_8
XFILLER_2_112 VDD VSS sg13g2_decap_8
XFILLER_3_679 VDD VSS sg13g2_decap_8
XFILLER_2_189 VDD VSS sg13g2_decap_8
XFILLER_78_469 VDD VSS sg13g2_decap_8
XFILLER_93_406 VDD VSS sg13g2_decap_8
XFILLER_65_119 VDD VSS sg13g2_decap_8
XFILLER_59_672 VDD VSS sg13g2_decap_8
XFILLER_48_63 VDD VSS sg13g2_decap_8
XFILLER_46_322 VDD VSS sg13g2_decap_8
XFILLER_58_182 VDD VSS sg13g2_decap_8
XFILLER_19_525 VDD VSS sg13g2_decap_8
XFILLER_74_686 VDD VSS sg13g2_decap_8
XFILLER_46_399 VDD VSS sg13g2_decap_8
XFILLER_61_336 VDD VSS sg13g2_decap_8
XFILLER_34_539 VDD VSS sg13g2_decap_8
XFILLER_73_196 VDD VSS sg13g2_decap_8
XFILLER_64_84 VDD VSS sg13g2_decap_8
XFILLER_15_742 VDD VSS sg13g2_decap_8
XFILLER_9_35 VDD VSS sg13g2_decap_8
XFILLER_14_252 VDD VSS sg13g2_decap_8
XFILLER_30_756 VDD VSS sg13g2_fill_1
XFILLER_6_462 VDD VSS sg13g2_decap_8
XFILLER_89_70 VDD VSS sg13g2_decap_8
XFILLER_69_436 VDD VSS sg13g2_decap_8
XFILLER_57_609 VDD VSS sg13g2_decap_8
XFILLER_84_406 VDD VSS sg13g2_decap_8
XFILLER_56_119 VDD VSS sg13g2_decap_8
XFILLER_37_322 VDD VSS sg13g2_decap_8
XFILLER_49_182 VDD VSS sg13g2_decap_8
XFILLER_65_675 VDD VSS sg13g2_decap_8
X_47_ VDD _61_/A _75_/A VSS sg13g2_inv_1
XFILLER_92_483 VDD VSS sg13g2_decap_8
XFILLER_80_623 VDD VSS sg13g2_decap_8
XFILLER_37_399 VDD VSS sg13g2_decap_8
XFILLER_25_539 VDD VSS sg13g2_decap_8
XFILLER_64_196 VDD VSS sg13g2_decap_8
XFILLER_52_336 VDD VSS sg13g2_decap_8
XFILLER_21_756 VDD VSS sg13g2_fill_1
XFILLER_20_266 VDD VSS sg13g2_decap_8
XFILLER_0_616 VDD VSS sg13g2_decap_8
XFILLER_88_756 VDD VSS sg13g2_fill_1
XFILLER_48_609 VDD VSS sg13g2_decap_8
XFILLER_87_266 VDD VSS sg13g2_decap_8
XFILLER_85_28 VDD VSS sg13g2_decap_8
XFILLER_47_119 VDD VSS sg13g2_decap_8
XFILLER_28_322 VDD VSS sg13g2_decap_8
XFILLER_18_77 VDD VSS sg13g2_decap_8
XFILLER_83_483 VDD VSS sg13g2_decap_8
XFILLER_56_686 VDD VSS sg13g2_decap_8
XFILLER_28_399 VDD VSS sg13g2_decap_8
XFILLER_16_539 VDD VSS sg13g2_decap_8
XFILLER_71_667 VDD VSS sg13g2_decap_8
XFILLER_70_133 VDD VSS sg13g2_decap_8
XFILLER_34_21 VDD VSS sg13g2_decap_8
XFILLER_43_336 VDD VSS sg13g2_decap_8
XFILLER_55_196 VDD VSS sg13g2_decap_8
XFILLER_12_756 VDD VSS sg13g2_fill_1
XFILLER_34_98 VDD VSS sg13g2_decap_8
XFILLER_11_266 VDD VSS sg13g2_decap_8
XFILLER_8_749 VDD VSS sg13g2_decap_8
XFILLER_50_42 VDD VSS sg13g2_decap_8
XFILLER_7_259 VDD VSS sg13g2_decap_8
XFILLER_3_476 VDD VSS sg13g2_decap_8
XFILLER_1_0 VDD VSS sg13g2_decap_8
XFILLER_79_756 VDD VSS sg13g2_fill_1
XFILLER_59_84 VDD VSS sg13g2_decap_8
XFILLER_39_609 VDD VSS sg13g2_decap_8
XFILLER_93_203 VDD VSS sg13g2_decap_8
XFILLER_78_266 VDD VSS sg13g2_decap_8
XFILLER_66_406 VDD VSS sg13g2_decap_8
XFILLER_38_119 VDD VSS sg13g2_decap_8
XFILLER_19_322 VDD VSS sg13g2_decap_8
XFILLER_74_483 VDD VSS sg13g2_decap_8
XFILLER_62_623 VDD VSS sg13g2_decap_8
XFILLER_47_686 VDD VSS sg13g2_decap_8
XFILLER_19_399 VDD VSS sg13g2_decap_8
XFILLER_34_336 VDD VSS sg13g2_decap_8
XFILLER_46_196 VDD VSS sg13g2_decap_8
XFILLER_61_133 VDD VSS sg13g2_decap_8
XFILLER_30_553 VDD VSS sg13g2_decap_8
XFILLER_34_0 VDD VSS sg13g2_decap_8
XFILLER_84_203 VDD VSS sg13g2_decap_8
XFILLER_57_406 VDD VSS sg13g2_decap_8
XFILLER_29_119 VDD VSS sg13g2_decap_8
XFILLER_72_409 VDD VSS sg13g2_decap_8
XFILLER_53_623 VDD VSS sg13g2_decap_8
XFILLER_1_91 VDD VSS sg13g2_decap_8
XFILLER_38_686 VDD VSS sg13g2_decap_8
XFILLER_92_280 VDD VSS sg13g2_decap_8
XFILLER_80_420 VDD VSS sg13g2_decap_8
XFILLER_25_336 VDD VSS sg13g2_decap_8
XFILLER_37_196 VDD VSS sg13g2_decap_8
XFILLER_52_133 VDD VSS sg13g2_decap_8
XFILLER_80_497 VDD VSS sg13g2_decap_8
XFILLER_21_553 VDD VSS sg13g2_decap_8
XFILLER_20_56 VDD VSS sg13g2_decap_8
XFILLER_0_413 VDD VSS sg13g2_decap_8
XFILLER_88_553 VDD VSS sg13g2_decap_8
Xhold21 _70_/Y VDD VSS _81_/D sg13g2_dlygate4sd3_1
XFILLER_29_21 VDD VSS sg13g2_decap_8
XFILLER_48_406 VDD VSS sg13g2_decap_8
XFILLER_76_748 VDD VSS sg13g2_decap_8
XFILLER_75_214 VDD VSS sg13g2_decap_8
XFILLER_91_707 VDD VSS sg13g2_decap_8
XFILLER_29_98 VDD VSS sg13g2_decap_8
XFILLER_90_217 VDD VSS sg13g2_decap_8
XFILLER_56_483 VDD VSS sg13g2_decap_8
XFILLER_29_686 VDD VSS sg13g2_decap_8
XFILLER_44_623 VDD VSS sg13g2_decap_8
XFILLER_83_280 VDD VSS sg13g2_decap_8
XFILLER_45_42 VDD VSS sg13g2_decap_8
XFILLER_16_336 VDD VSS sg13g2_decap_8
XFILLER_28_196 VDD VSS sg13g2_decap_8
XFILLER_43_133 VDD VSS sg13g2_decap_8
XFILLER_71_464 VDD VSS sg13g2_decap_8
XFILLER_12_553 VDD VSS sg13g2_decap_8
XFILLER_8_546 VDD VSS sg13g2_decap_8
XFILLER_61_63 VDD VSS sg13g2_decap_8
XFILLER_6_14 VDD VSS sg13g2_decap_8
XFILLER_3_273 VDD VSS sg13g2_decap_8
XFILLER_79_553 VDD VSS sg13g2_decap_8
XFILLER_39_406 VDD VSS sg13g2_decap_8
XFILLER_67_737 VDD VSS sg13g2_decap_8
XFILLER_66_203 VDD VSS sg13g2_decap_8
XFILLER_94_567 VDD VSS sg13g2_decap_8
XFILLER_82_707 VDD VSS sg13g2_decap_8
XFILLER_81_217 VDD VSS sg13g2_decap_8
XFILLER_47_483 VDD VSS sg13g2_decap_8
XFILLER_35_623 VDD VSS sg13g2_decap_8
XFILLER_62_420 VDD VSS sg13g2_decap_8
XFILLER_19_196 VDD VSS sg13g2_decap_8
XFILLER_34_133 VDD VSS sg13g2_decap_8
XFILLER_62_497 VDD VSS sg13g2_decap_8
XFILLER_50_637 VDD VSS sg13g2_decap_8
XFILLER_30_350 VDD VSS sg13g2_decap_8
XIO_BOND_outputs\[9\].output_pad output_PAD[9] bondpad_70x70_novias
XFILLER_57_203 VDD VSS sg13g2_decap_8
XFILLER_85_567 VDD VSS sg13g2_decap_8
XFILLER_72_217 VDD VSS sg13g2_decap_8
XFILLER_26_601 VDD VSS sg13g2_decap_8
XFILLER_38_483 VDD VSS sg13g2_decap_8
XFILLER_65_280 VDD VSS sg13g2_decap_8
XIO_BOND_inputs\[7\].input_pad input_PAD[7] bondpad_70x70_novias
XFILLER_25_133 VDD VSS sg13g2_decap_8
XFILLER_53_420 VDD VSS sg13g2_decap_8
XFILLER_26_678 VDD VSS sg13g2_decap_8
XFILLER_80_294 VDD VSS sg13g2_decap_8
XFILLER_53_497 VDD VSS sg13g2_decap_8
XFILLER_15_56 VDD VSS sg13g2_decap_8
XFILLER_41_637 VDD VSS sg13g2_decap_8
XFILLER_40_147 VDD VSS sg13g2_decap_8
XFILLER_21_350 VDD VSS sg13g2_decap_8
XFILLER_31_77 VDD VSS sg13g2_decap_8
XFILLER_1_700 VDD VSS sg13g2_decap_8
XFILLER_0_210 VDD VSS sg13g2_decap_8
XFILLER_88_350 VDD VSS sg13g2_decap_8
XFILLER_0_287 VDD VSS sg13g2_decap_8
XFILLER_48_203 VDD VSS sg13g2_decap_8
XFILLER_76_545 VDD VSS sg13g2_decap_8
XFILLER_64_707 VDD VSS sg13g2_decap_8
XFILLER_91_504 VDD VSS sg13g2_decap_8
XFILLER_63_217 VDD VSS sg13g2_decap_8
XFILLER_56_63 VDD VSS sg13g2_decap_8
XFILLER_72_740 VDD VSS sg13g2_decap_8
XFILLER_44_420 VDD VSS sg13g2_decap_8
XFILLER_56_280 VDD VSS sg13g2_decap_8
XFILLER_17_623 VDD VSS sg13g2_decap_8
XFILLER_29_483 VDD VSS sg13g2_decap_8
XFILLER_16_133 VDD VSS sg13g2_decap_8
XFILLER_32_637 VDD VSS sg13g2_decap_8
XFILLER_44_497 VDD VSS sg13g2_decap_8
XFILLER_72_84 VDD VSS sg13g2_decap_8
XFILLER_31_147 VDD VSS sg13g2_decap_8
XFILLER_12_350 VDD VSS sg13g2_decap_8
XFILLER_75_7 VDD VSS sg13g2_decap_8
XFILLER_8_343 VDD VSS sg13g2_decap_8
XFILLER_4_560 VDD VSS sg13g2_decap_8
XFILLER_79_350 VDD VSS sg13g2_decap_8
XFILLER_67_534 VDD VSS sg13g2_decap_8
XFILLER_39_203 VDD VSS sg13g2_decap_8
XFILLER_55_707 VDD VSS sg13g2_decap_8
XFILLER_82_504 VDD VSS sg13g2_decap_8
XFILLER_94_364 VDD VSS sg13g2_decap_8
XFILLER_54_217 VDD VSS sg13g2_decap_8
XFILLER_35_420 VDD VSS sg13g2_decap_8
XFILLER_47_280 VDD VSS sg13g2_decap_8
XFILLER_90_581 VDD VSS sg13g2_decap_8
XFILLER_50_434 VDD VSS sg13g2_decap_8
XFILLER_23_637 VDD VSS sg13g2_decap_8
XFILLER_35_497 VDD VSS sg13g2_decap_8
XFILLER_62_294 VDD VSS sg13g2_decap_8
XFILLER_22_147 VDD VSS sg13g2_decap_8
XFILLER_89_147 VDD VSS sg13g2_decap_8
XFILLER_77_309 VDD VSS sg13g2_decap_8
XFILLER_58_567 VDD VSS sg13g2_decap_8
XFILLER_46_707 VDD VSS sg13g2_decap_8
XFILLER_85_364 VDD VSS sg13g2_decap_8
XFILLER_93_28 VDD VSS sg13g2_decap_8
XFILLER_45_217 VDD VSS sg13g2_decap_8
XFILLER_73_548 VDD VSS sg13g2_decap_8
XFILLER_38_280 VDD VSS sg13g2_decap_8
XFILLER_81_581 VDD VSS sg13g2_decap_8
XFILLER_26_77 VDD VSS sg13g2_decap_8
XFILLER_26_475 VDD VSS sg13g2_decap_8
XFILLER_14_637 VDD VSS sg13g2_decap_8
XFILLER_13_147 VDD VSS sg13g2_decap_8
XFILLER_41_434 VDD VSS sg13g2_decap_8
XFILLER_53_294 VDD VSS sg13g2_decap_8
XFILLER_42_21 VDD VSS sg13g2_decap_8
XFILLER_42_98 VDD VSS sg13g2_decap_8
XFILLER_5_357 VDD VSS sg13g2_decap_8
XFILLER_1_574 VDD VSS sg13g2_decap_8
X_80_ _80__4/L_HI VSS VDD _80_/D _80_/Q _83_/CLK sg13g2_dfrbpq_1
XFILLER_76_320 VDD VSS sg13g2_decap_8
XFILLER_67_84 VDD VSS sg13g2_decap_8
XFILLER_49_567 VDD VSS sg13g2_decap_8
XFILLER_37_707 VDD VSS sg13g2_decap_8
XFILLER_64_504 VDD VSS sg13g2_decap_8
XFILLER_91_301 VDD VSS sg13g2_decap_8
XFILLER_36_217 VDD VSS sg13g2_decap_8
XFILLER_76_397 VDD VSS sg13g2_fill_2
XFILLER_17_420 VDD VSS sg13g2_decap_8
XFILLER_29_280 VDD VSS sg13g2_decap_8
XFILLER_91_378 VDD VSS sg13g2_decap_8
XFILLER_60_721 VDD VSS sg13g2_decap_8
XFILLER_17_497 VDD VSS sg13g2_decap_8
XFILLER_32_434 VDD VSS sg13g2_decap_8
XFILLER_44_294 VDD VSS sg13g2_decap_8
XFILLER_9_630 VDD VSS sg13g2_decap_8
XFILLER_8_140 VDD VSS sg13g2_decap_8
XFILLER_95_651 VDD VSS sg13g2_decap_8
XFILLER_67_331 VDD VSS sg13g2_decap_8
XFILLER_28_707 VDD VSS sg13g2_decap_8
XFILLER_94_161 VDD VSS sg13g2_decap_8
XFILLER_82_301 VDD VSS sg13g2_decap_8
XFILLER_55_504 VDD VSS sg13g2_decap_8
XFILLER_27_217 VDD VSS sg13g2_decap_8
XFILLER_82_378 VDD VSS sg13g2_decap_8
XFILLER_63_592 VDD VSS sg13g2_decap_8
XFILLER_51_721 VDD VSS sg13g2_decap_8
XFILLER_23_434 VDD VSS sg13g2_decap_8
XFILLER_35_294 VDD VSS sg13g2_decap_8
XFILLER_50_231 VDD VSS sg13g2_decap_8
XFILLER_12_35 VDD VSS sg13g2_decap_8
XFILLER_88_28 VDD VSS sg13g2_decap_8
XFILLER_5_7 VDD VSS sg13g2_decap_8
XFILLER_86_651 VDD VSS sg13g2_decap_8
XFILLER_85_161 VDD VSS sg13g2_decap_8
XFILLER_46_504 VDD VSS sg13g2_decap_8
XFILLER_37_21 VDD VSS sg13g2_decap_8
XFILLER_58_364 VDD VSS sg13g2_decap_8
XFILLER_19_707 VDD VSS sg13g2_decap_8
XFILLER_18_217 VDD VSS sg13g2_decap_8
XFILLER_61_518 VDD VSS sg13g2_decap_8
XFILLER_37_98 VDD VSS sg13g2_decap_8
XFILLER_54_581 VDD VSS sg13g2_decap_8
XFILLER_42_721 VDD VSS sg13g2_decap_8
XFILLER_53_42 VDD VSS sg13g2_decap_8
XFILLER_14_434 VDD VSS sg13g2_decap_8
XFILLER_41_231 VDD VSS sg13g2_decap_8
XFILLER_10_651 VDD VSS sg13g2_decap_8
XFILLER_6_644 VDD VSS sg13g2_decap_8
XFILLER_5_154 VDD VSS sg13g2_decap_8
XFILLER_69_629 VDD VSS sg13g2_decap_8
XFILLER_1_371 VDD VSS sg13g2_decap_8
XFILLER_38_7 VDD VSS sg13g2_decap_8
XFILLER_76_161 VDD VSS sg13g2_decap_8
X_63_ _75_/A VDD _64_/A VSS _66_/B _68_/D sg13g2_o21ai_1
XFILLER_64_301 VDD VSS sg13g2_decap_8
XFILLER_49_364 VDD VSS sg13g2_decap_8
XFILLER_37_504 VDD VSS sg13g2_decap_8
XFILLER_77_695 VDD VSS sg13g2_decap_8
XFILLER_92_665 VDD VSS sg13g2_decap_8
XFILLER_52_518 VDD VSS sg13g2_decap_8
XFILLER_91_175 VDD VSS sg13g2_decap_8
XFILLER_64_378 VDD VSS sg13g2_decap_8
XFILLER_33_721 VDD VSS sg13g2_decap_8
XFILLER_45_581 VDD VSS sg13g2_decap_8
XFILLER_17_294 VDD VSS sg13g2_decap_8
XFILLER_32_231 VDD VSS sg13g2_decap_8
XFILLER_60_595 VDD VSS sg13g2_decap_8
XFILLER_20_448 VDD VSS sg13g2_decap_8
XFILLER_64_0 VDD VSS sg13g2_decap_8
XFILLER_87_448 VDD VSS sg13g2_decap_8
XFILLER_4_91 VDD VSS sg13g2_decap_8
XFILLER_55_301 VDD VSS sg13g2_decap_8
XFILLER_28_504 VDD VSS sg13g2_decap_8
XFILLER_67_161 VDD VSS sg13g2_decap_8
XFILLER_83_665 VDD VSS sg13g2_decap_8
XFILLER_82_175 VDD VSS sg13g2_decap_8
XFILLER_55_378 VDD VSS sg13g2_decap_8
XFILLER_24_721 VDD VSS sg13g2_decap_8
XFILLER_36_581 VDD VSS sg13g2_decap_8
XFILLER_43_518 VDD VSS sg13g2_decap_8
XFILLER_70_348 VDD VSS sg13g2_decap_8
XFILLER_23_231 VDD VSS sg13g2_decap_8
XFILLER_51_595 VDD VSS sg13g2_decap_8
XFILLER_11_448 VDD VSS sg13g2_decap_8
XFILLER_23_56 VDD VSS sg13g2_decap_8
XFILLER_3_658 VDD VSS sg13g2_decap_8
XFILLER_2_168 VDD VSS sg13g2_decap_8
XFILLER_78_448 VDD VSS sg13g2_decap_8
XFILLER_48_42 VDD VSS sg13g2_decap_8
XFILLER_59_651 VDD VSS sg13g2_decap_8
XFILLER_19_504 VDD VSS sg13g2_decap_8
XFILLER_46_301 VDD VSS sg13g2_decap_8
XFILLER_58_161 VDD VSS sg13g2_decap_8
XFILLER_74_665 VDD VSS sg13g2_decap_8
XFILLER_0_49 VDD VSS sg13g2_decap_8
XFILLER_73_175 VDD VSS sg13g2_decap_8
XFILLER_64_63 VDD VSS sg13g2_decap_8
XFILLER_46_378 VDD VSS sg13g2_decap_8
XFILLER_61_315 VDD VSS sg13g2_decap_8
XFILLER_15_721 VDD VSS sg13g2_decap_8
XFILLER_27_581 VDD VSS sg13g2_decap_8
XFILLER_34_518 VDD VSS sg13g2_decap_8
XFILLER_14_231 VDD VSS sg13g2_decap_8
XFILLER_9_14 VDD VSS sg13g2_decap_8
XFILLER_30_735 VDD VSS sg13g2_decap_8
XFILLER_42_595 VDD VSS sg13g2_decap_8
XFILLER_80_84 VDD VSS sg13g2_decap_8
XFILLER_6_441 VDD VSS sg13g2_decap_8
XFILLER_69_415 VDD VSS sg13g2_decap_8
XFILLER_77_492 VDD VSS sg13g2_decap_8
XFILLER_37_301 VDD VSS sg13g2_decap_8
XFILLER_49_161 VDD VSS sg13g2_decap_8
XFILLER_65_654 VDD VSS sg13g2_decap_8
X_46_ VDD _60_/A _78_/Q VSS sg13g2_inv_1
XFILLER_80_602 VDD VSS sg13g2_decap_8
XFILLER_92_462 VDD VSS sg13g2_decap_8
XFILLER_64_175 VDD VSS sg13g2_decap_8
XFILLER_37_378 VDD VSS sg13g2_decap_8
XFILLER_52_315 VDD VSS sg13g2_decap_8
XFILLER_25_518 VDD VSS sg13g2_decap_8
XFILLER_18_581 VDD VSS sg13g2_decap_8
XFILLER_80_679 VDD VSS sg13g2_decap_8
XFILLER_60_392 VDD VSS sg13g2_decap_8
XFILLER_21_735 VDD VSS sg13g2_decap_8
XFILLER_33_595 VDD VSS sg13g2_decap_8
XFILLER_20_245 VDD VSS sg13g2_decap_8
XFILLER_88_735 VDD VSS sg13g2_decap_8
XFILLER_87_245 VDD VSS sg13g2_decap_8
XFILLER_28_301 VDD VSS sg13g2_decap_8
XFILLER_56_665 VDD VSS sg13g2_decap_8
XFILLER_18_56 VDD VSS sg13g2_decap_8
XFILLER_83_462 VDD VSS sg13g2_decap_8
XFILLER_28_378 VDD VSS sg13g2_decap_8
XFILLER_43_315 VDD VSS sg13g2_decap_8
XFILLER_55_175 VDD VSS sg13g2_decap_8
XFILLER_16_518 VDD VSS sg13g2_decap_8
XFILLER_71_646 VDD VSS sg13g2_decap_8
XFILLER_70_112 VDD VSS sg13g2_decap_8
XFILLER_12_735 VDD VSS sg13g2_decap_8
XFILLER_34_77 VDD VSS sg13g2_decap_8
XFILLER_51_392 VDD VSS sg13g2_decap_8
XFILLER_24_595 VDD VSS sg13g2_decap_8
XFILLER_8_728 VDD VSS sg13g2_decap_8
XFILLER_11_245 VDD VSS sg13g2_decap_8
XFILLER_7_238 VDD VSS sg13g2_decap_8
XFILLER_50_21 VDD VSS sg13g2_decap_8
XFILLER_50_98 VDD VSS sg13g2_decap_8
XFILLER_79_735 VDD VSS sg13g2_decap_8
XFILLER_3_455 VDD VSS sg13g2_decap_8
XFILLER_78_245 VDD VSS sg13g2_decap_8
XFILLER_59_63 VDD VSS sg13g2_decap_8
XFILLER_94_749 VDD VSS sg13g2_decap_8
XFILLER_19_301 VDD VSS sg13g2_decap_8
XFILLER_93_259 VDD VSS sg13g2_decap_8
XFILLER_47_665 VDD VSS sg13g2_decap_8
XFILLER_62_602 VDD VSS sg13g2_decap_8
XFILLER_74_462 VDD VSS sg13g2_decap_8
XFILLER_75_95 VDD VSS sg13g2_decap_8
XFILLER_19_378 VDD VSS sg13g2_decap_8
XFILLER_34_315 VDD VSS sg13g2_decap_8
XFILLER_46_175 VDD VSS sg13g2_decap_8
XFILLER_61_112 VDD VSS sg13g2_decap_8
XFILLER_62_679 VDD VSS sg13g2_decap_8
XFILLER_61_189 VDD VSS sg13g2_decap_8
XFILLER_15_595 VDD VSS sg13g2_decap_8
XFILLER_42_392 VDD VSS sg13g2_decap_8
XFILLER_30_532 VDD VSS sg13g2_decap_8
XFILLER_27_0 VDD VSS sg13g2_decap_8
XFILLER_85_749 VDD VSS sg13g2_decap_8
XFILLER_69_289 VDD VSS sg13g2_decap_8
XFILLER_84_259 VDD VSS sg13g2_decap_8
XFILLER_38_665 VDD VSS sg13g2_decap_8
XFILLER_65_462 VDD VSS sg13g2_decap_8
XFILLER_53_602 VDD VSS sg13g2_decap_8
XFILLER_1_70 VDD VSS sg13g2_decap_8
XIO_BOND_inputs\[6\].input_pad input_PAD[6] bondpad_70x70_novias
XFILLER_25_315 VDD VSS sg13g2_decap_8
XFILLER_37_175 VDD VSS sg13g2_decap_8
XFILLER_52_112 VDD VSS sg13g2_decap_8
XFILLER_80_476 VDD VSS sg13g2_decap_8
XFILLER_53_679 VDD VSS sg13g2_decap_8
XFILLER_40_329 VDD VSS sg13g2_decap_8
XFILLER_52_189 VDD VSS sg13g2_decap_8
XFILLER_33_392 VDD VSS sg13g2_decap_8
XFILLER_21_532 VDD VSS sg13g2_decap_8
XFILLER_20_35 VDD VSS sg13g2_decap_8
XFILLER_88_532 VDD VSS sg13g2_decap_8
XFILLER_76_727 VDD VSS sg13g2_decap_8
Xhold22 _83_/Q VDD VSS _43_/A sg13g2_dlygate4sd3_1
XFILLER_0_469 VDD VSS sg13g2_decap_8
Xhold11 hold11/A VDD VSS _75_/A sg13g2_dlygate4sd3_1
XFILLER_75_237 VDD VSS sg13g2_fill_1
XFILLER_29_77 VDD VSS sg13g2_decap_8
XFILLER_29_665 VDD VSS sg13g2_decap_8
XFILLER_45_21 VDD VSS sg13g2_decap_8
XFILLER_16_315 VDD VSS sg13g2_decap_8
XFILLER_28_175 VDD VSS sg13g2_decap_8
XFILLER_56_462 VDD VSS sg13g2_decap_8
XFILLER_44_602 VDD VSS sg13g2_decap_8
XFILLER_71_443 VDD VSS sg13g2_decap_8
XFILLER_43_112 VDD VSS sg13g2_decap_8
XFILLER_45_98 VDD VSS sg13g2_decap_8
XFILLER_44_679 VDD VSS sg13g2_decap_8
XFILLER_31_329 VDD VSS sg13g2_decap_8
XFILLER_43_189 VDD VSS sg13g2_decap_8
XFILLER_12_532 VDD VSS sg13g2_decap_8
XFILLER_61_42 VDD VSS sg13g2_decap_8
XFILLER_24_392 VDD VSS sg13g2_decap_8
XFILLER_8_525 VDD VSS sg13g2_decap_8
XFILLER_4_742 VDD VSS sg13g2_decap_8
XFILLER_3_252 VDD VSS sg13g2_decap_8
XFILLER_79_532 VDD VSS sg13g2_decap_8
XFILLER_67_716 VDD VSS sg13g2_decap_8
XFILLER_20_7 VDD VSS sg13g2_decap_8
XFILLER_94_546 VDD VSS sg13g2_decap_8
XFILLER_66_259 VDD VSS sg13g2_decap_8
XFILLER_47_462 VDD VSS sg13g2_decap_8
XFILLER_35_602 VDD VSS sg13g2_decap_8
XFILLER_19_175 VDD VSS sg13g2_decap_8
XFILLER_34_112 VDD VSS sg13g2_decap_8
XFILLER_62_476 VDD VSS sg13g2_decap_8
XFILLER_50_616 VDD VSS sg13g2_decap_8
XFILLER_35_679 VDD VSS sg13g2_decap_8
XFILLER_22_329 VDD VSS sg13g2_decap_8
XFILLER_34_189 VDD VSS sg13g2_decap_8
XFILLER_15_392 VDD VSS sg13g2_decap_8
XFILLER_89_329 VDD VSS sg13g2_decap_8
XFILLER_58_749 VDD VSS sg13g2_decap_8
XFILLER_85_546 VDD VSS sg13g2_decap_8
XFILLER_57_259 VDD VSS sg13g2_decap_8
XFILLER_38_462 VDD VSS sg13g2_decap_8
XFILLER_25_112 VDD VSS sg13g2_decap_8
XFILLER_26_657 VDD VSS sg13g2_decap_8
XFILLER_53_476 VDD VSS sg13g2_decap_8
XFILLER_41_616 VDD VSS sg13g2_decap_8
XFILLER_80_273 VDD VSS sg13g2_decap_8
XFILLER_13_329 VDD VSS sg13g2_decap_8
XFILLER_15_35 VDD VSS sg13g2_decap_8
XFILLER_25_189 VDD VSS sg13g2_decap_8
XFILLER_40_126 VDD VSS sg13g2_decap_8
XFILLER_31_56 VDD VSS sg13g2_decap_8
XFILLER_5_539 VDD VSS sg13g2_decap_8
XFILLER_1_756 VDD VSS sg13g2_fill_1
XFILLER_76_524 VDD VSS sg13g2_decap_8
XFILLER_49_749 VDD VSS sg13g2_decap_8
XFILLER_0_266 VDD VSS sg13g2_decap_8
XFILLER_48_259 VDD VSS sg13g2_decap_8
XFILLER_56_42 VDD VSS sg13g2_decap_8
XFILLER_29_462 VDD VSS sg13g2_decap_8
XFILLER_17_602 VDD VSS sg13g2_decap_8
XFILLER_16_112 VDD VSS sg13g2_decap_8
XFILLER_17_679 VDD VSS sg13g2_decap_8
XFILLER_71_284 VDD VSS sg13g2_fill_1
XFILLER_16_189 VDD VSS sg13g2_decap_8
XFILLER_44_476 VDD VSS sg13g2_decap_8
XFILLER_32_616 VDD VSS sg13g2_decap_8
XFILLER_72_63 VDD VSS sg13g2_decap_8
XFILLER_31_126 VDD VSS sg13g2_decap_8
XFILLER_8_322 VDD VSS sg13g2_decap_8
XFILLER_40_693 VDD VSS sg13g2_decap_8
XFILLER_68_7 VDD VSS sg13g2_decap_8
XFILLER_8_399 VDD VSS sg13g2_decap_8
XFILLER_67_513 VDD VSS sg13g2_decap_8
XFILLER_94_343 VDD VSS sg13g2_decap_8
XFILLER_39_259 VDD VSS sg13g2_decap_8
XFILLER_90_560 VDD VSS sg13g2_decap_8
XFILLER_62_273 VDD VSS sg13g2_decap_8
XFILLER_35_476 VDD VSS sg13g2_decap_8
XFILLER_50_413 VDD VSS sg13g2_decap_8
XFILLER_23_616 VDD VSS sg13g2_decap_8
XFILLER_94_0 VDD VSS sg13g2_decap_8
XFILLER_22_126 VDD VSS sg13g2_decap_8
XFILLER_31_693 VDD VSS sg13g2_decap_8
XFILLER_7_91 VDD VSS sg13g2_decap_8
XFILLER_89_126 VDD VSS sg13g2_decap_8
XFILLER_85_343 VDD VSS sg13g2_decap_8
XFILLER_58_546 VDD VSS sg13g2_decap_8
XFILLER_73_527 VDD VSS sg13g2_decap_8
XFILLER_66_590 VDD VSS sg13g2_decap_8
XFILLER_26_56 VDD VSS sg13g2_decap_8
XFILLER_26_454 VDD VSS sg13g2_decap_8
XFILLER_81_560 VDD VSS sg13g2_decap_8
XFILLER_41_413 VDD VSS sg13g2_decap_8
XFILLER_53_273 VDD VSS sg13g2_decap_8
XFILLER_14_616 VDD VSS sg13g2_decap_8
XFILLER_13_126 VDD VSS sg13g2_decap_8
XFILLER_9_119 VDD VSS sg13g2_decap_8
XFILLER_42_77 VDD VSS sg13g2_decap_8
XFILLER_22_693 VDD VSS sg13g2_decap_8
XFILLER_5_336 VDD VSS sg13g2_decap_8
XFILLER_1_553 VDD VSS sg13g2_decap_8
XFILLER_89_693 VDD VSS sg13g2_decap_8
XFILLER_3_49 VDD VSS sg13g2_decap_8
XFILLER_67_63 VDD VSS sg13g2_decap_8
XFILLER_49_546 VDD VSS sg13g2_decap_8
XFILLER_76_376 VDD VSS sg13g2_decap_8
XFILLER_91_357 VDD VSS sg13g2_decap_8
XFILLER_83_84 VDD VSS sg13g2_decap_8
XFILLER_60_700 VDD VSS sg13g2_decap_8
XFILLER_17_476 VDD VSS sg13g2_decap_8
XFILLER_32_413 VDD VSS sg13g2_decap_8
XFILLER_44_273 VDD VSS sg13g2_decap_8
XFILLER_72_593 VDD VSS sg13g2_decap_8
XFILLER_13_693 VDD VSS sg13g2_decap_8
XFILLER_40_490 VDD VSS sg13g2_decap_8
XFILLER_9_686 VDD VSS sg13g2_decap_8
XFILLER_8_196 VDD VSS sg13g2_decap_8
XFILLER_95_630 VDD VSS sg13g2_decap_8
XFILLER_67_310 VDD VSS sg13g2_decap_8
XFILLER_94_140 VDD VSS sg13g2_decap_8
XFILLER_67_387 VDD VSS sg13g2_decap_8
XFILLER_70_519 VDD VSS sg13g2_decap_8
XFILLER_82_357 VDD VSS sg13g2_decap_8
XFILLER_63_571 VDD VSS sg13g2_decap_8
XFILLER_51_700 VDD VSS sg13g2_decap_8
XFILLER_23_413 VDD VSS sg13g2_decap_8
XFILLER_35_273 VDD VSS sg13g2_decap_8
XFILLER_50_210 VDD VSS sg13g2_decap_8
XFILLER_50_287 VDD VSS sg13g2_decap_8
XFILLER_12_14 VDD VSS sg13g2_decap_8
XFILLER_31_490 VDD VSS sg13g2_decap_8
XFILLER_86_630 VDD VSS sg13g2_decap_8
XFILLER_85_140 VDD VSS sg13g2_decap_8
XFILLER_58_343 VDD VSS sg13g2_decap_8
XFILLER_37_77 VDD VSS sg13g2_decap_8
XFILLER_54_560 VDD VSS sg13g2_decap_8
XFILLER_14_413 VDD VSS sg13g2_decap_8
XFILLER_26_273 VDD VSS sg13g2_decap_8
XFILLER_42_700 VDD VSS sg13g2_decap_8
XFILLER_53_21 VDD VSS sg13g2_decap_8
XFILLER_41_210 VDD VSS sg13g2_decap_8
XFILLER_53_98 VDD VSS sg13g2_decap_8
XFILLER_41_287 VDD VSS sg13g2_decap_8
XFILLER_10_630 VDD VSS sg13g2_decap_8
XFILLER_22_490 VDD VSS sg13g2_decap_8
XFILLER_6_623 VDD VSS sg13g2_decap_8
XFILLER_5_133 VDD VSS sg13g2_decap_8
XFILLER_69_608 VDD VSS sg13g2_decap_8
XFILLER_78_84 VDD VSS sg13g2_decap_8
XFILLER_1_350 VDD VSS sg13g2_decap_8
XFILLER_89_490 VDD VSS sg13g2_decap_8
XFILLER_77_674 VDD VSS sg13g2_decap_8
XFILLER_76_140 VDD VSS sg13g2_decap_8
X_62_ _78_/Q _66_/D _66_/B _65_/B VDD VSS sg13g2_nand3_1
XFILLER_49_343 VDD VSS sg13g2_decap_8
XFILLER_92_644 VDD VSS sg13g2_decap_8
XFILLER_91_154 VDD VSS sg13g2_decap_8
XFILLER_64_357 VDD VSS sg13g2_decap_8
XFILLER_17_273 VDD VSS sg13g2_decap_8
XFILLER_33_700 VDD VSS sg13g2_decap_8
XFILLER_45_560 VDD VSS sg13g2_decap_8
XFILLER_32_210 VDD VSS sg13g2_decap_8
XFILLER_60_574 VDD VSS sg13g2_decap_8
XFILLER_20_427 VDD VSS sg13g2_decap_8
XFILLER_32_287 VDD VSS sg13g2_decap_8
XFILLER_13_490 VDD VSS sg13g2_decap_8
XFILLER_9_483 VDD VSS sg13g2_decap_8
XFILLER_57_0 VDD VSS sg13g2_decap_8
XFILLER_87_427 VDD VSS sg13g2_decap_8
XFILLER_4_70 VDD VSS sg13g2_decap_8
XFILLER_67_140 VDD VSS sg13g2_decap_8
XFILLER_68_685 VDD VSS sg13g2_decap_8
XFILLER_83_644 VDD VSS sg13g2_decap_8
XFILLER_55_357 VDD VSS sg13g2_decap_8
XFILLER_82_154 VDD VSS sg13g2_decap_8
XFILLER_70_327 VDD VSS sg13g2_decap_8
XFILLER_24_700 VDD VSS sg13g2_decap_8
XFILLER_36_560 VDD VSS sg13g2_decap_8
XFILLER_23_210 VDD VSS sg13g2_decap_8
XFILLER_51_574 VDD VSS sg13g2_decap_8
XFILLER_11_427 VDD VSS sg13g2_decap_8
XFILLER_23_35 VDD VSS sg13g2_decap_8
XFILLER_23_287 VDD VSS sg13g2_decap_8
XFILLER_3_637 VDD VSS sg13g2_decap_8
XFILLER_2_147 VDD VSS sg13g2_decap_8
XFILLER_78_427 VDD VSS sg13g2_decap_8
XFILLER_59_630 VDD VSS sg13g2_decap_8
XFILLER_48_21 VDD VSS sg13g2_decap_8
XFILLER_58_140 VDD VSS sg13g2_decap_8
XFILLER_48_98 VDD VSS sg13g2_decap_8
XFILLER_74_644 VDD VSS sg13g2_decap_8
XFILLER_0_28 VDD VSS sg13g2_decap_8
XFILLER_46_357 VDD VSS sg13g2_decap_8
XFILLER_73_154 VDD VSS sg13g2_decap_8
XFILLER_64_42 VDD VSS sg13g2_decap_8
XFILLER_15_700 VDD VSS sg13g2_decap_8
XFILLER_27_560 VDD VSS sg13g2_decap_8
XFILLER_14_210 VDD VSS sg13g2_decap_8
XFILLER_30_714 VDD VSS sg13g2_decap_8
XFILLER_42_574 VDD VSS sg13g2_decap_8
XFILLER_14_287 VDD VSS sg13g2_decap_8
XFILLER_80_63 VDD VSS sg13g2_decap_8
XFILLER_6_420 VDD VSS sg13g2_decap_8
XFILLER_50_7 VDD VSS sg13g2_decap_8
XFILLER_6_497 VDD VSS sg13g2_decap_8
XFILLER_49_140 VDD VSS sg13g2_decap_8
XFILLER_65_633 VDD VSS sg13g2_decap_8
XFILLER_77_471 VDD VSS sg13g2_decap_8
XIO_BOND_inputs\[5\].input_pad input_PAD[5] bondpad_70x70_novias
XFILLER_92_441 VDD VSS sg13g2_decap_8
X_45_ VDD _74_/C _45_/A VSS sg13g2_inv_1
XFILLER_37_357 VDD VSS sg13g2_decap_8
XFILLER_64_154 VDD VSS sg13g2_decap_8
XFILLER_18_560 VDD VSS sg13g2_decap_8
XFILLER_80_658 VDD VSS sg13g2_decap_8
XFILLER_21_714 VDD VSS sg13g2_decap_8
XFILLER_20_224 VDD VSS sg13g2_decap_8
XFILLER_60_371 VDD VSS sg13g2_decap_8
XFILLER_33_574 VDD VSS sg13g2_decap_8
XFILLER_9_280 VDD VSS sg13g2_decap_8
XFILLER_88_714 VDD VSS sg13g2_decap_8
XFILLER_87_224 VDD VSS sg13g2_decap_8
XFILLER_68_482 VDD VSS sg13g2_decap_8
XFILLER_18_35 VDD VSS sg13g2_decap_8
XFILLER_83_441 VDD VSS sg13g2_decap_8
XFILLER_56_644 VDD VSS sg13g2_decap_8
XFILLER_28_357 VDD VSS sg13g2_decap_8
XFILLER_71_625 VDD VSS sg13g2_decap_8
XFILLER_55_154 VDD VSS sg13g2_decap_8
XFILLER_70_168 VDD VSS sg13g2_decap_8
XFILLER_12_714 VDD VSS sg13g2_decap_8
XFILLER_34_56 VDD VSS sg13g2_decap_8
XFILLER_51_371 VDD VSS sg13g2_decap_8
XFILLER_24_574 VDD VSS sg13g2_decap_8
XFILLER_8_707 VDD VSS sg13g2_decap_8
XFILLER_11_224 VDD VSS sg13g2_decap_8
XFILLER_7_217 VDD VSS sg13g2_decap_8
XFILLER_50_77 VDD VSS sg13g2_decap_8
XFILLER_3_434 VDD VSS sg13g2_decap_8
XFILLER_79_714 VDD VSS sg13g2_decap_8
XFILLER_59_42 VDD VSS sg13g2_decap_8
XFILLER_78_224 VDD VSS sg13g2_decap_8
XFILLER_94_728 VDD VSS sg13g2_decap_8
XFILLER_93_238 VDD VSS sg13g2_decap_8
XFILLER_74_430 VDD VSS sg13g2_decap_8
XFILLER_47_644 VDD VSS sg13g2_decap_8
XFILLER_19_357 VDD VSS sg13g2_decap_8
XFILLER_75_74 VDD VSS sg13g2_decap_8
XFILLER_46_154 VDD VSS sg13g2_decap_8
XFILLER_62_658 VDD VSS sg13g2_decap_8
XFILLER_61_168 VDD VSS sg13g2_decap_8
XFILLER_70_680 VDD VSS sg13g2_decap_8
XFILLER_91_84 VDD VSS sg13g2_decap_8
XFILLER_42_371 VDD VSS sg13g2_decap_8
XFILLER_15_574 VDD VSS sg13g2_decap_8
XFILLER_30_511 VDD VSS sg13g2_decap_8
XFILLER_30_588 VDD VSS sg13g2_decap_8
XFILLER_6_294 VDD VSS sg13g2_decap_8
XFILLER_69_224 VDD VSS sg13g2_decap_8
XFILLER_69_268 VDD VSS sg13g2_decap_8
XFILLER_85_728 VDD VSS sg13g2_decap_8
XFILLER_84_238 VDD VSS sg13g2_decap_8
XFILLER_65_441 VDD VSS sg13g2_decap_8
XFILLER_38_644 VDD VSS sg13g2_decap_8
XFILLER_37_154 VDD VSS sg13g2_decap_8
XFILLER_53_658 VDD VSS sg13g2_decap_8
XFILLER_80_455 VDD VSS sg13g2_decap_8
XFILLER_40_308 VDD VSS sg13g2_decap_8
XFILLER_52_168 VDD VSS sg13g2_decap_8
XFILLER_33_371 VDD VSS sg13g2_decap_8
XFILLER_21_511 VDD VSS sg13g2_decap_8
XFILLER_21_588 VDD VSS sg13g2_decap_8
XFILLER_20_14 VDD VSS sg13g2_decap_8
XFILLER_88_511 VDD VSS sg13g2_decap_8
XFILLER_76_706 VDD VSS sg13g2_decap_8
Xhold23 _80_/Q VDD VSS hold23/X sg13g2_dlygate4sd3_1
Xhold12 _71_/Y VDD VSS _72_/B1 sg13g2_dlygate4sd3_1
XFILLER_0_448 VDD VSS sg13g2_decap_8
XFILLER_88_588 VDD VSS sg13g2_decap_8
XFILLER_29_56 VDD VSS sg13g2_decap_8
XFILLER_56_441 VDD VSS sg13g2_decap_8
XFILLER_29_644 VDD VSS sg13g2_decap_8
XFILLER_28_154 VDD VSS sg13g2_decap_8
XFILLER_71_422 VDD VSS sg13g2_decap_8
XFILLER_44_658 VDD VSS sg13g2_decap_8
XFILLER_45_77 VDD VSS sg13g2_decap_8
XFILLER_31_308 VDD VSS sg13g2_decap_8
XFILLER_43_168 VDD VSS sg13g2_decap_8
XFILLER_71_499 VDD VSS sg13g2_decap_8
XFILLER_12_511 VDD VSS sg13g2_decap_8
XFILLER_24_371 VDD VSS sg13g2_decap_8
XFILLER_8_504 VDD VSS sg13g2_decap_8
XFILLER_61_21 VDD VSS sg13g2_decap_8
XFILLER_12_588 VDD VSS sg13g2_decap_8
XFILLER_61_98 VDD VSS sg13g2_decap_8
XFILLER_6_49 VDD VSS sg13g2_decap_8
XFILLER_4_721 VDD VSS sg13g2_decap_8
XFILLER_3_231 VDD VSS sg13g2_decap_8
XFILLER_79_511 VDD VSS sg13g2_decap_8
XFILLER_10_91 VDD VSS sg13g2_decap_8
XFILLER_94_525 VDD VSS sg13g2_decap_8
XFILLER_79_588 VDD VSS sg13g2_decap_8
XFILLER_66_238 VDD VSS sg13g2_decap_8
XFILLER_86_84 VDD VSS sg13g2_decap_8
XFILLER_13_7 VDD VSS sg13g2_decap_8
XFILLER_47_441 VDD VSS sg13g2_decap_8
XFILLER_19_154 VDD VSS sg13g2_decap_8
XFILLER_90_742 VDD VSS sg13g2_decap_8
XFILLER_74_293 VDD VSS sg13g2_decap_4
XFILLER_62_455 VDD VSS sg13g2_fill_2
XFILLER_35_658 VDD VSS sg13g2_decap_8
XFILLER_15_371 VDD VSS sg13g2_decap_8
XFILLER_22_308 VDD VSS sg13g2_decap_8
XFILLER_34_168 VDD VSS sg13g2_decap_8
XFILLER_30_385 VDD VSS sg13g2_decap_8
XFILLER_7_581 VDD VSS sg13g2_decap_8
XFILLER_89_308 VDD VSS sg13g2_decap_8
XFILLER_85_525 VDD VSS sg13g2_decap_8
XFILLER_58_728 VDD VSS sg13g2_decap_8
XFILLER_73_709 VDD VSS sg13g2_decap_8
XFILLER_57_238 VDD VSS sg13g2_decap_8
XFILLER_38_441 VDD VSS sg13g2_decap_8
XFILLER_81_742 VDD VSS sg13g2_decap_8
XFILLER_26_636 VDD VSS sg13g2_decap_8
XFILLER_80_252 VDD VSS sg13g2_decap_8
XFILLER_15_14 VDD VSS sg13g2_decap_8
XFILLER_53_455 VDD VSS sg13g2_decap_8
XFILLER_13_308 VDD VSS sg13g2_decap_8
XFILLER_40_105 VDD VSS sg13g2_decap_8
XFILLER_25_168 VDD VSS sg13g2_decap_8
XFILLER_31_35 VDD VSS sg13g2_decap_8
XFILLER_21_385 VDD VSS sg13g2_decap_8
XFILLER_5_518 VDD VSS sg13g2_decap_8
XFILLER_1_735 VDD VSS sg13g2_decap_8
XFILLER_0_245 VDD VSS sg13g2_decap_8
XFILLER_76_503 VDD VSS sg13g2_decap_8
XFILLER_88_385 VDD VSS sg13g2_decap_8
XFILLER_49_728 VDD VSS sg13g2_decap_8
XFILLER_56_21 VDD VSS sg13g2_decap_8
XFILLER_48_238 VDD VSS sg13g2_decap_8
XFILLER_29_441 VDD VSS sg13g2_decap_8
XFILLER_91_539 VDD VSS sg13g2_decap_8
XFILLER_56_98 VDD VSS sg13g2_decap_8
XFILLER_44_455 VDD VSS sg13g2_decap_8
XFILLER_17_658 VDD VSS sg13g2_decap_8
XFILLER_71_263 VDD VSS sg13g2_decap_8
XFILLER_72_42 VDD VSS sg13g2_decap_8
XFILLER_31_105 VDD VSS sg13g2_decap_8
XFILLER_16_168 VDD VSS sg13g2_decap_8
XFILLER_8_301 VDD VSS sg13g2_decap_8
XFILLER_40_672 VDD VSS sg13g2_decap_8
XFILLER_12_385 VDD VSS sg13g2_decap_8
XFILLER_8_378 VDD VSS sg13g2_decap_8
XFILLER_4_595 VDD VSS sg13g2_decap_8
XFILLER_79_385 VDD VSS sg13g2_decap_8
XFILLER_94_322 VDD VSS sg13g2_decap_8
XFILLER_39_238 VDD VSS sg13g2_decap_8
XFILLER_67_569 VDD VSS sg13g2_decap_8
XFILLER_82_539 VDD VSS sg13g2_decap_8
XFILLER_94_399 VDD VSS sg13g2_decap_8
XFILLER_63_753 VDD VSS sg13g2_decap_4
XFILLER_35_455 VDD VSS sg13g2_decap_8
XFILLER_62_252 VDD VSS sg13g2_decap_8
XFILLER_22_105 VDD VSS sg13g2_decap_8
XFILLER_87_0 VDD VSS sg13g2_decap_8
XFILLER_50_469 VDD VSS sg13g2_decap_8
XFILLER_31_672 VDD VSS sg13g2_decap_8
XFILLER_30_182 VDD VSS sg13g2_decap_8
XFILLER_7_70 VDD VSS sg13g2_decap_8
XFILLER_89_105 VDD VSS sg13g2_decap_8
XFILLER_58_525 VDD VSS sg13g2_decap_8
XFILLER_85_322 VDD VSS sg13g2_decap_8
XFILLER_73_506 VDD VSS sg13g2_decap_8
XFILLER_85_399 VDD VSS sg13g2_decap_8
XFILLER_54_742 VDD VSS sg13g2_decap_8
XFILLER_26_35 VDD VSS sg13g2_decap_8
XFILLER_26_433 VDD VSS sg13g2_decap_8
XFILLER_13_105 VDD VSS sg13g2_decap_8
XFILLER_53_252 VDD VSS sg13g2_decap_8
XFILLER_41_469 VDD VSS sg13g2_decap_8
XFILLER_42_56 VDD VSS sg13g2_decap_8
XFILLER_22_672 VDD VSS sg13g2_decap_8
XFILLER_21_182 VDD VSS sg13g2_decap_8
XFILLER_5_315 VDD VSS sg13g2_decap_8
XFILLER_1_532 VDD VSS sg13g2_decap_8
XFILLER_3_28 VDD VSS sg13g2_decap_8
XFILLER_89_672 VDD VSS sg13g2_decap_8
XFILLER_95_119 VDD VSS sg13g2_decap_8
XFILLER_88_182 VDD VSS sg13g2_decap_8
XFILLER_67_42 VDD VSS sg13g2_decap_8
XFILLER_49_525 VDD VSS sg13g2_decap_8
XFILLER_76_355 VDD VSS sg13g2_decap_8
XFILLER_64_539 VDD VSS sg13g2_decap_8
XFILLER_91_336 VDD VSS sg13g2_decap_8
XFILLER_17_455 VDD VSS sg13g2_decap_8
XFILLER_45_742 VDD VSS sg13g2_decap_8
XFILLER_72_572 VDD VSS sg13g2_decap_8
XFILLER_83_63 VDD VSS sg13g2_decap_8
XFILLER_44_252 VDD VSS sg13g2_decap_8
XFILLER_60_756 VDD VSS sg13g2_fill_1
XFILLER_32_469 VDD VSS sg13g2_decap_8
XFILLER_20_609 VDD VSS sg13g2_decap_8
XFILLER_80_7 VDD VSS sg13g2_decap_8
XFILLER_13_672 VDD VSS sg13g2_decap_8
XFILLER_9_665 VDD VSS sg13g2_decap_8
XFILLER_12_182 VDD VSS sg13g2_decap_8
XFILLER_8_175 VDD VSS sg13g2_decap_8
XFILLER_87_609 VDD VSS sg13g2_decap_8
XFILLER_4_392 VDD VSS sg13g2_decap_8
XFILLER_86_119 VDD VSS sg13g2_decap_8
XFILLER_79_182 VDD VSS sg13g2_decap_8
XFILLER_67_366 VDD VSS sg13g2_decap_8
XFILLER_95_686 VDD VSS sg13g2_decap_8
XFILLER_82_336 VDD VSS sg13g2_decap_8
XFILLER_55_539 VDD VSS sg13g2_decap_8
XFILLER_94_196 VDD VSS sg13g2_decap_8
XFILLER_36_742 VDD VSS sg13g2_decap_8
XFILLER_63_550 VDD VSS sg13g2_decap_8
XFILLER_35_252 VDD VSS sg13g2_decap_8
XFILLER_51_756 VDD VSS sg13g2_fill_1
XFILLER_11_609 VDD VSS sg13g2_decap_8
XFILLER_23_469 VDD VSS sg13g2_decap_8
XFILLER_50_266 VDD VSS sg13g2_decap_8
XFILLER_10_119 VDD VSS sg13g2_decap_8
XFILLER_2_329 VDD VSS sg13g2_decap_8
XFILLER_78_609 VDD VSS sg13g2_decap_8
XFILLER_77_119 VDD VSS sg13g2_decap_8
XFILLER_58_322 VDD VSS sg13g2_decap_8
XFILLER_86_686 VDD VSS sg13g2_decap_8
XFILLER_73_325 VDD VSS sg13g2_decap_8
XFILLER_46_539 VDD VSS sg13g2_decap_8
XFILLER_37_56 VDD VSS sg13g2_decap_8
XFILLER_58_399 VDD VSS sg13g2_decap_8
XFILLER_85_196 VDD VSS sg13g2_decap_8
XFILLER_27_742 VDD VSS sg13g2_decap_8
XFILLER_26_252 VDD VSS sg13g2_decap_8
XFILLER_42_756 VDD VSS sg13g2_fill_1
XFILLER_53_77 VDD VSS sg13g2_decap_8
XFILLER_14_469 VDD VSS sg13g2_decap_8
XFILLER_41_266 VDD VSS sg13g2_decap_8
XFILLER_6_602 VDD VSS sg13g2_decap_8
XFILLER_10_686 VDD VSS sg13g2_decap_8
XFILLER_5_112 VDD VSS sg13g2_decap_8
XFILLER_6_679 VDD VSS sg13g2_decap_8
XFILLER_5_189 VDD VSS sg13g2_decap_8
XFILLER_68_119 VDD VSS sg13g2_decap_8
XFILLER_78_63 VDD VSS sg13g2_decap_8
XFILLER_49_322 VDD VSS sg13g2_decap_8
XFILLER_77_653 VDD VSS sg13g2_decap_8
X_61_ _61_/A _61_/B _68_/D _61_/Y VDD VSS sg13g2_nor3_1
XIO_BOND_inputs\[4\].input_pad input_PAD[4] bondpad_70x70_novias
XFILLER_92_623 VDD VSS sg13g2_decap_8
XFILLER_49_399 VDD VSS sg13g2_decap_8
XFILLER_37_539 VDD VSS sg13g2_decap_8
XFILLER_91_133 VDD VSS sg13g2_decap_8
XFILLER_76_196 VDD VSS sg13g2_decap_8
XFILLER_64_336 VDD VSS sg13g2_decap_8
XFILLER_94_84 VDD VSS sg13g2_decap_8
XFILLER_18_742 VDD VSS sg13g2_decap_8
XFILLER_17_252 VDD VSS sg13g2_decap_8
XFILLER_33_756 VDD VSS sg13g2_fill_1
XFILLER_60_553 VDD VSS sg13g2_decap_8
XFILLER_20_406 VDD VSS sg13g2_decap_8
XFILLER_32_266 VDD VSS sg13g2_decap_8
XFILLER_9_462 VDD VSS sg13g2_decap_8
XFILLER_87_406 VDD VSS sg13g2_decap_8
XFILLER_59_119 VDD VSS sg13g2_decap_8
XFILLER_68_664 VDD VSS sg13g2_decap_8
XFILLER_95_483 VDD VSS sg13g2_decap_8
XFILLER_83_623 VDD VSS sg13g2_decap_8
XFILLER_28_539 VDD VSS sg13g2_decap_8
XFILLER_82_133 VDD VSS sg13g2_decap_8
XFILLER_55_336 VDD VSS sg13g2_decap_8
XFILLER_70_306 VDD VSS sg13g2_decap_8
XFILLER_51_553 VDD VSS sg13g2_decap_8
XFILLER_11_406 VDD VSS sg13g2_decap_8
XFILLER_24_756 VDD VSS sg13g2_fill_1
XFILLER_23_14 VDD VSS sg13g2_decap_8
XFILLER_23_266 VDD VSS sg13g2_decap_8
XFILLER_3_616 VDD VSS sg13g2_decap_8
XFILLER_2_126 VDD VSS sg13g2_decap_8
XFILLER_78_406 VDD VSS sg13g2_decap_8
XFILLER_86_483 VDD VSS sg13g2_decap_8
XFILLER_74_623 VDD VSS sg13g2_decap_8
XFILLER_59_686 VDD VSS sg13g2_decap_8
XFILLER_48_77 VDD VSS sg13g2_decap_8
XFILLER_19_539 VDD VSS sg13g2_decap_8
XFILLER_73_133 VDD VSS sg13g2_decap_8
XFILLER_64_21 VDD VSS sg13g2_decap_8
XFILLER_46_336 VDD VSS sg13g2_decap_8
XFILLER_58_196 VDD VSS sg13g2_decap_8
XFILLER_64_32 VDD VSS sg13g2_fill_1
XFILLER_64_98 VDD VSS sg13g2_decap_8
XFILLER_15_756 VDD VSS sg13g2_fill_1
XFILLER_42_553 VDD VSS sg13g2_decap_8
XFILLER_80_42 VDD VSS sg13g2_decap_8
XFILLER_9_49 VDD VSS sg13g2_decap_8
XFILLER_14_266 VDD VSS sg13g2_decap_8
XFILLER_10_483 VDD VSS sg13g2_decap_8
XFILLER_13_91 VDD VSS sg13g2_decap_8
XFILLER_6_476 VDD VSS sg13g2_decap_8
XFILLER_89_84 VDD VSS sg13g2_decap_8
XFILLER_43_7 VDD VSS sg13g2_decap_8
XFILLER_2_693 VDD VSS sg13g2_decap_8
XFILLER_65_612 VDD VSS sg13g2_decap_8
XFILLER_92_420 VDD VSS sg13g2_decap_8
X_44_ VDD _74_/B _82_/Q VSS sg13g2_inv_1
XFILLER_64_133 VDD VSS sg13g2_decap_8
XFILLER_37_336 VDD VSS sg13g2_decap_8
XFILLER_49_196 VDD VSS sg13g2_decap_8
XFILLER_65_689 VDD VSS sg13g2_decap_8
XFILLER_92_497 VDD VSS sg13g2_decap_8
XFILLER_80_637 VDD VSS sg13g2_decap_8
XFILLER_60_350 VDD VSS sg13g2_decap_8
XFILLER_33_553 VDD VSS sg13g2_decap_8
XFILLER_20_203 VDD VSS sg13g2_decap_8
XFILLER_87_203 VDD VSS sg13g2_decap_8
XFILLER_75_409 VDD VSS sg13g2_decap_8
XFILLER_68_461 VDD VSS sg13g2_decap_8
XFILLER_56_623 VDD VSS sg13g2_decap_8
XFILLER_18_14 VDD VSS sg13g2_decap_8
XFILLER_95_280 VDD VSS sg13g2_decap_8
XFILLER_83_420 VDD VSS sg13g2_decap_8
XFILLER_28_336 VDD VSS sg13g2_decap_8
XFILLER_55_133 VDD VSS sg13g2_decap_8
XFILLER_71_604 VDD VSS sg13g2_decap_8
XFILLER_83_497 VDD VSS sg13g2_decap_8
XFILLER_70_147 VDD VSS sg13g2_decap_8
XFILLER_34_35 VDD VSS sg13g2_decap_8
XFILLER_24_553 VDD VSS sg13g2_decap_8
XFILLER_11_203 VDD VSS sg13g2_decap_8
XFILLER_51_350 VDD VSS sg13g2_decap_8
XFILLER_50_56 VDD VSS sg13g2_decap_8
XFILLER_3_413 VDD VSS sg13g2_decap_8
XFILLER_59_21 VDD VSS sg13g2_decap_8
XFILLER_78_203 VDD VSS sg13g2_decap_8
XFILLER_94_707 VDD VSS sg13g2_decap_8
XFILLER_59_98 VDD VSS sg13g2_decap_8
XFILLER_93_217 VDD VSS sg13g2_decap_8
XFILLER_59_483 VDD VSS sg13g2_decap_8
XFILLER_47_623 VDD VSS sg13g2_decap_8
XFILLER_86_280 VDD VSS sg13g2_decap_8
XFILLER_75_53 VDD VSS sg13g2_decap_8
XFILLER_19_336 VDD VSS sg13g2_decap_8
XFILLER_46_133 VDD VSS sg13g2_decap_8
XFILLER_74_497 VDD VSS sg13g2_decap_8
XFILLER_62_637 VDD VSS sg13g2_decap_8
XFILLER_61_147 VDD VSS sg13g2_decap_8
XFILLER_15_553 VDD VSS sg13g2_decap_8
XFILLER_91_63 VDD VSS sg13g2_decap_8
XFILLER_42_350 VDD VSS sg13g2_decap_8
XFILLER_30_567 VDD VSS sg13g2_decap_8
XFILLER_10_280 VDD VSS sg13g2_decap_8
XFILLER_6_273 VDD VSS sg13g2_decap_8
XFILLER_69_203 VDD VSS sg13g2_decap_8
XFILLER_85_707 VDD VSS sg13g2_decap_8
XFILLER_69_247 VDD VSS sg13g2_decap_8
XFILLER_2_490 VDD VSS sg13g2_decap_8
XFILLER_84_217 VDD VSS sg13g2_decap_8
XFILLER_38_623 VDD VSS sg13g2_decap_8
XFILLER_65_420 VDD VSS sg13g2_decap_8
XFILLER_37_133 VDD VSS sg13g2_decap_8
XFILLER_65_475 VDD VSS sg13g2_fill_2
XFILLER_65_486 VDD VSS sg13g2_decap_8
XFILLER_92_294 VDD VSS sg13g2_decap_8
XFILLER_80_434 VDD VSS sg13g2_decap_8
XFILLER_53_637 VDD VSS sg13g2_decap_8
XFILLER_52_147 VDD VSS sg13g2_decap_8
XFILLER_33_350 VDD VSS sg13g2_decap_8
XFILLER_21_567 VDD VSS sg13g2_decap_8
XFILLER_0_427 VDD VSS sg13g2_decap_8
XFILLER_88_567 VDD VSS sg13g2_decap_8
Xhold13 _72_/Y VDD VSS _82_/D sg13g2_dlygate4sd3_1
XFILLER_29_35 VDD VSS sg13g2_decap_8
Xhold24 _65_/Y VDD VSS _67_/B sg13g2_dlygate4sd3_1
XFILLER_75_228 VDD VSS sg13g2_decap_8
XFILLER_56_420 VDD VSS sg13g2_decap_8
XFILLER_29_623 VDD VSS sg13g2_decap_8
XFILLER_28_133 VDD VSS sg13g2_decap_8
XFILLER_83_294 VDD VSS sg13g2_decap_8
XFILLER_56_497 VDD VSS sg13g2_decap_8
XFILLER_45_56 VDD VSS sg13g2_decap_8
XFILLER_44_637 VDD VSS sg13g2_decap_8
XFILLER_43_147 VDD VSS sg13g2_decap_8
XFILLER_71_478 VDD VSS sg13g2_decap_8
XFILLER_24_350 VDD VSS sg13g2_decap_8
Xoutputs\[2\].output_pad _78_/Q IOVDD IOVSS output_PAD[2] VDD VSS sg13g2_IOPadOut30mA
XFILLER_12_567 VDD VSS sg13g2_decap_8
XFILLER_61_77 VDD VSS sg13g2_decap_8
XFILLER_4_700 VDD VSS sg13g2_decap_8
XFILLER_6_28 VDD VSS sg13g2_decap_8
XFILLER_3_210 VDD VSS sg13g2_decap_8
XFILLER_3_287 VDD VSS sg13g2_decap_8
XFILLER_10_70 VDD VSS sg13g2_decap_8
XFILLER_79_567 VDD VSS sg13g2_decap_8
XFILLER_94_504 VDD VSS sg13g2_decap_8
XFILLER_66_217 VDD VSS sg13g2_decap_8
XFILLER_86_63 VDD VSS sg13g2_decap_8
XFILLER_47_420 VDD VSS sg13g2_decap_8
XFILLER_59_280 VDD VSS sg13g2_decap_8
XFILLER_74_250 VDD VSS sg13g2_fill_2
XFILLER_19_133 VDD VSS sg13g2_decap_8
XFILLER_90_721 VDD VSS sg13g2_decap_8
XFILLER_74_272 VDD VSS sg13g2_decap_8
XFILLER_47_497 VDD VSS sg13g2_decap_8
XFILLER_35_637 VDD VSS sg13g2_decap_8
XFILLER_62_434 VDD VSS sg13g2_decap_8
XFILLER_34_147 VDD VSS sg13g2_decap_8
XFILLER_15_350 VDD VSS sg13g2_decap_8
XFILLER_30_364 VDD VSS sg13g2_decap_8
XFILLER_7_560 VDD VSS sg13g2_decap_8
XFILLER_58_707 VDD VSS sg13g2_decap_8
XFILLER_32_0 VDD VSS sg13g2_decap_8
XFILLER_85_504 VDD VSS sg13g2_decap_8
XFILLER_57_217 VDD VSS sg13g2_decap_8
XFILLER_38_420 VDD VSS sg13g2_decap_8
XFILLER_66_751 VDD VSS sg13g2_decap_4
XFILLER_93_581 VDD VSS sg13g2_decap_8
XFILLER_81_721 VDD VSS sg13g2_decap_8
XFILLER_26_615 VDD VSS sg13g2_decap_8
XFILLER_38_497 VDD VSS sg13g2_decap_8
XFILLER_80_231 VDD VSS sg13g2_decap_8
XFILLER_65_294 VDD VSS sg13g2_decap_8
XFILLER_25_147 VDD VSS sg13g2_decap_8
XFILLER_53_434 VDD VSS sg13g2_decap_8
XFILLER_21_364 VDD VSS sg13g2_decap_8
XFILLER_31_14 VDD VSS sg13g2_decap_8
XFILLER_1_714 VDD VSS sg13g2_decap_8
XFILLER_49_707 VDD VSS sg13g2_decap_8
XFILLER_0_224 VDD VSS sg13g2_decap_8
XFILLER_88_364 VDD VSS sg13g2_decap_8
XFILLER_48_217 VDD VSS sg13g2_decap_8
XFILLER_76_559 VDD VSS sg13g2_decap_8
XFILLER_29_420 VDD VSS sg13g2_decap_8
XFILLER_91_518 VDD VSS sg13g2_decap_8
XFILLER_84_581 VDD VSS sg13g2_decap_8
XFILLER_56_77 VDD VSS sg13g2_decap_8
XFILLER_17_637 VDD VSS sg13g2_decap_8
XFILLER_29_497 VDD VSS sg13g2_decap_8
XFILLER_72_754 VDD VSS sg13g2_fill_2
XFILLER_71_242 VDD VSS sg13g2_decap_8
XFILLER_16_147 VDD VSS sg13g2_decap_8
XFILLER_44_434 VDD VSS sg13g2_decap_8
XFILLER_56_294 VDD VSS sg13g2_decap_8
XFILLER_72_21 VDD VSS sg13g2_decap_8
XFILLER_72_98 VDD VSS sg13g2_decap_8
XFILLER_40_651 VDD VSS sg13g2_decap_8
XFILLER_12_364 VDD VSS sg13g2_decap_8
XFILLER_8_357 VDD VSS sg13g2_decap_8
XFILLER_21_91 VDD VSS sg13g2_decap_8
XFILLER_4_574 VDD VSS sg13g2_decap_8
XFILLER_94_301 VDD VSS sg13g2_decap_8
XFILLER_79_364 VDD VSS sg13g2_decap_8
XFILLER_67_548 VDD VSS sg13g2_decap_8
XFILLER_39_217 VDD VSS sg13g2_decap_8
XFILLER_82_518 VDD VSS sg13g2_decap_8
XFILLER_94_378 VDD VSS sg13g2_decap_8
XFILLER_75_592 VDD VSS sg13g2_decap_8
XFILLER_63_732 VDD VSS sg13g2_decap_8
XFILLER_62_231 VDD VSS sg13g2_decap_8
XFILLER_35_434 VDD VSS sg13g2_decap_8
XFILLER_47_294 VDD VSS sg13g2_decap_8
XFILLER_90_595 VDD VSS sg13g2_decap_8
XFILLER_50_448 VDD VSS sg13g2_decap_8
XFILLER_31_651 VDD VSS sg13g2_decap_8
XFILLER_30_161 VDD VSS sg13g2_decap_8
XFILLER_85_301 VDD VSS sg13g2_decap_8
XFILLER_58_504 VDD VSS sg13g2_decap_8
XFILLER_85_378 VDD VSS sg13g2_decap_8
XFILLER_54_721 VDD VSS sg13g2_decap_8
XFILLER_26_14 VDD VSS sg13g2_decap_8
XFILLER_26_412 VDD VSS sg13g2_decap_8
XFILLER_38_294 VDD VSS sg13g2_decap_8
XFILLER_53_231 VDD VSS sg13g2_decap_8
XFILLER_26_489 VDD VSS sg13g2_decap_8
XFILLER_81_595 VDD VSS sg13g2_decap_8
XFILLER_41_448 VDD VSS sg13g2_decap_8
XFILLER_42_35 VDD VSS sg13g2_decap_8
XFILLER_22_651 VDD VSS sg13g2_decap_8
XFILLER_21_161 VDD VSS sg13g2_decap_8
XFILLER_1_511 VDD VSS sg13g2_decap_8
XFILLER_89_651 VDD VSS sg13g2_decap_8
XFILLER_67_21 VDD VSS sg13g2_decap_8
XFILLER_49_504 VDD VSS sg13g2_decap_8
XFILLER_88_161 VDD VSS sg13g2_decap_8
XFILLER_76_334 VDD VSS sg13g2_decap_8
XFILLER_1_588 VDD VSS sg13g2_decap_8
XIO_BOND_inputs\[3\].input_pad input_PAD[3] bondpad_70x70_novias
XFILLER_67_98 VDD VSS sg13g2_decap_8
XFILLER_64_518 VDD VSS sg13g2_decap_8
XFILLER_91_315 VDD VSS sg13g2_decap_8
XFILLER_57_581 VDD VSS sg13g2_decap_8
XFILLER_45_721 VDD VSS sg13g2_decap_8
XFILLER_83_42 VDD VSS sg13g2_decap_8
XFILLER_17_434 VDD VSS sg13g2_decap_8
XFILLER_29_294 VDD VSS sg13g2_decap_8
XFILLER_44_231 VDD VSS sg13g2_decap_8
XFILLER_72_551 VDD VSS sg13g2_decap_8
XFILLER_60_735 VDD VSS sg13g2_decap_8
XFILLER_32_448 VDD VSS sg13g2_decap_8
XFILLER_13_651 VDD VSS sg13g2_decap_8
XFILLER_16_91 VDD VSS sg13g2_decap_8
XFILLER_9_644 VDD VSS sg13g2_decap_8
XFILLER_12_161 VDD VSS sg13g2_decap_8
XFILLER_73_7 VDD VSS sg13g2_decap_8
XFILLER_8_154 VDD VSS sg13g2_decap_8
XFILLER_4_371 VDD VSS sg13g2_decap_8
XFILLER_79_161 VDD VSS sg13g2_decap_8
XFILLER_95_665 VDD VSS sg13g2_decap_8
XFILLER_67_345 VDD VSS sg13g2_decap_8
XFILLER_94_175 VDD VSS sg13g2_decap_8
XFILLER_82_315 VDD VSS sg13g2_decap_8
XFILLER_55_518 VDD VSS sg13g2_decap_8
XFILLER_48_581 VDD VSS sg13g2_decap_8
XFILLER_36_721 VDD VSS sg13g2_decap_8
XFILLER_35_231 VDD VSS sg13g2_decap_8
XFILLER_90_392 VDD VSS sg13g2_decap_8
XFILLER_51_735 VDD VSS sg13g2_decap_8
XFILLER_23_448 VDD VSS sg13g2_decap_8
XFILLER_50_245 VDD VSS sg13g2_decap_8
XFILLER_12_49 VDD VSS sg13g2_decap_8
XFILLER_2_308 VDD VSS sg13g2_decap_8
XFILLER_58_301 VDD VSS sg13g2_decap_8
XFILLER_86_665 VDD VSS sg13g2_decap_8
XFILLER_85_175 VDD VSS sg13g2_decap_8
XFILLER_73_304 VDD VSS sg13g2_decap_8
XFILLER_46_518 VDD VSS sg13g2_decap_8
XFILLER_37_35 VDD VSS sg13g2_decap_8
XFILLER_58_378 VDD VSS sg13g2_decap_8
XFILLER_27_721 VDD VSS sg13g2_decap_8
XFILLER_39_581 VDD VSS sg13g2_decap_8
XFILLER_26_231 VDD VSS sg13g2_decap_8
XFILLER_81_392 VDD VSS sg13g2_decap_8
XFILLER_54_595 VDD VSS sg13g2_decap_8
XFILLER_42_735 VDD VSS sg13g2_decap_8
XFILLER_53_56 VDD VSS sg13g2_decap_8
XFILLER_14_448 VDD VSS sg13g2_decap_8
XFILLER_41_245 VDD VSS sg13g2_decap_8
XFILLER_10_665 VDD VSS sg13g2_decap_8
XFILLER_6_658 VDD VSS sg13g2_decap_8
XFILLER_5_168 VDD VSS sg13g2_decap_8
XFILLER_78_42 VDD VSS sg13g2_decap_8
XFILLER_77_632 VDD VSS sg13g2_decap_8
XFILLER_1_385 VDD VSS sg13g2_decap_8
XFILLER_49_301 VDD VSS sg13g2_decap_8
X_60_ _60_/A _60_/B _60_/C _60_/D _68_/D VDD VSS sg13g2_nor4_1
XFILLER_92_602 VDD VSS sg13g2_decap_8
XFILLER_76_175 VDD VSS sg13g2_decap_8
XFILLER_64_315 VDD VSS sg13g2_decap_8
XFILLER_94_63 VDD VSS sg13g2_decap_8
XFILLER_49_378 VDD VSS sg13g2_decap_8
XFILLER_37_518 VDD VSS sg13g2_decap_8
XFILLER_91_112 VDD VSS sg13g2_decap_8
XFILLER_18_721 VDD VSS sg13g2_decap_8
XFILLER_92_679 VDD VSS sg13g2_decap_8
XFILLER_17_231 VDD VSS sg13g2_decap_8
XFILLER_91_189 VDD VSS sg13g2_decap_8
XFILLER_72_381 VDD VSS sg13g2_decap_8
XFILLER_60_532 VDD VSS sg13g2_decap_8
XFILLER_33_735 VDD VSS sg13g2_decap_8
XFILLER_45_595 VDD VSS sg13g2_decap_8
XFILLER_32_245 VDD VSS sg13g2_decap_8
XFILLER_9_441 VDD VSS sg13g2_decap_8
XFILLER_68_643 VDD VSS sg13g2_decap_8
XFILLER_83_602 VDD VSS sg13g2_decap_8
XFILLER_95_462 VDD VSS sg13g2_decap_8
XFILLER_67_175 VDD VSS sg13g2_decap_8
XFILLER_55_315 VDD VSS sg13g2_decap_8
XFILLER_28_518 VDD VSS sg13g2_decap_8
XFILLER_82_112 VDD VSS sg13g2_decap_8
XFILLER_83_679 VDD VSS sg13g2_decap_8
XFILLER_82_189 VDD VSS sg13g2_decap_8
XFILLER_51_532 VDD VSS sg13g2_decap_8
XFILLER_24_735 VDD VSS sg13g2_decap_8
XFILLER_36_595 VDD VSS sg13g2_decap_8
XFILLER_63_392 VDD VSS sg13g2_decap_8
XFILLER_23_245 VDD VSS sg13g2_decap_8
Xoutputs\[7\].output_pad _83_/Q IOVDD IOVSS output_PAD[7] VDD VSS sg13g2_IOPadOut30mA
XFILLER_2_105 VDD VSS sg13g2_decap_8
XFILLER_3_7 VDD VSS sg13g2_decap_8
XFILLER_59_665 VDD VSS sg13g2_decap_8
XFILLER_48_56 VDD VSS sg13g2_decap_8
XFILLER_74_602 VDD VSS sg13g2_decap_8
XFILLER_86_462 VDD VSS sg13g2_decap_8
XFILLER_46_315 VDD VSS sg13g2_decap_8
XFILLER_58_175 VDD VSS sg13g2_decap_8
XFILLER_19_518 VDD VSS sg13g2_decap_8
XFILLER_73_112 VDD VSS sg13g2_decap_8
XFILLER_74_679 VDD VSS sg13g2_decap_8
XFILLER_73_189 VDD VSS sg13g2_decap_8
XFILLER_64_77 VDD VSS sg13g2_decap_8
XFILLER_61_329 VDD VSS sg13g2_decap_8
XFILLER_15_735 VDD VSS sg13g2_decap_8
XFILLER_27_595 VDD VSS sg13g2_decap_8
XFILLER_14_245 VDD VSS sg13g2_decap_8
XFILLER_54_392 VDD VSS sg13g2_decap_8
XFILLER_42_532 VDD VSS sg13g2_decap_8
XFILLER_80_21 VDD VSS sg13g2_decap_8
XFILLER_9_28 VDD VSS sg13g2_decap_8
XFILLER_30_749 VDD VSS sg13g2_decap_8
XFILLER_80_98 VDD VSS sg13g2_decap_8
XFILLER_10_462 VDD VSS sg13g2_decap_8
XFILLER_13_70 VDD VSS sg13g2_decap_8
XFILLER_6_455 VDD VSS sg13g2_decap_8
XFILLER_89_63 VDD VSS sg13g2_decap_8
XFILLER_69_429 VDD VSS sg13g2_decap_8
XFILLER_2_672 VDD VSS sg13g2_decap_8
XFILLER_36_7 VDD VSS sg13g2_decap_8
XFILLER_1_182 VDD VSS sg13g2_decap_8
X_43_ VDD _74_/A _43_/A VSS sg13g2_inv_1
XFILLER_37_315 VDD VSS sg13g2_decap_8
XFILLER_49_175 VDD VSS sg13g2_decap_8
XFILLER_64_112 VDD VSS sg13g2_decap_8
XFILLER_80_616 VDD VSS sg13g2_decap_8
XFILLER_65_668 VDD VSS sg13g2_decap_8
XFILLER_92_476 VDD VSS sg13g2_decap_8
XFILLER_64_189 VDD VSS sg13g2_decap_8
XFILLER_52_329 VDD VSS sg13g2_decap_8
XFILLER_18_595 VDD VSS sg13g2_decap_8
XFILLER_45_392 VDD VSS sg13g2_decap_8
XFILLER_33_532 VDD VSS sg13g2_decap_8
XFILLER_21_749 VDD VSS sg13g2_decap_8
XFILLER_20_259 VDD VSS sg13g2_decap_8
XFILLER_62_0 VDD VSS sg13g2_decap_8
XFILLER_0_609 VDD VSS sg13g2_decap_8
XFILLER_88_749 VDD VSS sg13g2_decap_8
XFILLER_87_259 VDD VSS sg13g2_decap_8
XFILLER_68_440 VDD VSS sg13g2_decap_8
XFILLER_56_602 VDD VSS sg13g2_decap_8
XFILLER_28_315 VDD VSS sg13g2_decap_8
XFILLER_55_112 VDD VSS sg13g2_decap_8
XFILLER_83_476 VDD VSS sg13g2_decap_8
XFILLER_56_679 VDD VSS sg13g2_decap_8
XFILLER_70_126 VDD VSS sg13g2_decap_8
XFILLER_43_329 VDD VSS sg13g2_decap_8
XFILLER_55_189 VDD VSS sg13g2_decap_8
XFILLER_34_14 VDD VSS sg13g2_decap_8
XFILLER_36_392 VDD VSS sg13g2_decap_8
XFILLER_24_532 VDD VSS sg13g2_decap_8
XFILLER_12_749 VDD VSS sg13g2_decap_8
XFILLER_11_259 VDD VSS sg13g2_decap_8
XFILLER_50_35 VDD VSS sg13g2_decap_8
XFILLER_3_469 VDD VSS sg13g2_decap_8
XFILLER_79_749 VDD VSS sg13g2_decap_8
XFILLER_59_77 VDD VSS sg13g2_decap_8
XFILLER_78_259 VDD VSS sg13g2_decap_8
XFILLER_75_21 VDD VSS sg13g2_decap_8
XFILLER_47_602 VDD VSS sg13g2_decap_8
XFILLER_59_462 VDD VSS sg13g2_decap_8
XFILLER_19_315 VDD VSS sg13g2_decap_8
XFILLER_46_112 VDD VSS sg13g2_decap_8
XFILLER_62_616 VDD VSS sg13g2_decap_8
XFILLER_74_476 VDD VSS sg13g2_decap_8
XFILLER_47_679 VDD VSS sg13g2_decap_8
XFILLER_34_329 VDD VSS sg13g2_decap_8
XFILLER_46_189 VDD VSS sg13g2_decap_8
XFILLER_61_126 VDD VSS sg13g2_decap_8
XFILLER_91_42 VDD VSS sg13g2_decap_8
XFILLER_27_392 VDD VSS sg13g2_decap_8
XFILLER_15_532 VDD VSS sg13g2_decap_8
XFILLER_30_546 VDD VSS sg13g2_decap_8
XFILLER_24_91 VDD VSS sg13g2_decap_8
XFILLER_7_742 VDD VSS sg13g2_decap_8
XFILLER_6_252 VDD VSS sg13g2_decap_8
XFILLER_38_602 VDD VSS sg13g2_decap_8
XFILLER_77_281 VDD VSS sg13g2_decap_8
XFILLER_37_112 VDD VSS sg13g2_decap_8
XFILLER_38_679 VDD VSS sg13g2_decap_8
XFILLER_92_273 VDD VSS sg13g2_decap_8
XFILLER_80_413 VDD VSS sg13g2_decap_8
XFILLER_53_616 VDD VSS sg13g2_decap_8
XFILLER_1_84 VDD VSS sg13g2_decap_8
XFILLER_25_329 VDD VSS sg13g2_decap_8
XFILLER_37_189 VDD VSS sg13g2_decap_8
XFILLER_18_392 VDD VSS sg13g2_decap_8
XFILLER_52_126 VDD VSS sg13g2_decap_8
XFILLER_61_693 VDD VSS sg13g2_decap_8
XFILLER_21_546 VDD VSS sg13g2_decap_8
XFILLER_20_49 VDD VSS sg13g2_decap_8
XFILLER_0_406 VDD VSS sg13g2_decap_8
XFILLER_88_546 VDD VSS sg13g2_decap_8
Xhold14 hold14/A VDD VSS _52_/A sg13g2_dlygate4sd3_1
XFILLER_29_14 VDD VSS sg13g2_decap_8
XFILLER_75_207 VDD VSS sg13g2_decap_8
Xhold25 _78_/Q VDD VSS _59_/A sg13g2_dlygate4sd3_1
XFILLER_29_602 VDD VSS sg13g2_decap_8
XFILLER_28_112 VDD VSS sg13g2_decap_8
XFILLER_29_679 VDD VSS sg13g2_decap_8
XFILLER_83_273 VDD VSS sg13g2_decap_8
XFILLER_45_35 VDD VSS sg13g2_decap_8
XFILLER_16_329 VDD VSS sg13g2_decap_8
XFILLER_28_189 VDD VSS sg13g2_decap_8
XFILLER_56_476 VDD VSS sg13g2_decap_8
XFILLER_44_616 VDD VSS sg13g2_decap_8
XFILLER_71_457 VDD VSS sg13g2_decap_8
XFILLER_43_126 VDD VSS sg13g2_decap_8
XFILLER_52_693 VDD VSS sg13g2_decap_8
XFILLER_12_546 VDD VSS sg13g2_decap_8
XFILLER_61_56 VDD VSS sg13g2_decap_8
XFILLER_8_539 VDD VSS sg13g2_decap_8
XFILLER_4_756 VDD VSS sg13g2_fill_1
XFILLER_3_266 VDD VSS sg13g2_decap_8
XFILLER_79_546 VDD VSS sg13g2_decap_8
XFILLER_86_42 VDD VSS sg13g2_decap_8
XFILLER_19_112 VDD VSS sg13g2_decap_8
XFILLER_90_700 VDD VSS sg13g2_decap_8
XFILLER_19_91 VDD VSS sg13g2_decap_8
XFILLER_62_413 VDD VSS sg13g2_decap_8
XFILLER_19_189 VDD VSS sg13g2_decap_8
XFILLER_47_476 VDD VSS sg13g2_decap_8
XFILLER_35_616 VDD VSS sg13g2_decap_8
XFILLER_62_457 VDD VSS sg13g2_fill_1
XFILLER_34_126 VDD VSS sg13g2_decap_8
XFILLER_43_693 VDD VSS sg13g2_decap_8
XFILLER_30_343 VDD VSS sg13g2_decap_8
XFILLER_25_0 VDD VSS sg13g2_decap_8
XFILLER_66_730 VDD VSS sg13g2_decap_8
XFILLER_93_560 VDD VSS sg13g2_decap_8
XFILLER_81_700 VDD VSS sg13g2_decap_8
XFILLER_65_273 VDD VSS sg13g2_decap_8
XFILLER_38_476 VDD VSS sg13g2_decap_8
XFILLER_53_413 VDD VSS sg13g2_decap_8
XFILLER_80_210 VDD VSS sg13g2_decap_8
XFILLER_25_126 VDD VSS sg13g2_decap_8
XFILLER_80_287 VDD VSS sg13g2_decap_8
XFILLER_61_490 VDD VSS sg13g2_decap_8
XFILLER_15_49 VDD VSS sg13g2_decap_8
XFILLER_34_693 VDD VSS sg13g2_decap_8
XFILLER_21_343 VDD VSS sg13g2_decap_8
XFILLER_0_203 VDD VSS sg13g2_decap_8
XFILLER_88_343 VDD VSS sg13g2_decap_8
XIO_BOND_inputs\[2\].input_pad input_PAD[2] bondpad_70x70_novias
XFILLER_76_538 VDD VSS sg13g2_decap_8
XFILLER_56_56 VDD VSS sg13g2_decap_8
XFILLER_84_560 VDD VSS sg13g2_decap_8
XFILLER_29_476 VDD VSS sg13g2_decap_8
XFILLER_44_413 VDD VSS sg13g2_decap_8
XFILLER_56_273 VDD VSS sg13g2_decap_8
XFILLER_17_616 VDD VSS sg13g2_decap_8
XFILLER_72_733 VDD VSS sg13g2_decap_8
XFILLER_71_210 VDD VSS sg13g2_fill_2
XFILLER_16_126 VDD VSS sg13g2_decap_8
XFILLER_72_77 VDD VSS sg13g2_decap_8
XFILLER_52_490 VDD VSS sg13g2_decap_8
XFILLER_25_693 VDD VSS sg13g2_decap_8
XFILLER_40_630 VDD VSS sg13g2_decap_8
XFILLER_12_343 VDD VSS sg13g2_decap_8
XFILLER_8_336 VDD VSS sg13g2_decap_8
XFILLER_21_70 VDD VSS sg13g2_decap_8
XFILLER_4_553 VDD VSS sg13g2_decap_8
XFILLER_79_343 VDD VSS sg13g2_decap_8
XFILLER_67_527 VDD VSS sg13g2_decap_8
XFILLER_94_357 VDD VSS sg13g2_decap_8
XFILLER_75_571 VDD VSS sg13g2_decap_8
XFILLER_63_711 VDD VSS sg13g2_decap_8
XFILLER_35_413 VDD VSS sg13g2_decap_8
XFILLER_47_273 VDD VSS sg13g2_decap_8
XFILLER_62_210 VDD VSS sg13g2_decap_8
XFILLER_90_574 VDD VSS sg13g2_decap_8
XFILLER_62_287 VDD VSS sg13g2_decap_8
XFILLER_50_427 VDD VSS sg13g2_decap_8
XFILLER_16_693 VDD VSS sg13g2_decap_8
XFILLER_31_630 VDD VSS sg13g2_decap_8
XFILLER_43_490 VDD VSS sg13g2_decap_8
XFILLER_30_140 VDD VSS sg13g2_decap_8
XIO_CORNER_NORTH_EAST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XFILLER_85_357 VDD VSS sg13g2_decap_8
XFILLER_54_700 VDD VSS sg13g2_decap_8
XFILLER_38_273 VDD VSS sg13g2_decap_8
XFILLER_53_210 VDD VSS sg13g2_decap_8
XFILLER_81_574 VDD VSS sg13g2_decap_8
XFILLER_26_468 VDD VSS sg13g2_decap_8
XFILLER_41_427 VDD VSS sg13g2_decap_8
XFILLER_53_287 VDD VSS sg13g2_decap_8
XFILLER_42_14 VDD VSS sg13g2_decap_8
XFILLER_22_630 VDD VSS sg13g2_decap_8
XFILLER_34_490 VDD VSS sg13g2_decap_8
XFILLER_21_140 VDD VSS sg13g2_decap_8
XFILLER_89_630 VDD VSS sg13g2_decap_8
XFILLER_88_140 VDD VSS sg13g2_decap_8
XFILLER_1_567 VDD VSS sg13g2_decap_8
XFILLER_76_313 VDD VSS sg13g2_decap_8
XFILLER_67_77 VDD VSS sg13g2_decap_8
XFILLER_57_560 VDD VSS sg13g2_decap_8
XFILLER_17_413 VDD VSS sg13g2_decap_8
XFILLER_29_273 VDD VSS sg13g2_decap_8
XFILLER_45_700 VDD VSS sg13g2_decap_8
XFILLER_72_530 VDD VSS sg13g2_decap_8
XFILLER_83_21 VDD VSS sg13g2_decap_8
XFILLER_44_210 VDD VSS sg13g2_decap_8
XFILLER_60_714 VDD VSS sg13g2_decap_8
XFILLER_83_98 VDD VSS sg13g2_decap_8
XFILLER_16_70 VDD VSS sg13g2_decap_8
XFILLER_32_427 VDD VSS sg13g2_decap_8
XFILLER_44_287 VDD VSS sg13g2_decap_8
XFILLER_13_630 VDD VSS sg13g2_decap_8
XFILLER_25_490 VDD VSS sg13g2_decap_8
XFILLER_9_623 VDD VSS sg13g2_decap_8
XFILLER_12_140 VDD VSS sg13g2_decap_8
XFILLER_8_133 VDD VSS sg13g2_decap_8
XFILLER_66_7 VDD VSS sg13g2_decap_8
XFILLER_32_91 VDD VSS sg13g2_decap_8
XFILLER_4_350 VDD VSS sg13g2_decap_8
XFILLER_79_140 VDD VSS sg13g2_decap_8
XFILLER_67_324 VDD VSS sg13g2_decap_8
XFILLER_95_644 VDD VSS sg13g2_decap_8
XFILLER_94_154 VDD VSS sg13g2_decap_8
XFILLER_48_560 VDD VSS sg13g2_decap_8
XFILLER_36_700 VDD VSS sg13g2_decap_8
XFILLER_35_210 VDD VSS sg13g2_decap_8
XFILLER_51_714 VDD VSS sg13g2_decap_8
XFILLER_63_585 VDD VSS sg13g2_decap_8
XFILLER_90_371 VDD VSS sg13g2_decap_8
XFILLER_23_427 VDD VSS sg13g2_decap_8
XFILLER_35_287 VDD VSS sg13g2_decap_8
XFILLER_50_224 VDD VSS sg13g2_decap_8
XFILLER_92_0 VDD VSS sg13g2_decap_8
XFILLER_16_490 VDD VSS sg13g2_decap_8
XFILLER_12_28 VDD VSS sg13g2_decap_8
XFILLER_86_644 VDD VSS sg13g2_decap_8
XFILLER_37_14 VDD VSS sg13g2_decap_8
XFILLER_58_357 VDD VSS sg13g2_decap_8
XFILLER_85_154 VDD VSS sg13g2_decap_8
XFILLER_27_700 VDD VSS sg13g2_decap_8
XFILLER_39_560 VDD VSS sg13g2_decap_8
XFILLER_26_210 VDD VSS sg13g2_decap_8
XFILLER_42_714 VDD VSS sg13g2_decap_8
XFILLER_81_371 VDD VSS sg13g2_decap_8
XFILLER_54_574 VDD VSS sg13g2_decap_8
XFILLER_53_35 VDD VSS sg13g2_decap_8
XFILLER_14_427 VDD VSS sg13g2_decap_8
XFILLER_26_287 VDD VSS sg13g2_decap_4
XFILLER_41_224 VDD VSS sg13g2_decap_8
XFILLER_10_644 VDD VSS sg13g2_decap_8
XFILLER_6_637 VDD VSS sg13g2_decap_8
XFILLER_5_147 VDD VSS sg13g2_decap_8
XFILLER_78_21 VDD VSS sg13g2_decap_8
XFILLER_77_611 VDD VSS sg13g2_decap_8
XFILLER_78_98 VDD VSS sg13g2_decap_8
XFILLER_1_364 VDD VSS sg13g2_decap_8
XFILLER_49_357 VDD VSS sg13g2_decap_8
XFILLER_77_688 VDD VSS sg13g2_decap_8
XFILLER_76_154 VDD VSS sg13g2_decap_8
XFILLER_94_42 VDD VSS sg13g2_decap_8
XFILLER_18_700 VDD VSS sg13g2_decap_8
XFILLER_92_658 VDD VSS sg13g2_decap_8
XFILLER_17_210 VDD VSS sg13g2_decap_8
XFILLER_91_168 VDD VSS sg13g2_decap_8
XFILLER_60_511 VDD VSS sg13g2_decap_8
XFILLER_27_91 VDD VSS sg13g2_decap_8
XFILLER_17_287 VDD VSS sg13g2_decap_8
XFILLER_33_714 VDD VSS sg13g2_decap_8
XFILLER_45_574 VDD VSS sg13g2_decap_8
XFILLER_32_224 VDD VSS sg13g2_decap_8
XFILLER_60_588 VDD VSS sg13g2_decap_8
XFILLER_9_420 VDD VSS sg13g2_decap_8
XFILLER_9_497 VDD VSS sg13g2_decap_8
XFILLER_68_622 VDD VSS sg13g2_decap_8
XFILLER_4_84 VDD VSS sg13g2_decap_8
XFILLER_95_441 VDD VSS sg13g2_decap_8
XFILLER_68_699 VDD VSS sg13g2_decap_8
XFILLER_67_154 VDD VSS sg13g2_decap_8
XFILLER_83_658 VDD VSS sg13g2_decap_8
XFILLER_82_168 VDD VSS sg13g2_decap_8
XFILLER_63_371 VDD VSS sg13g2_decap_8
XFILLER_51_511 VDD VSS sg13g2_decap_8
XFILLER_24_714 VDD VSS sg13g2_decap_8
XFILLER_36_574 VDD VSS sg13g2_decap_8
XFILLER_23_224 VDD VSS sg13g2_decap_8
XFILLER_51_588 VDD VSS sg13g2_decap_8
XFILLER_23_49 VDD VSS sg13g2_decap_8
XFILLER_86_441 VDD VSS sg13g2_decap_8
XFILLER_59_644 VDD VSS sg13g2_decap_8
XFILLER_48_35 VDD VSS sg13g2_decap_8
XFILLER_58_154 VDD VSS sg13g2_decap_8
XFILLER_74_658 VDD VSS sg13g2_decap_8
XFILLER_73_168 VDD VSS sg13g2_decap_8
XFILLER_61_308 VDD VSS sg13g2_decap_8
XFILLER_64_56 VDD VSS sg13g2_decap_8
XFILLER_54_371 VDD VSS sg13g2_decap_8
XFILLER_15_714 VDD VSS sg13g2_decap_8
XFILLER_27_574 VDD VSS sg13g2_decap_8
XFILLER_42_511 VDD VSS sg13g2_decap_8
XFILLER_14_224 VDD VSS sg13g2_decap_8
XFILLER_30_728 VDD VSS sg13g2_decap_8
XFILLER_42_588 VDD VSS sg13g2_decap_8
XFILLER_80_77 VDD VSS sg13g2_decap_8
XFILLER_10_441 VDD VSS sg13g2_decap_8
XFILLER_6_434 VDD VSS sg13g2_decap_8
XFILLER_89_42 VDD VSS sg13g2_decap_8
XFILLER_69_408 VDD VSS sg13g2_decap_8
XFILLER_2_651 VDD VSS sg13g2_decap_8
XFILLER_1_161 VDD VSS sg13g2_decap_8
XFILLER_29_7 VDD VSS sg13g2_decap_8
XFILLER_49_154 VDD VSS sg13g2_decap_8
XFILLER_77_485 VDD VSS sg13g2_decap_8
XFILLER_65_647 VDD VSS sg13g2_decap_8
XFILLER_92_455 VDD VSS sg13g2_decap_8
XFILLER_64_168 VDD VSS sg13g2_decap_8
XFILLER_52_308 VDD VSS sg13g2_decap_8
XFILLER_45_371 VDD VSS sg13g2_decap_8
XFILLER_18_574 VDD VSS sg13g2_decap_8
XFILLER_33_511 VDD VSS sg13g2_decap_8
XFILLER_21_728 VDD VSS sg13g2_decap_8
XFILLER_33_588 VDD VSS sg13g2_decap_8
XFILLER_20_238 VDD VSS sg13g2_decap_8
XFILLER_60_385 VDD VSS sg13g2_decap_8
XFILLER_9_294 VDD VSS sg13g2_decap_8
XFILLER_55_0 VDD VSS sg13g2_decap_8
XFILLER_88_728 VDD VSS sg13g2_decap_8
XFILLER_87_238 VDD VSS sg13g2_decap_8
XFILLER_68_496 VDD VSS sg13g2_decap_8
XFILLER_18_49 VDD VSS sg13g2_decap_8
XFILLER_83_455 VDD VSS sg13g2_decap_8
XFILLER_56_658 VDD VSS sg13g2_decap_8
XFILLER_43_308 VDD VSS sg13g2_decap_8
XFILLER_71_639 VDD VSS sg13g2_decap_8
XFILLER_70_105 VDD VSS sg13g2_decap_8
XFILLER_36_371 VDD VSS sg13g2_decap_8
XFILLER_55_168 VDD VSS sg13g2_decap_8
XFILLER_24_511 VDD VSS sg13g2_decap_8
XFILLER_12_728 VDD VSS sg13g2_decap_8
XFILLER_24_588 VDD VSS sg13g2_decap_8
XFILLER_11_238 VDD VSS sg13g2_decap_8
XFILLER_51_385 VDD VSS sg13g2_decap_8
XFILLER_50_14 VDD VSS sg13g2_decap_8
XFILLER_3_448 VDD VSS sg13g2_decap_8
XFILLER_79_728 VDD VSS sg13g2_decap_8
XFILLER_59_56 VDD VSS sg13g2_decap_8
XFILLER_78_238 VDD VSS sg13g2_decap_8
XFILLER_59_441 VDD VSS sg13g2_decap_8
XFILLER_74_444 VDD VSS sg13g2_fill_1
XFILLER_74_455 VDD VSS sg13g2_decap_8
XFILLER_75_88 VDD VSS sg13g2_decap_8
XFILLER_47_658 VDD VSS sg13g2_decap_8
XFILLER_61_105 VDD VSS sg13g2_decap_8
XFILLER_27_371 VDD VSS sg13g2_decap_8
XFILLER_34_308 VDD VSS sg13g2_decap_8
XFILLER_46_168 VDD VSS sg13g2_decap_8
XFILLER_15_511 VDD VSS sg13g2_decap_8
XFILLER_91_21 VDD VSS sg13g2_decap_8
XFILLER_15_588 VDD VSS sg13g2_decap_8
XFILLER_70_694 VDD VSS sg13g2_decap_8
XFILLER_91_98 VDD VSS sg13g2_decap_8
XFILLER_42_385 VDD VSS sg13g2_decap_8
XFILLER_30_525 VDD VSS sg13g2_decap_8
XFILLER_24_70 VDD VSS sg13g2_decap_8
XFILLER_7_721 VDD VSS sg13g2_decap_8
XFILLER_6_231 VDD VSS sg13g2_decap_8
XFILLER_40_91 VDD VSS sg13g2_decap_8
XFILLER_69_238 VDD VSS sg13g2_fill_2
XFILLER_93_742 VDD VSS sg13g2_decap_8
XFILLER_77_260 VDD VSS sg13g2_decap_8
XFILLER_92_252 VDD VSS sg13g2_decap_8
XFILLER_65_455 VDD VSS sg13g2_decap_8
XFILLER_1_63 VDD VSS sg13g2_decap_8
XFILLER_38_658 VDD VSS sg13g2_decap_8
XFILLER_52_105 VDD VSS sg13g2_decap_8
XFILLER_18_371 VDD VSS sg13g2_decap_8
XFILLER_25_308 VDD VSS sg13g2_decap_8
XFILLER_37_168 VDD VSS sg13g2_decap_8
XFILLER_80_469 VDD VSS sg13g2_decap_8
XFILLER_61_672 VDD VSS sg13g2_decap_8
XFILLER_33_385 VDD VSS sg13g2_decap_8
XFILLER_60_182 VDD VSS sg13g2_decap_8
XFILLER_21_525 VDD VSS sg13g2_decap_8
XFILLER_20_28 VDD VSS sg13g2_decap_8
XFILLER_88_525 VDD VSS sg13g2_decap_8
XIO_BOND_inputs\[1\].input_pad input_PAD[1] bondpad_70x70_novias
Xhold26 _59_/Y VDD VSS _61_/B sg13g2_dlygate4sd3_1
Xhold15 _49_/Y VDD VSS _60_/C sg13g2_dlygate4sd3_1
XFILLER_84_742 VDD VSS sg13g2_decap_8
XFILLER_68_293 VDD VSS sg13g2_decap_8
XFILLER_56_455 VDD VSS sg13g2_decap_8
XFILLER_29_658 VDD VSS sg13g2_decap_8
XFILLER_83_252 VDD VSS sg13g2_decap_8
XFILLER_43_105 VDD VSS sg13g2_decap_8
XFILLER_45_14 VDD VSS sg13g2_decap_8
XFILLER_16_308 VDD VSS sg13g2_decap_8
XFILLER_28_168 VDD VSS sg13g2_decap_8
XFILLER_71_436 VDD VSS sg13g2_decap_8
XFILLER_52_672 VDD VSS sg13g2_decap_8
XFILLER_12_525 VDD VSS sg13g2_decap_8
XFILLER_24_385 VDD VSS sg13g2_decap_8
XFILLER_51_182 VDD VSS sg13g2_decap_8
XFILLER_8_518 VDD VSS sg13g2_decap_8
XFILLER_61_35 VDD VSS sg13g2_decap_8
XFILLER_4_735 VDD VSS sg13g2_decap_8
XFILLER_3_245 VDD VSS sg13g2_decap_8
XFILLER_79_525 VDD VSS sg13g2_decap_8
XFILLER_86_21 VDD VSS sg13g2_decap_8
XFILLER_67_709 VDD VSS sg13g2_decap_8
XFILLER_94_539 VDD VSS sg13g2_decap_8
XFILLER_86_98 VDD VSS sg13g2_decap_8
XFILLER_75_753 VDD VSS sg13g2_decap_4
XFILLER_19_70 VDD VSS sg13g2_decap_8
XFILLER_47_455 VDD VSS sg13g2_decap_8
XFILLER_74_252 VDD VSS sg13g2_fill_1
XFILLER_34_105 VDD VSS sg13g2_decap_8
XFILLER_19_168 VDD VSS sg13g2_decap_8
XFILLER_90_756 VDD VSS sg13g2_fill_1
XFILLER_62_469 VDD VSS sg13g2_decap_8
XFILLER_50_609 VDD VSS sg13g2_decap_8
XFILLER_43_672 VDD VSS sg13g2_decap_8
XFILLER_70_491 VDD VSS sg13g2_decap_8
XFILLER_70_480 VDD VSS sg13g2_fill_1
XFILLER_35_91 VDD VSS sg13g2_decap_8
XFILLER_15_385 VDD VSS sg13g2_decap_8
XFILLER_30_322 VDD VSS sg13g2_decap_8
XFILLER_42_182 VDD VSS sg13g2_decap_8
XFILLER_30_399 VDD VSS sg13g2_decap_8
XFILLER_7_595 VDD VSS sg13g2_decap_8
XFILLER_85_539 VDD VSS sg13g2_decap_8
XFILLER_18_0 VDD VSS sg13g2_decap_8
XFILLER_38_455 VDD VSS sg13g2_decap_8
XFILLER_65_252 VDD VSS sg13g2_decap_8
XFILLER_25_105 VDD VSS sg13g2_decap_8
XFILLER_81_756 VDD VSS sg13g2_fill_1
XFILLER_80_266 VDD VSS sg13g2_decap_8
XFILLER_15_28 VDD VSS sg13g2_decap_8
XFILLER_53_469 VDD VSS sg13g2_decap_8
XFILLER_41_609 VDD VSS sg13g2_decap_8
XFILLER_40_119 VDD VSS sg13g2_decap_8
XFILLER_34_672 VDD VSS sg13g2_decap_8
XFILLER_21_322 VDD VSS sg13g2_decap_8
XFILLER_33_182 VDD VSS sg13g2_decap_8
XFILLER_31_49 VDD VSS sg13g2_decap_8
XFILLER_21_399 VDD VSS sg13g2_decap_8
XFILLER_88_322 VDD VSS sg13g2_decap_8
XFILLER_1_749 VDD VSS sg13g2_decap_8
XFILLER_76_517 VDD VSS sg13g2_decap_8
XFILLER_0_259 VDD VSS sg13g2_decap_8
XFILLER_69_580 VDD VSS sg13g2_decap_8
XFILLER_88_399 VDD VSS sg13g2_decap_8
XFILLER_57_742 VDD VSS sg13g2_decap_8
XFILLER_56_35 VDD VSS sg13g2_decap_8
XFILLER_29_455 VDD VSS sg13g2_decap_8
XFILLER_72_712 VDD VSS sg13g2_decap_8
XFILLER_16_105 VDD VSS sg13g2_decap_8
XFILLER_56_252 VDD VSS sg13g2_decap_8
XFILLER_72_756 VDD VSS sg13g2_fill_1
XFILLER_71_222 VDD VSS sg13g2_fill_1
XFILLER_44_469 VDD VSS sg13g2_decap_8
XFILLER_32_609 VDD VSS sg13g2_decap_8
XFILLER_71_277 VDD VSS sg13g2_decap_8
XFILLER_72_56 VDD VSS sg13g2_decap_8
XFILLER_31_119 VDD VSS sg13g2_decap_8
XFILLER_25_672 VDD VSS sg13g2_decap_8
XFILLER_12_322 VDD VSS sg13g2_decap_8
XFILLER_24_182 VDD VSS sg13g2_decap_8
XFILLER_8_315 VDD VSS sg13g2_decap_8
XFILLER_40_686 VDD VSS sg13g2_decap_8
XFILLER_12_399 VDD VSS sg13g2_decap_8
XFILLER_4_532 VDD VSS sg13g2_decap_8
XFILLER_79_322 VDD VSS sg13g2_decap_8
XFILLER_67_506 VDD VSS sg13g2_decap_8
XFILLER_79_399 VDD VSS sg13g2_decap_8
XFILLER_94_336 VDD VSS sg13g2_decap_8
XFILLER_48_742 VDD VSS sg13g2_decap_8
XFILLER_11_7 VDD VSS sg13g2_decap_8
XFILLER_75_550 VDD VSS sg13g2_decap_8
XFILLER_47_252 VDD VSS sg13g2_decap_8
XFILLER_90_553 VDD VSS sg13g2_decap_8
XFILLER_62_266 VDD VSS sg13g2_decap_8
XFILLER_35_469 VDD VSS sg13g2_decap_8
XFILLER_50_406 VDD VSS sg13g2_decap_8
XFILLER_23_609 VDD VSS sg13g2_decap_8
XFILLER_22_119 VDD VSS sg13g2_decap_8
XFILLER_16_672 VDD VSS sg13g2_decap_8
XFILLER_15_182 VDD VSS sg13g2_decap_8
XFILLER_31_686 VDD VSS sg13g2_decap_8
XFILLER_30_196 VDD VSS sg13g2_decap_8
XFILLER_7_392 VDD VSS sg13g2_decap_8
XFILLER_7_84 VDD VSS sg13g2_decap_8
XFILLER_89_119 VDD VSS sg13g2_decap_8
XFILLER_58_539 VDD VSS sg13g2_decap_8
XFILLER_85_336 VDD VSS sg13g2_decap_8
XFILLER_39_742 VDD VSS sg13g2_decap_8
XFILLER_38_252 VDD VSS sg13g2_decap_8
XFILLER_66_583 VDD VSS sg13g2_decap_8
XFILLER_54_756 VDD VSS sg13g2_fill_1
XFILLER_26_447 VDD VSS sg13g2_decap_8
XFILLER_81_553 VDD VSS sg13g2_decap_8
XFILLER_26_49 VDD VSS sg13g2_decap_8
XFILLER_41_406 VDD VSS sg13g2_decap_8
XFILLER_53_266 VDD VSS sg13g2_decap_8
XFILLER_14_609 VDD VSS sg13g2_decap_8
XFILLER_13_119 VDD VSS sg13g2_decap_8
XFILLER_22_686 VDD VSS sg13g2_decap_8
XFILLER_21_196 VDD VSS sg13g2_decap_8
XFILLER_5_329 VDD VSS sg13g2_decap_8
XFILLER_1_546 VDD VSS sg13g2_decap_8
XFILLER_89_686 VDD VSS sg13g2_decap_8
XFILLER_67_56 VDD VSS sg13g2_decap_8
XFILLER_49_539 VDD VSS sg13g2_decap_8
XFILLER_88_196 VDD VSS sg13g2_decap_8
XFILLER_76_369 VDD VSS sg13g2_decap_8
XFILLER_29_252 VDD VSS sg13g2_decap_8
XFILLER_83_77 VDD VSS sg13g2_decap_8
XFILLER_17_469 VDD VSS sg13g2_decap_8
XFILLER_32_406 VDD VSS sg13g2_decap_8
XFILLER_45_756 VDD VSS sg13g2_fill_1
XFILLER_72_586 VDD VSS sg13g2_decap_8
XFILLER_44_266 VDD VSS sg13g2_decap_8
XFILLER_9_602 VDD VSS sg13g2_decap_8
XFILLER_13_686 VDD VSS sg13g2_decap_8
XFILLER_8_112 VDD VSS sg13g2_decap_8
XFILLER_12_196 VDD VSS sg13g2_decap_8
XFILLER_40_483 VDD VSS sg13g2_decap_8
XFILLER_9_679 VDD VSS sg13g2_decap_8
XFILLER_32_70 VDD VSS sg13g2_decap_8
XFILLER_8_189 VDD VSS sg13g2_decap_8
XFILLER_59_7 VDD VSS sg13g2_decap_8
XFILLER_95_623 VDD VSS sg13g2_decap_8
XFILLER_67_303 VDD VSS sg13g2_decap_8
XFILLER_94_133 VDD VSS sg13g2_decap_8
XFILLER_79_196 VDD VSS sg13g2_decap_8
XFILLER_63_564 VDD VSS sg13g2_decap_8
XFILLER_90_350 VDD VSS sg13g2_decap_8
XFILLER_36_756 VDD VSS sg13g2_fill_1
XFILLER_23_406 VDD VSS sg13g2_decap_8
XFILLER_35_266 VDD VSS sg13g2_decap_8
XFILLER_50_203 VDD VSS sg13g2_decap_8
XFILLER_85_0 VDD VSS sg13g2_decap_8
XFILLER_31_483 VDD VSS sg13g2_decap_8
XFILLER_86_623 VDD VSS sg13g2_decap_8
XFILLER_85_133 VDD VSS sg13g2_decap_8
XFILLER_58_336 VDD VSS sg13g2_decap_8
XFILLER_73_339 VDD VSS sg13g2_decap_4
XFILLER_81_350 VDD VSS sg13g2_decap_8
XFILLER_54_553 VDD VSS sg13g2_decap_8
XFILLER_27_756 VDD VSS sg13g2_fill_1
XFILLER_53_14 VDD VSS sg13g2_decap_8
XFILLER_14_406 VDD VSS sg13g2_decap_8
XFILLER_26_266 VDD VSS sg13g2_decap_8
XFILLER_41_203 VDD VSS sg13g2_decap_8
XFILLER_10_623 VDD VSS sg13g2_decap_8
XFILLER_22_483 VDD VSS sg13g2_decap_8
XFILLER_6_616 VDD VSS sg13g2_decap_8
XFILLER_5_126 VDD VSS sg13g2_decap_8
XFILLER_1_343 VDD VSS sg13g2_decap_8
XFILLER_89_483 VDD VSS sg13g2_decap_8
XFILLER_78_77 VDD VSS sg13g2_decap_8
XFILLER_76_133 VDD VSS sg13g2_decap_8
XFILLER_49_336 VDD VSS sg13g2_decap_8
XFILLER_77_667 VDD VSS sg13g2_decap_8
XFILLER_94_21 VDD VSS sg13g2_decap_8
XFILLER_92_637 VDD VSS sg13g2_decap_8
XFILLER_91_147 VDD VSS sg13g2_decap_8
XFILLER_94_98 VDD VSS sg13g2_decap_8
XFILLER_27_70 VDD VSS sg13g2_decap_8
XFILLER_18_756 VDD VSS sg13g2_fill_1
XFILLER_45_553 VDD VSS sg13g2_decap_8
XFILLER_17_266 VDD VSS sg13g2_decap_8
XFILLER_32_203 VDD VSS sg13g2_decap_8
X_76__3 VDD VSS _76__3/L_HI sg13g2_tiehi
XFILLER_60_567 VDD VSS sg13g2_decap_8
XFILLER_13_483 VDD VSS sg13g2_decap_8
XFILLER_43_91 VDD VSS sg13g2_decap_8
XFILLER_40_280 VDD VSS sg13g2_decap_8
XFILLER_9_476 VDD VSS sg13g2_decap_8
XFILLER_5_693 VDD VSS sg13g2_decap_8
XFILLER_68_601 VDD VSS sg13g2_decap_8
XFILLER_4_63 VDD VSS sg13g2_decap_8
XFILLER_95_420 VDD VSS sg13g2_decap_8
XFILLER_67_133 VDD VSS sg13g2_decap_8
XFILLER_68_678 VDD VSS sg13g2_decap_8
XFILLER_95_497 VDD VSS sg13g2_decap_8
XFILLER_83_637 VDD VSS sg13g2_decap_8
XFILLER_82_147 VDD VSS sg13g2_decap_8
XFILLER_36_553 VDD VSS sg13g2_decap_8
XFILLER_63_350 VDD VSS sg13g2_decap_8
XFILLER_23_203 VDD VSS sg13g2_decap_8
XFILLER_51_567 VDD VSS sg13g2_decap_8
XFILLER_23_28 VDD VSS sg13g2_decap_8
XFILLER_31_280 VDD VSS sg13g2_decap_8
XFILLER_59_623 VDD VSS sg13g2_decap_8
XFILLER_48_14 VDD VSS sg13g2_decap_8
XFILLER_86_420 VDD VSS sg13g2_decap_8
XFILLER_58_133 VDD VSS sg13g2_decap_8
XFILLER_86_497 VDD VSS sg13g2_decap_8
XFILLER_74_637 VDD VSS sg13g2_decap_8
XFILLER_73_147 VDD VSS sg13g2_decap_8
XFILLER_27_553 VDD VSS sg13g2_decap_8
XFILLER_14_203 VDD VSS sg13g2_decap_8
XFILLER_54_350 VDD VSS sg13g2_decap_8
XFILLER_30_707 VDD VSS sg13g2_decap_8
XFILLER_42_567 VDD VSS sg13g2_decap_8
XFILLER_80_56 VDD VSS sg13g2_decap_8
XFILLER_10_420 VDD VSS sg13g2_decap_8
XFILLER_22_280 VDD VSS sg13g2_decap_8
XFILLER_6_413 VDD VSS sg13g2_decap_8
XFILLER_89_21 VDD VSS sg13g2_decap_8
XFILLER_10_497 VDD VSS sg13g2_decap_8
XFILLER_89_98 VDD VSS sg13g2_decap_8
XFILLER_2_630 VDD VSS sg13g2_decap_8
XFILLER_1_140 VDD VSS sg13g2_decap_8
XFILLER_89_280 VDD VSS sg13g2_decap_8
XFILLER_77_464 VDD VSS sg13g2_decap_8
XFILLER_77_442 VDD VSS sg13g2_decap_8
XFILLER_49_133 VDD VSS sg13g2_decap_8
XFILLER_65_626 VDD VSS sg13g2_decap_8
XFILLER_92_434 VDD VSS sg13g2_decap_8
XFILLER_64_147 VDD VSS sg13g2_decap_8
XFILLER_38_91 VDD VSS sg13g2_decap_8
XFILLER_18_553 VDD VSS sg13g2_decap_8
XFILLER_73_681 VDD VSS sg13g2_decap_8
XFILLER_45_350 VDD VSS sg13g2_decap_8
XFILLER_60_364 VDD VSS sg13g2_decap_8
XFILLER_21_707 VDD VSS sg13g2_decap_8
XFILLER_33_567 VDD VSS sg13g2_decap_8
XFILLER_20_217 VDD VSS sg13g2_decap_8
XFILLER_13_280 VDD VSS sg13g2_decap_8
XFILLER_9_273 VDD VSS sg13g2_decap_8
XFILLER_88_707 VDD VSS sg13g2_decap_8
XIO_BOND_inputs\[0\].input_pad input_PAD[0] bondpad_70x70_novias
XFILLER_5_490 VDD VSS sg13g2_decap_8
XFILLER_48_0 VDD VSS sg13g2_decap_8
XFILLER_87_217 VDD VSS sg13g2_decap_8
XFILLER_83_434 VDD VSS sg13g2_decap_8
XFILLER_68_475 VDD VSS sg13g2_decap_8
XFILLER_56_637 VDD VSS sg13g2_decap_8
XFILLER_18_28 VDD VSS sg13g2_decap_8
XFILLER_95_294 VDD VSS sg13g2_decap_8
XFILLER_55_147 VDD VSS sg13g2_decap_8
XFILLER_71_618 VDD VSS sg13g2_decap_8
XFILLER_36_350 VDD VSS sg13g2_decap_8
XFILLER_12_707 VDD VSS sg13g2_decap_8
XFILLER_34_49 VDD VSS sg13g2_decap_8
XFILLER_51_364 VDD VSS sg13g2_decap_8
XFILLER_24_567 VDD VSS sg13g2_decap_8
XFILLER_11_217 VDD VSS sg13g2_decap_8
XFILLER_3_427 VDD VSS sg13g2_decap_8
XFILLER_79_707 VDD VSS sg13g2_decap_8
XFILLER_78_217 VDD VSS sg13g2_decap_8
XFILLER_59_35 VDD VSS sg13g2_decap_8
XFILLER_59_420 VDD VSS sg13g2_decap_8
XFILLER_74_423 VDD VSS sg13g2_decap_8
XFILLER_59_497 VDD VSS sg13g2_decap_8
XFILLER_47_637 VDD VSS sg13g2_decap_8
XFILLER_86_294 VDD VSS sg13g2_decap_8
XFILLER_75_67 VDD VSS sg13g2_decap_8
XFILLER_46_147 VDD VSS sg13g2_decap_8
XFILLER_27_350 VDD VSS sg13g2_decap_8
XFILLER_70_673 VDD VSS sg13g2_decap_8
XFILLER_42_364 VDD VSS sg13g2_decap_8
XFILLER_15_567 VDD VSS sg13g2_decap_8
XFILLER_30_504 VDD VSS sg13g2_decap_8
XFILLER_91_77 VDD VSS sg13g2_decap_8
XFILLER_7_700 VDD VSS sg13g2_decap_8
XFILLER_6_210 VDD VSS sg13g2_decap_8
XFILLER_10_294 VDD VSS sg13g2_decap_8
XFILLER_6_287 VDD VSS sg13g2_decap_8
XFILLER_40_70 VDD VSS sg13g2_decap_8
XFILLER_69_217 VDD VSS sg13g2_decap_8
XFILLER_41_7 VDD VSS sg13g2_decap_8
XFILLER_93_721 VDD VSS sg13g2_decap_8
XFILLER_38_637 VDD VSS sg13g2_decap_8
XFILLER_92_231 VDD VSS sg13g2_decap_8
XFILLER_65_434 VDD VSS sg13g2_decap_8
XFILLER_1_42 VDD VSS sg13g2_decap_8
XFILLER_37_147 VDD VSS sg13g2_decap_8
XFILLER_18_350 VDD VSS sg13g2_decap_8
XFILLER_80_448 VDD VSS sg13g2_decap_8
XFILLER_61_651 VDD VSS sg13g2_decap_8
XFILLER_33_364 VDD VSS sg13g2_decap_8
XFILLER_21_504 VDD VSS sg13g2_decap_8
XFILLER_60_161 VDD VSS sg13g2_decap_8
XFILLER_88_504 VDD VSS sg13g2_decap_8
Xhold16 _50_/Y VDD VSS _55_/A2 sg13g2_dlygate4sd3_1
Xhold27 _61_/Y VDD VSS _78_/D sg13g2_dlygate4sd3_1
XFILLER_29_49 VDD VSS sg13g2_decap_8
XFILLER_84_721 VDD VSS sg13g2_decap_8
XFILLER_68_272 VDD VSS sg13g2_decap_8
XFILLER_29_637 VDD VSS sg13g2_decap_8
XFILLER_83_231 VDD VSS sg13g2_decap_8
XFILLER_28_147 VDD VSS sg13g2_decap_8
XFILLER_56_434 VDD VSS sg13g2_decap_8
XFILLER_52_651 VDD VSS sg13g2_decap_8
XFILLER_12_504 VDD VSS sg13g2_decap_8
XFILLER_61_14 VDD VSS sg13g2_decap_8
XFILLER_24_364 VDD VSS sg13g2_decap_8
XFILLER_51_161 VDD VSS sg13g2_decap_8
XFILLER_20_581 VDD VSS sg13g2_decap_8
XFILLER_4_714 VDD VSS sg13g2_decap_8
XFILLER_3_224 VDD VSS sg13g2_decap_8
XFILLER_79_504 VDD VSS sg13g2_decap_8
XFILLER_10_84 VDD VSS sg13g2_decap_8
XFILLER_94_518 VDD VSS sg13g2_decap_8
XFILLER_87_581 VDD VSS sg13g2_decap_8
XFILLER_75_732 VDD VSS sg13g2_decap_8
XFILLER_86_77 VDD VSS sg13g2_decap_8
XFILLER_74_231 VDD VSS sg13g2_decap_4
XFILLER_19_147 VDD VSS sg13g2_decap_8
XFILLER_47_434 VDD VSS sg13g2_decap_8
XFILLER_59_294 VDD VSS sg13g2_decap_8
XFILLER_90_735 VDD VSS sg13g2_decap_8
XFILLER_74_297 VDD VSS sg13g2_fill_1
XFILLER_74_286 VDD VSS sg13g2_decap_8
XFILLER_62_448 VDD VSS sg13g2_decap_8
XFILLER_35_70 VDD VSS sg13g2_decap_8
XFILLER_43_651 VDD VSS sg13g2_decap_8
XFILLER_15_364 VDD VSS sg13g2_decap_8
XFILLER_30_301 VDD VSS sg13g2_decap_8
XFILLER_42_161 VDD VSS sg13g2_decap_8
XFILLER_89_7 VDD VSS sg13g2_decap_8
XFILLER_30_378 VDD VSS sg13g2_decap_8
XFILLER_11_581 VDD VSS sg13g2_decap_8
XFILLER_51_91 VDD VSS sg13g2_decap_8
XFILLER_7_574 VDD VSS sg13g2_decap_8
XFILLER_85_518 VDD VSS sg13g2_decap_8
XFILLER_78_581 VDD VSS sg13g2_decap_8
XFILLER_65_231 VDD VSS sg13g2_decap_8
XFILLER_38_434 VDD VSS sg13g2_decap_8
XFILLER_26_629 VDD VSS sg13g2_decap_8
XFILLER_93_595 VDD VSS sg13g2_decap_8
XFILLER_81_735 VDD VSS sg13g2_decap_8
XFILLER_53_448 VDD VSS sg13g2_decap_8
XFILLER_80_245 VDD VSS sg13g2_decap_8
XFILLER_34_651 VDD VSS sg13g2_decap_8
XFILLER_21_301 VDD VSS sg13g2_decap_8
XFILLER_33_161 VDD VSS sg13g2_decap_8
XFILLER_21_378 VDD VSS sg13g2_decap_8
XFILLER_31_28 VDD VSS sg13g2_decap_8
XIO_BOND_outputs\[0\].output_pad output_PAD[0] bondpad_70x70_novias
XFILLER_88_301 VDD VSS sg13g2_decap_8
XFILLER_1_728 VDD VSS sg13g2_decap_8
XFILLER_0_238 VDD VSS sg13g2_decap_8
XFILLER_88_378 VDD VSS sg13g2_decap_8
XFILLER_57_721 VDD VSS sg13g2_decap_8
XFILLER_56_14 VDD VSS sg13g2_decap_8
XFILLER_29_434 VDD VSS sg13g2_decap_8
XFILLER_56_231 VDD VSS sg13g2_decap_8
XFILLER_84_595 VDD VSS sg13g2_decap_8
XFILLER_71_212 VDD VSS sg13g2_fill_1
XFILLER_44_448 VDD VSS sg13g2_decap_8
XFILLER_71_256 VDD VSS sg13g2_decap_8
XFILLER_25_651 VDD VSS sg13g2_decap_8
XFILLER_71_289 VDD VSS sg13g2_fill_1
XFILLER_72_35 VDD VSS sg13g2_decap_8
XFILLER_12_301 VDD VSS sg13g2_decap_8
XFILLER_24_161 VDD VSS sg13g2_decap_8
XFILLER_12_378 VDD VSS sg13g2_decap_8
XFILLER_40_665 VDD VSS sg13g2_decap_8
XFILLER_4_511 VDD VSS sg13g2_decap_8
XFILLER_79_301 VDD VSS sg13g2_decap_8
XFILLER_4_588 VDD VSS sg13g2_decap_8
XFILLER_94_315 VDD VSS sg13g2_decap_8
XFILLER_79_378 VDD VSS sg13g2_decap_8
XFILLER_48_721 VDD VSS sg13g2_decap_8
XFILLER_47_231 VDD VSS sg13g2_decap_8
XFILLER_90_532 VDD VSS sg13g2_decap_8
XFILLER_63_746 VDD VSS sg13g2_decap_8
XFILLER_62_245 VDD VSS sg13g2_decap_8
XFILLER_46_91 VDD VSS sg13g2_decap_8
XFILLER_35_448 VDD VSS sg13g2_decap_8
XFILLER_16_651 VDD VSS sg13g2_decap_8
XFILLER_15_161 VDD VSS sg13g2_decap_8
XFILLER_31_665 VDD VSS sg13g2_decap_8
XFILLER_30_175 VDD VSS sg13g2_decap_8
XFILLER_7_63 VDD VSS sg13g2_decap_8
XFILLER_7_371 VDD VSS sg13g2_decap_8
XFILLER_30_0 VDD VSS sg13g2_decap_8
XFILLER_85_315 VDD VSS sg13g2_decap_8
XFILLER_58_518 VDD VSS sg13g2_decap_8
XFILLER_39_721 VDD VSS sg13g2_decap_8
XFILLER_66_562 VDD VSS sg13g2_decap_8
XFILLER_38_231 VDD VSS sg13g2_decap_8
XFILLER_81_532 VDD VSS sg13g2_decap_8
XFILLER_93_392 VDD VSS sg13g2_decap_8
XFILLER_54_735 VDD VSS sg13g2_decap_8
XFILLER_26_28 VDD VSS sg13g2_decap_8
XFILLER_26_426 VDD VSS sg13g2_decap_8
XFILLER_53_245 VDD VSS sg13g2_decap_8
XFILLER_42_49 VDD VSS sg13g2_decap_8
XFILLER_22_665 VDD VSS sg13g2_decap_8
XFILLER_21_175 VDD VSS sg13g2_decap_8
XFILLER_5_308 VDD VSS sg13g2_decap_8
XFILLER_1_525 VDD VSS sg13g2_decap_8
XFILLER_89_665 VDD VSS sg13g2_decap_8
XFILLER_88_175 VDD VSS sg13g2_decap_8
XFILLER_67_35 VDD VSS sg13g2_decap_8
XFILLER_49_518 VDD VSS sg13g2_decap_8
XFILLER_76_348 VDD VSS sg13g2_decap_8
XFILLER_29_231 VDD VSS sg13g2_decap_8
XFILLER_91_329 VDD VSS sg13g2_decap_8
XFILLER_57_595 VDD VSS sg13g2_decap_8
XFILLER_45_735 VDD VSS sg13g2_decap_8
XFILLER_72_565 VDD VSS sg13g2_decap_8
XFILLER_84_392 VDD VSS sg13g2_decap_8
XFILLER_83_56 VDD VSS sg13g2_decap_8
XFILLER_17_448 VDD VSS sg13g2_decap_8
XFILLER_44_245 VDD VSS sg13g2_decap_8
XFILLER_60_749 VDD VSS sg13g2_decap_8
XFILLER_13_665 VDD VSS sg13g2_decap_8
XFILLER_40_462 VDD VSS sg13g2_decap_8
XFILLER_9_658 VDD VSS sg13g2_decap_8
XFILLER_12_175 VDD VSS sg13g2_decap_8
XFILLER_8_168 VDD VSS sg13g2_decap_8
XFILLER_4_385 VDD VSS sg13g2_decap_8
XFILLER_95_602 VDD VSS sg13g2_decap_8
XFILLER_79_175 VDD VSS sg13g2_decap_8
XFILLER_94_112 VDD VSS sg13g2_decap_8
XFILLER_95_679 VDD VSS sg13g2_decap_8
XFILLER_67_359 VDD VSS sg13g2_decap_8
XFILLER_94_189 VDD VSS sg13g2_decap_8
XFILLER_82_329 VDD VSS sg13g2_decap_8
XFILLER_75_381 VDD VSS sg13g2_decap_8
XFILLER_48_595 VDD VSS sg13g2_decap_8
XFILLER_36_735 VDD VSS sg13g2_decap_8
XFILLER_63_543 VDD VSS sg13g2_decap_8
XFILLER_35_245 VDD VSS sg13g2_decap_8
XFILLER_51_749 VDD VSS sg13g2_decap_8
XFILLER_31_462 VDD VSS sg13g2_decap_8
XFILLER_50_259 VDD VSS sg13g2_decap_8
XFILLER_78_0 VDD VSS sg13g2_decap_8
XFILLER_86_602 VDD VSS sg13g2_decap_8
XFILLER_58_315 VDD VSS sg13g2_decap_8
XFILLER_85_112 VDD VSS sg13g2_decap_8
XFILLER_86_679 VDD VSS sg13g2_decap_8
XFILLER_37_49 VDD VSS sg13g2_decap_8
XFILLER_85_189 VDD VSS sg13g2_decap_8
XFILLER_73_318 VDD VSS sg13g2_decap_8
XFILLER_27_735 VDD VSS sg13g2_decap_8
XFILLER_39_595 VDD VSS sg13g2_decap_8
XFILLER_66_392 VDD VSS sg13g2_decap_8
XFILLER_54_532 VDD VSS sg13g2_decap_8
XFILLER_26_245 VDD VSS sg13g2_decap_8
XFILLER_42_749 VDD VSS sg13g2_decap_8
XFILLER_10_602 VDD VSS sg13g2_decap_8
XFILLER_22_462 VDD VSS sg13g2_decap_8
XFILLER_41_259 VDD VSS sg13g2_decap_8
XFILLER_10_679 VDD VSS sg13g2_decap_8
XFILLER_5_105 VDD VSS sg13g2_decap_8
XFILLER_78_56 VDD VSS sg13g2_decap_8
XFILLER_1_322 VDD VSS sg13g2_decap_8
XFILLER_89_462 VDD VSS sg13g2_decap_8
XFILLER_49_315 VDD VSS sg13g2_decap_8
XFILLER_77_646 VDD VSS sg13g2_decap_8
XFILLER_76_112 VDD VSS sg13g2_decap_8
XFILLER_1_399 VDD VSS sg13g2_decap_8
XFILLER_92_616 VDD VSS sg13g2_decap_8
XFILLER_91_126 VDD VSS sg13g2_decap_8
XFILLER_76_189 VDD VSS sg13g2_decap_8
XFILLER_64_329 VDD VSS sg13g2_decap_8
XFILLER_94_77 VDD VSS sg13g2_decap_8
XFILLER_18_735 VDD VSS sg13g2_decap_8
XFILLER_17_245 VDD VSS sg13g2_decap_8
XFILLER_57_392 VDD VSS sg13g2_decap_8
XFILLER_45_532 VDD VSS sg13g2_decap_8
XFILLER_72_395 VDD VSS sg13g2_decap_8
XFILLER_60_546 VDD VSS sg13g2_decap_8
XFILLER_33_749 VDD VSS sg13g2_decap_8
XFILLER_32_259 VDD VSS sg13g2_decap_8
XFILLER_13_462 VDD VSS sg13g2_decap_8
XFILLER_43_70 VDD VSS sg13g2_decap_8
XFILLER_71_7 VDD VSS sg13g2_decap_8
XFILLER_9_455 VDD VSS sg13g2_decap_8
XFILLER_5_672 VDD VSS sg13g2_decap_8
XFILLER_4_182 VDD VSS sg13g2_decap_8
XFILLER_4_42 VDD VSS sg13g2_decap_8
XFILLER_68_657 VDD VSS sg13g2_decap_8
XFILLER_67_112 VDD VSS sg13g2_decap_8
XFILLER_83_616 VDD VSS sg13g2_decap_8
XFILLER_95_476 VDD VSS sg13g2_decap_8
XFILLER_82_126 VDD VSS sg13g2_decap_8
XFILLER_67_189 VDD VSS sg13g2_decap_8
XFILLER_55_329 VDD VSS sg13g2_decap_8
XFILLER_48_392 VDD VSS sg13g2_decap_8
XFILLER_36_532 VDD VSS sg13g2_decap_8
XFILLER_91_693 VDD VSS sg13g2_decap_8
XFILLER_51_546 VDD VSS sg13g2_decap_8
XFILLER_24_749 VDD VSS sg13g2_decap_8
XFILLER_23_259 VDD VSS sg13g2_decap_8
XFILLER_3_609 VDD VSS sg13g2_decap_8
XFILLER_2_119 VDD VSS sg13g2_decap_8
XFILLER_59_602 VDD VSS sg13g2_decap_8
XFILLER_58_112 VDD VSS sg13g2_decap_8
XFILLER_74_616 VDD VSS sg13g2_decap_8
XFILLER_59_679 VDD VSS sg13g2_decap_8
XFILLER_86_476 VDD VSS sg13g2_decap_8
XFILLER_73_126 VDD VSS sg13g2_decap_8
XFILLER_46_329 VDD VSS sg13g2_decap_8
XFILLER_58_189 VDD VSS sg13g2_decap_8
XFILLER_64_14 VDD VSS sg13g2_decap_8
XFILLER_39_392 VDD VSS sg13g2_decap_8
XFILLER_27_532 VDD VSS sg13g2_decap_8
XFILLER_82_693 VDD VSS sg13g2_decap_8
XFILLER_15_749 VDD VSS sg13g2_decap_8
XFILLER_42_546 VDD VSS sg13g2_decap_8
XFILLER_14_259 VDD VSS sg13g2_decap_8
XFILLER_80_35 VDD VSS sg13g2_decap_8
XFILLER_10_476 VDD VSS sg13g2_decap_8
XFILLER_13_84 VDD VSS sg13g2_decap_8
XFILLER_6_469 VDD VSS sg13g2_decap_8
XFILLER_89_77 VDD VSS sg13g2_decap_8
XFILLER_8_0 VDD VSS sg13g2_decap_8
XFILLER_77_421 VDD VSS sg13g2_decap_8
XFILLER_2_686 VDD VSS sg13g2_decap_8
XFILLER_49_112 VDD VSS sg13g2_decap_8
XFILLER_65_605 VDD VSS sg13g2_decap_8
XFILLER_1_196 VDD VSS sg13g2_decap_8
XFILLER_92_413 VDD VSS sg13g2_decap_8
XFILLER_38_70 VDD VSS sg13g2_decap_8
XFILLER_37_329 VDD VSS sg13g2_decap_8
XFILLER_49_189 VDD VSS sg13g2_decap_8
XFILLER_64_126 VDD VSS sg13g2_decap_8
XFILLER_18_532 VDD VSS sg13g2_decap_8
XFILLER_73_660 VDD VSS sg13g2_decap_8
XFILLER_33_546 VDD VSS sg13g2_decap_8
XFILLER_54_91 VDD VSS sg13g2_decap_8
XFILLER_60_343 VDD VSS sg13g2_decap_8
XFILLER_9_252 VDD VSS sg13g2_decap_8
XIO_BOND_outputs\[5\].output_pad output_PAD[5] bondpad_70x70_novias
XFILLER_68_454 VDD VSS sg13g2_decap_8
XFILLER_95_273 VDD VSS sg13g2_decap_8
XFILLER_83_413 VDD VSS sg13g2_decap_8
XFILLER_56_616 VDD VSS sg13g2_decap_8
XFILLER_28_329 VDD VSS sg13g2_decap_8
XFILLER_55_126 VDD VSS sg13g2_decap_8
XFILLER_91_490 VDD VSS sg13g2_decap_8
XFILLER_64_693 VDD VSS sg13g2_decap_8
XFILLER_34_28 VDD VSS sg13g2_decap_8
XFILLER_24_546 VDD VSS sg13g2_decap_8
XFILLER_51_343 VDD VSS sg13g2_decap_8
XFILLER_50_49 VDD VSS sg13g2_decap_8
XFILLER_3_406 VDD VSS sg13g2_decap_8
XFILLER_59_14 VDD VSS sg13g2_decap_8
XFILLER_1_7 VDD VSS sg13g2_decap_8
XFILLER_86_273 VDD VSS sg13g2_decap_8
XFILLER_74_402 VDD VSS sg13g2_decap_8
XFILLER_75_46 VDD VSS sg13g2_decap_8
XFILLER_47_616 VDD VSS sg13g2_decap_8
XFILLER_19_329 VDD VSS sg13g2_decap_8
XFILLER_59_476 VDD VSS sg13g2_decap_8
XFILLER_46_126 VDD VSS sg13g2_decap_8
XFILLER_82_490 VDD VSS sg13g2_decap_8
XFILLER_55_693 VDD VSS sg13g2_decap_8
XFILLER_70_652 VDD VSS sg13g2_decap_8
XFILLER_91_56 VDD VSS sg13g2_decap_8
XFILLER_42_343 VDD VSS sg13g2_decap_8
XFILLER_15_546 VDD VSS sg13g2_decap_8
XFILLER_7_756 VDD VSS sg13g2_fill_1
XFILLER_10_273 VDD VSS sg13g2_decap_8
XFILLER_6_266 VDD VSS sg13g2_decap_8
XFILLER_2_483 VDD VSS sg13g2_decap_8
XFILLER_34_7 VDD VSS sg13g2_decap_8
XFILLER_49_91 VDD VSS sg13g2_decap_8
XFILLER_93_700 VDD VSS sg13g2_decap_8
XFILLER_65_413 VDD VSS sg13g2_decap_8
XFILLER_1_21 VDD VSS sg13g2_decap_8
XFILLER_38_616 VDD VSS sg13g2_decap_8
XFILLER_92_210 VDD VSS sg13g2_decap_8
XFILLER_77_295 VDD VSS sg13g2_decap_8
XFILLER_37_126 VDD VSS sg13g2_decap_8
XFILLER_1_98 VDD VSS sg13g2_decap_8
XFILLER_92_287 VDD VSS sg13g2_decap_8
XFILLER_80_427 VDD VSS sg13g2_decap_8
XFILLER_61_630 VDD VSS sg13g2_decap_8
XFILLER_46_693 VDD VSS sg13g2_decap_8
XFILLER_33_343 VDD VSS sg13g2_decap_8
XFILLER_60_140 VDD VSS sg13g2_decap_8
XFILLER_60_0 VDD VSS sg13g2_decap_8
XFILLER_69_741 VDD VSS sg13g2_decap_8
Xhold17 _54_/Y VDD VSS _76_/D sg13g2_dlygate4sd3_1
Xhold28 _49_/D VDD VSS _52_/B sg13g2_dlygate4sd3_1
XFILLER_29_28 VDD VSS sg13g2_decap_8
XFILLER_84_700 VDD VSS sg13g2_decap_8
XFILLER_68_251 VDD VSS sg13g2_decap_8
XFILLER_56_413 VDD VSS sg13g2_decap_8
XFILLER_29_616 VDD VSS sg13g2_decap_8
XFILLER_83_210 VDD VSS sg13g2_decap_8
XFILLER_28_126 VDD VSS sg13g2_decap_8
XFILLER_83_287 VDD VSS sg13g2_decap_8
XFILLER_45_49 VDD VSS sg13g2_decap_8
XFILLER_37_693 VDD VSS sg13g2_decap_8
XFILLER_64_490 VDD VSS sg13g2_decap_8
XFILLER_52_630 VDD VSS sg13g2_decap_8
XFILLER_24_343 VDD VSS sg13g2_decap_8
XFILLER_51_140 VDD VSS sg13g2_decap_8
XFILLER_20_560 VDD VSS sg13g2_decap_8
XFILLER_3_203 VDD VSS sg13g2_decap_8
XFILLER_10_63 VDD VSS sg13g2_decap_8
XFILLER_86_56 VDD VSS sg13g2_decap_8
XFILLER_87_560 VDD VSS sg13g2_decap_8
XFILLER_75_711 VDD VSS sg13g2_decap_8
XFILLER_47_413 VDD VSS sg13g2_decap_8
XFILLER_59_273 VDD VSS sg13g2_decap_8
XFILLER_74_210 VDD VSS sg13g2_decap_8
XFILLER_19_126 VDD VSS sg13g2_decap_8
XFILLER_90_714 VDD VSS sg13g2_decap_8
XFILLER_62_427 VDD VSS sg13g2_decap_8
XFILLER_28_693 VDD VSS sg13g2_decap_8
XFILLER_55_490 VDD VSS sg13g2_decap_8
XFILLER_15_343 VDD VSS sg13g2_decap_8
XFILLER_43_630 VDD VSS sg13g2_decap_8
XFILLER_42_140 VDD VSS sg13g2_decap_8
XFILLER_11_560 VDD VSS sg13g2_decap_8
XFILLER_30_357 VDD VSS sg13g2_decap_8
XFILLER_51_70 VDD VSS sg13g2_decap_8
XFILLER_7_553 VDD VSS sg13g2_decap_8
XFILLER_2_280 VDD VSS sg13g2_decap_8
XFILLER_78_560 VDD VSS sg13g2_decap_8
XFILLER_38_413 VDD VSS sg13g2_decap_8
XFILLER_66_755 VDD VSS sg13g2_fill_2
XFILLER_66_744 VDD VSS sg13g2_decap_8
XFILLER_65_210 VDD VSS sg13g2_decap_8
XFILLER_93_574 VDD VSS sg13g2_decap_8
XFILLER_81_714 VDD VSS sg13g2_decap_8
XFILLER_26_608 VDD VSS sg13g2_decap_8
XFILLER_80_224 VDD VSS sg13g2_decap_8
XFILLER_65_287 VDD VSS sg13g2_decap_8
XFILLER_53_427 VDD VSS sg13g2_decap_8
XFILLER_19_693 VDD VSS sg13g2_decap_8
XFILLER_46_490 VDD VSS sg13g2_decap_8
XFILLER_34_630 VDD VSS sg13g2_decap_8
XFILLER_33_140 VDD VSS sg13g2_decap_8
XFILLER_21_357 VDD VSS sg13g2_decap_8
XFILLER_1_707 VDD VSS sg13g2_decap_8
XFILLER_0_217 VDD VSS sg13g2_decap_8
XFILLER_88_357 VDD VSS sg13g2_decap_8
XFILLER_57_700 VDD VSS sg13g2_decap_8
XFILLER_29_413 VDD VSS sg13g2_decap_8
XFILLER_56_210 VDD VSS sg13g2_decap_8
XFILLER_84_574 VDD VSS sg13g2_decap_8
XFILLER_72_747 VDD VSS sg13g2_decap_8
XFILLER_44_427 VDD VSS sg13g2_decap_8
XFILLER_56_287 VDD VSS sg13g2_decap_8
XFILLER_71_235 VDD VSS sg13g2_decap_8
XFILLER_72_14 VDD VSS sg13g2_decap_8
XFILLER_25_630 VDD VSS sg13g2_decap_8
XFILLER_37_490 VDD VSS sg13g2_decap_8
XFILLER_24_140 VDD VSS sg13g2_decap_8
XFILLER_40_644 VDD VSS sg13g2_decap_8
XFILLER_12_357 VDD VSS sg13g2_decap_8
XFILLER_4_567 VDD VSS sg13g2_decap_8
XFILLER_21_84 VDD VSS sg13g2_decap_8
XFILLER_79_357 VDD VSS sg13g2_decap_8
XFILLER_48_700 VDD VSS sg13g2_decap_8
XFILLER_47_210 VDD VSS sg13g2_decap_8
XFILLER_90_511 VDD VSS sg13g2_decap_8
XFILLER_75_585 VDD VSS sg13g2_decap_8
XFILLER_63_725 VDD VSS sg13g2_decap_8
XFILLER_62_224 VDD VSS sg13g2_decap_8
XFILLER_46_70 VDD VSS sg13g2_decap_8
XFILLER_35_427 VDD VSS sg13g2_decap_8
XFILLER_47_287 VDD VSS sg13g2_decap_8
XFILLER_16_630 VDD VSS sg13g2_decap_8
XFILLER_28_490 VDD VSS sg13g2_decap_8
XFILLER_90_588 VDD VSS sg13g2_decap_8
XFILLER_15_140 VDD VSS sg13g2_decap_8
XFILLER_31_644 VDD VSS sg13g2_decap_8
XFILLER_62_91 VDD VSS sg13g2_decap_8
XFILLER_30_154 VDD VSS sg13g2_decap_8
XFILLER_7_350 VDD VSS sg13g2_decap_8
XFILLER_7_42 VDD VSS sg13g2_decap_8
XFILLER_23_0 VDD VSS sg13g2_decap_8
XFILLER_39_700 VDD VSS sg13g2_decap_8
XFILLER_38_210 VDD VSS sg13g2_decap_8
XFILLER_66_541 VDD VSS sg13g2_decap_8
XFILLER_81_511 VDD VSS sg13g2_decap_8
XFILLER_93_371 VDD VSS sg13g2_decap_8
XFILLER_54_714 VDD VSS sg13g2_decap_8
XFILLER_26_405 VDD VSS sg13g2_decap_8
XFILLER_38_287 VDD VSS sg13g2_decap_8
XFILLER_53_224 VDD VSS sg13g2_decap_8
XFILLER_19_490 VDD VSS sg13g2_decap_8
XFILLER_81_588 VDD VSS sg13g2_decap_8
XFILLER_22_644 VDD VSS sg13g2_decap_8
XFILLER_42_28 VDD VSS sg13g2_decap_8
XFILLER_21_154 VDD VSS sg13g2_decap_8
XFILLER_1_504 VDD VSS sg13g2_decap_8
XIO_CORNER_SOUTH_EAST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XFILLER_89_644 VDD VSS sg13g2_decap_8
XFILLER_67_14 VDD VSS sg13g2_decap_8
XFILLER_88_154 VDD VSS sg13g2_decap_8
XFILLER_76_327 VDD VSS sg13g2_decap_8
XFILLER_29_210 VDD VSS sg13g2_decap_8
XFILLER_91_308 VDD VSS sg13g2_decap_8
XFILLER_84_371 VDD VSS sg13g2_decap_8
XFILLER_83_35 VDD VSS sg13g2_decap_8
XFILLER_57_574 VDD VSS sg13g2_decap_8
XFILLER_17_427 VDD VSS sg13g2_decap_8
XFILLER_29_287 VDD VSS sg13g2_decap_8
XFILLER_45_714 VDD VSS sg13g2_decap_8
XFILLER_72_544 VDD VSS sg13g2_decap_8
XFILLER_44_224 VDD VSS sg13g2_decap_8
XFILLER_60_728 VDD VSS sg13g2_decap_8
XFILLER_13_644 VDD VSS sg13g2_decap_8
XFILLER_16_84 VDD VSS sg13g2_decap_8
XFILLER_12_154 VDD VSS sg13g2_decap_8
XFILLER_40_441 VDD VSS sg13g2_decap_8
XFILLER_9_637 VDD VSS sg13g2_decap_8
XFILLER_8_147 VDD VSS sg13g2_decap_8
XFILLER_4_364 VDD VSS sg13g2_decap_8
XFILLER_79_154 VDD VSS sg13g2_decap_8
XFILLER_95_658 VDD VSS sg13g2_decap_8
XFILLER_67_338 VDD VSS sg13g2_decap_8
XFILLER_0_581 VDD VSS sg13g2_decap_8
XFILLER_94_168 VDD VSS sg13g2_decap_8
XFILLER_82_308 VDD VSS sg13g2_decap_8
XFILLER_63_522 VDD VSS sg13g2_decap_8
XFILLER_75_360 VDD VSS sg13g2_decap_8
XFILLER_48_574 VDD VSS sg13g2_decap_8
XFILLER_57_91 VDD VSS sg13g2_decap_8
XFILLER_36_714 VDD VSS sg13g2_decap_8
XFILLER_35_224 VDD VSS sg13g2_decap_8
XFILLER_51_728 VDD VSS sg13g2_decap_8
XFILLER_63_599 VDD VSS sg13g2_decap_8
XFILLER_90_385 VDD VSS sg13g2_decap_8
XFILLER_50_238 VDD VSS sg13g2_decap_8
XFILLER_31_441 VDD VSS sg13g2_decap_8
XFILLER_86_658 VDD VSS sg13g2_decap_8
XFILLER_85_168 VDD VSS sg13g2_decap_8
XFILLER_37_28 VDD VSS sg13g2_decap_8
XFILLER_66_371 VDD VSS sg13g2_decap_8
XFILLER_54_511 VDD VSS sg13g2_decap_8
XFILLER_27_714 VDD VSS sg13g2_decap_8
XFILLER_39_574 VDD VSS sg13g2_decap_8
XFILLER_26_224 VDD VSS sg13g2_decap_8
XFILLER_54_588 VDD VSS sg13g2_decap_8
XFILLER_42_728 VDD VSS sg13g2_decap_8
XFILLER_81_385 VDD VSS sg13g2_decap_8
XFILLER_53_49 VDD VSS sg13g2_decap_8
XFILLER_41_238 VDD VSS sg13g2_decap_8
XFILLER_22_441 VDD VSS sg13g2_decap_8
XFILLER_10_658 VDD VSS sg13g2_decap_8
XFILLER_1_301 VDD VSS sg13g2_decap_8
XFILLER_89_441 VDD VSS sg13g2_decap_8
XFILLER_78_35 VDD VSS sg13g2_decap_8
XFILLER_77_625 VDD VSS sg13g2_decap_8
XFILLER_1_378 VDD VSS sg13g2_decap_8
XFILLER_64_308 VDD VSS sg13g2_decap_8
XFILLER_76_168 VDD VSS sg13g2_decap_8
XFILLER_94_56 VDD VSS sg13g2_decap_8
XFILLER_91_105 VDD VSS sg13g2_decap_8
XFILLER_57_371 VDD VSS sg13g2_decap_8
XFILLER_18_714 VDD VSS sg13g2_decap_8
XFILLER_45_511 VDD VSS sg13g2_decap_8
XFILLER_17_224 VDD VSS sg13g2_decap_8
XFILLER_72_374 VDD VSS sg13g2_decap_8
XFILLER_33_728 VDD VSS sg13g2_decap_8
XFILLER_45_588 VDD VSS sg13g2_decap_8
XFILLER_60_525 VDD VSS sg13g2_decap_8
XFILLER_32_238 VDD VSS sg13g2_decap_8
XFILLER_13_441 VDD VSS sg13g2_decap_8
XFILLER_9_434 VDD VSS sg13g2_decap_8
XFILLER_64_7 VDD VSS sg13g2_decap_8
XFILLER_5_651 VDD VSS sg13g2_decap_8
XFILLER_4_161 VDD VSS sg13g2_decap_8
XFILLER_4_21 VDD VSS sg13g2_decap_8
XFILLER_68_636 VDD VSS sg13g2_decap_8
XFILLER_4_98 VDD VSS sg13g2_decap_8
XFILLER_95_455 VDD VSS sg13g2_decap_8
XFILLER_67_168 VDD VSS sg13g2_decap_8
XFILLER_82_105 VDD VSS sg13g2_decap_8
XFILLER_48_371 VDD VSS sg13g2_decap_8
XFILLER_55_308 VDD VSS sg13g2_decap_8
XFILLER_36_511 VDD VSS sg13g2_decap_8
XFILLER_91_672 VDD VSS sg13g2_decap_8
XFILLER_24_728 VDD VSS sg13g2_decap_8
XFILLER_36_588 VDD VSS sg13g2_decap_8
XFILLER_90_182 VDD VSS sg13g2_decap_8
XFILLER_63_385 VDD VSS sg13g2_decap_8
XFILLER_51_525 VDD VSS sg13g2_decap_8
XFILLER_23_238 VDD VSS sg13g2_decap_8
XFILLER_90_0 VDD VSS sg13g2_decap_8
XFILLER_48_49 VDD VSS sg13g2_decap_8
XFILLER_86_455 VDD VSS sg13g2_decap_8
XFILLER_59_658 VDD VSS sg13g2_decap_8
XFILLER_73_105 VDD VSS sg13g2_decap_8
XFILLER_39_371 VDD VSS sg13g2_decap_8
XFILLER_46_308 VDD VSS sg13g2_decap_8
XFILLER_58_168 VDD VSS sg13g2_decap_8
XFILLER_27_511 VDD VSS sg13g2_decap_8
XFILLER_82_672 VDD VSS sg13g2_decap_8
XFILLER_15_728 VDD VSS sg13g2_decap_8
XFILLER_81_182 VDD VSS sg13g2_decap_8
XFILLER_14_238 VDD VSS sg13g2_decap_8
XFILLER_54_385 VDD VSS sg13g2_decap_8
XFILLER_27_588 VDD VSS sg13g2_decap_8
XFILLER_42_525 VDD VSS sg13g2_decap_8
XFILLER_80_14 VDD VSS sg13g2_decap_8
XFILLER_10_455 VDD VSS sg13g2_decap_8
XFILLER_13_63 VDD VSS sg13g2_decap_8
XFILLER_6_448 VDD VSS sg13g2_decap_8
XFILLER_89_56 VDD VSS sg13g2_decap_8
XFILLER_2_665 VDD VSS sg13g2_decap_8
XFILLER_1_175 VDD VSS sg13g2_decap_8
XFILLER_77_499 VDD VSS sg13g2_decap_8
XFILLER_64_105 VDD VSS sg13g2_decap_8
XFILLER_37_308 VDD VSS sg13g2_decap_8
XFILLER_49_168 VDD VSS sg13g2_decap_8
XFILLER_18_511 VDD VSS sg13g2_decap_8
XFILLER_80_609 VDD VSS sg13g2_decap_8
XFILLER_92_469 VDD VSS sg13g2_decap_8
XFILLER_72_182 VDD VSS sg13g2_decap_8
XFILLER_45_385 VDD VSS sg13g2_decap_8
XFILLER_60_322 VDD VSS sg13g2_decap_8
XFILLER_18_588 VDD VSS sg13g2_decap_8
XFILLER_33_525 VDD VSS sg13g2_decap_8
XFILLER_54_70 VDD VSS sg13g2_decap_8
XFILLER_60_399 VDD VSS sg13g2_decap_8
XFILLER_9_231 VDD VSS sg13g2_decap_8
XFILLER_70_91 VDD VSS sg13g2_decap_8
XFILLER_68_433 VDD VSS sg13g2_decap_8
XFILLER_95_252 VDD VSS sg13g2_decap_8
XFILLER_55_105 VDD VSS sg13g2_decap_8
XFILLER_28_308 VDD VSS sg13g2_decap_8
XFILLER_64_672 VDD VSS sg13g2_decap_8
XFILLER_83_469 VDD VSS sg13g2_decap_8
XFILLER_70_119 VDD VSS sg13g2_decap_8
XFILLER_63_182 VDD VSS sg13g2_decap_8
XFILLER_36_385 VDD VSS sg13g2_decap_8
XFILLER_51_322 VDD VSS sg13g2_decap_8
XFILLER_24_525 VDD VSS sg13g2_decap_8
XFILLER_51_399 VDD VSS sg13g2_decap_8
XFILLER_20_742 VDD VSS sg13g2_decap_8
XFILLER_50_28 VDD VSS sg13g2_decap_8
XFILLER_87_742 VDD VSS sg13g2_decap_8
XFILLER_59_455 VDD VSS sg13g2_decap_8
XFILLER_86_252 VDD VSS sg13g2_decap_8
XFILLER_75_14 VDD VSS sg13g2_decap_8
XFILLER_46_105 VDD VSS sg13g2_decap_8
XFILLER_19_308 VDD VSS sg13g2_decap_8
XFILLER_62_609 VDD VSS sg13g2_decap_8
XFILLER_74_469 VDD VSS sg13g2_decap_8
XFILLER_55_672 VDD VSS sg13g2_decap_8
XFILLER_27_385 VDD VSS sg13g2_decap_8
XFILLER_61_119 VDD VSS sg13g2_decap_8
XFILLER_15_525 VDD VSS sg13g2_decap_8
XFILLER_70_631 VDD VSS sg13g2_decap_8
XFILLER_91_35 VDD VSS sg13g2_decap_8
XFILLER_42_322 VDD VSS sg13g2_decap_8
XFILLER_54_182 VDD VSS sg13g2_decap_8
XFILLER_11_742 VDD VSS sg13g2_decap_8
XFILLER_24_84 VDD VSS sg13g2_decap_8
XFILLER_42_399 VDD VSS sg13g2_decap_8
XFILLER_30_539 VDD VSS sg13g2_decap_8
XFILLER_10_252 VDD VSS sg13g2_decap_8
XFILLER_7_735 VDD VSS sg13g2_decap_8
XFILLER_6_245 VDD VSS sg13g2_decap_8
XFILLER_2_462 VDD VSS sg13g2_decap_8
XFILLER_78_742 VDD VSS sg13g2_decap_8
XFILLER_27_7 VDD VSS sg13g2_decap_8
XFILLER_49_70 VDD VSS sg13g2_decap_8
XFILLER_77_274 VDD VSS sg13g2_decap_8
XFILLER_37_105 VDD VSS sg13g2_decap_8
XFILLER_93_756 VDD VSS sg13g2_fill_1
XFILLER_92_266 VDD VSS sg13g2_decap_8
XFILLER_80_406 VDD VSS sg13g2_decap_8
XFILLER_65_469 VDD VSS sg13g2_fill_2
XFILLER_53_609 VDD VSS sg13g2_decap_8
XFILLER_1_77 VDD VSS sg13g2_decap_8
XFILLER_65_91 VDD VSS sg13g2_decap_8
XFILLER_46_672 VDD VSS sg13g2_decap_8
XFILLER_18_385 VDD VSS sg13g2_decap_8
XFILLER_52_119 VDD VSS sg13g2_decap_8
XFILLER_33_322 VDD VSS sg13g2_decap_8
XFILLER_45_182 VDD VSS sg13g2_decap_8
XFILLER_61_686 VDD VSS sg13g2_decap_8
XFILLER_33_399 VDD VSS sg13g2_decap_8
XFILLER_60_196 VDD VSS sg13g2_decap_8
XFILLER_21_539 VDD VSS sg13g2_decap_8
XFILLER_53_0 VDD VSS sg13g2_decap_8
XFILLER_88_539 VDD VSS sg13g2_decap_8
XFILLER_69_720 VDD VSS sg13g2_decap_8
Xhold18 _79_/Q VDD VSS _66_/B sg13g2_dlygate4sd3_1
Xhold29 _52_/Y VDD VSS _57_/B sg13g2_dlygate4sd3_1
XFILLER_68_230 VDD VSS sg13g2_decap_8
XFILLER_28_105 VDD VSS sg13g2_decap_8
XFILLER_84_756 VDD VSS sg13g2_fill_1
XFILLER_83_266 VDD VSS sg13g2_decap_8
XFILLER_45_28 VDD VSS sg13g2_decap_8
XFILLER_56_469 VDD VSS sg13g2_decap_8
XFILLER_44_609 VDD VSS sg13g2_decap_8
XFILLER_43_119 VDD VSS sg13g2_decap_8
XFILLER_37_672 VDD VSS sg13g2_decap_8
XFILLER_24_322 VDD VSS sg13g2_decap_8
XFILLER_36_182 VDD VSS sg13g2_decap_8
XFILLER_52_686 VDD VSS sg13g2_decap_8
XFILLER_12_539 VDD VSS sg13g2_decap_8
XFILLER_61_49 VDD VSS sg13g2_decap_8
XFILLER_24_399 VDD VSS sg13g2_decap_8
XFILLER_51_196 VDD VSS sg13g2_decap_8
XFILLER_4_749 VDD VSS sg13g2_decap_8
XFILLER_3_259 VDD VSS sg13g2_decap_8
XFILLER_10_42 VDD VSS sg13g2_decap_8
XFILLER_79_539 VDD VSS sg13g2_decap_8
XFILLER_86_35 VDD VSS sg13g2_decap_8
XFILLER_19_105 VDD VSS sg13g2_decap_8
XFILLER_59_252 VDD VSS sg13g2_decap_8
XFILLER_62_406 VDD VSS sg13g2_decap_8
XFILLER_19_84 VDD VSS sg13g2_decap_8
XFILLER_47_469 VDD VSS sg13g2_decap_8
XFILLER_35_609 VDD VSS sg13g2_decap_8
XFILLER_34_119 VDD VSS sg13g2_decap_8
XFILLER_28_672 VDD VSS sg13g2_decap_8
XFILLER_15_322 VDD VSS sg13g2_decap_8
XFILLER_27_182 VDD VSS sg13g2_decap_8
XFILLER_43_686 VDD VSS sg13g2_decap_8
XFILLER_15_399 VDD VSS sg13g2_decap_8
XFILLER_30_336 VDD VSS sg13g2_decap_8
XFILLER_42_196 VDD VSS sg13g2_decap_8
XFILLER_7_532 VDD VSS sg13g2_decap_8
XFILLER_66_723 VDD VSS sg13g2_decap_8
XFILLER_93_553 VDD VSS sg13g2_decap_8
XFILLER_65_266 VDD VSS sg13g2_decap_8
XFILLER_38_469 VDD VSS sg13g2_decap_8
XFILLER_53_406 VDD VSS sg13g2_decap_8
XFILLER_80_203 VDD VSS sg13g2_decap_8
XFILLER_25_119 VDD VSS sg13g2_decap_8
XFILLER_19_672 VDD VSS sg13g2_decap_8
XFILLER_18_182 VDD VSS sg13g2_decap_8
XFILLER_34_686 VDD VSS sg13g2_decap_8
XFILLER_61_483 VDD VSS sg13g2_decap_8
XFILLER_21_336 VDD VSS sg13g2_decap_8
XFILLER_33_196 VDD VSS sg13g2_decap_8
XFILLER_88_336 VDD VSS sg13g2_decap_8
XFILLER_69_594 VDD VSS sg13g2_decap_8
XFILLER_84_553 VDD VSS sg13g2_decap_8
XFILLER_57_756 VDD VSS sg13g2_fill_1
XFILLER_56_49 VDD VSS sg13g2_decap_8
XFILLER_29_469 VDD VSS sg13g2_decap_8
XFILLER_17_609 VDD VSS sg13g2_decap_8
XIO_CORNER_NORTH_WEST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XFILLER_72_726 VDD VSS sg13g2_decap_8
XFILLER_71_203 VDD VSS sg13g2_decap_8
XFILLER_16_119 VDD VSS sg13g2_decap_8
XFILLER_44_406 VDD VSS sg13g2_decap_8
XFILLER_56_266 VDD VSS sg13g2_decap_8
XFILLER_25_686 VDD VSS sg13g2_decap_8
XFILLER_52_483 VDD VSS sg13g2_decap_8
XFILLER_12_336 VDD VSS sg13g2_decap_8
XFILLER_24_196 VDD VSS sg13g2_decap_8
XFILLER_40_623 VDD VSS sg13g2_decap_8
X_77__10 VDD VSS _77__10/L_HI sg13g2_tiehi
XFILLER_8_329 VDD VSS sg13g2_decap_8
XFILLER_21_63 VDD VSS sg13g2_decap_8
XFILLER_4_546 VDD VSS sg13g2_decap_8
XFILLER_79_336 VDD VSS sg13g2_decap_8
XFILLER_75_564 VDD VSS sg13g2_decap_8
XFILLER_63_704 VDD VSS sg13g2_decap_8
XFILLER_48_756 VDD VSS sg13g2_fill_1
XFILLER_62_203 VDD VSS sg13g2_decap_8
XFILLER_35_406 VDD VSS sg13g2_decap_8
XFILLER_47_266 VDD VSS sg13g2_decap_8
XFILLER_90_567 VDD VSS sg13g2_decap_8
XFILLER_16_686 VDD VSS sg13g2_decap_8
XFILLER_94_7 VDD VSS sg13g2_decap_8
XFILLER_15_196 VDD VSS sg13g2_decap_8
XFILLER_31_623 VDD VSS sg13g2_decap_8
XFILLER_43_483 VDD VSS sg13g2_decap_8
XFILLER_70_291 VDD VSS sg13g2_decap_4
XFILLER_62_70 VDD VSS sg13g2_decap_8
XFILLER_30_133 VDD VSS sg13g2_decap_8
XFILLER_7_21 VDD VSS sg13g2_decap_8
XFILLER_7_98 VDD VSS sg13g2_decap_8
XFILLER_66_520 VDD VSS sg13g2_decap_8
XFILLER_16_0 VDD VSS sg13g2_decap_8
XFILLER_39_756 VDD VSS sg13g2_fill_1
XFILLER_66_597 VDD VSS sg13g2_decap_8
XFILLER_93_350 VDD VSS sg13g2_decap_8
XFILLER_38_266 VDD VSS sg13g2_decap_8
XFILLER_53_203 VDD VSS sg13g2_decap_8
XFILLER_81_567 VDD VSS sg13g2_decap_8
XFILLER_61_280 VDD VSS sg13g2_decap_8
XFILLER_22_623 VDD VSS sg13g2_decap_8
XFILLER_34_483 VDD VSS sg13g2_decap_8
XFILLER_21_133 VDD VSS sg13g2_decap_8
XFILLER_89_623 VDD VSS sg13g2_decap_8
XFILLER_88_133 VDD VSS sg13g2_decap_8
XFILLER_76_306 VDD VSS sg13g2_decap_8
XFILLER_69_380 VDD VSS sg13g2_decap_8
XFILLER_57_553 VDD VSS sg13g2_decap_8
XFILLER_72_523 VDD VSS sg13g2_decap_8
XFILLER_84_350 VDD VSS sg13g2_decap_8
XFILLER_83_14 VDD VSS sg13g2_decap_8
XFILLER_17_406 VDD VSS sg13g2_decap_8
XFILLER_29_266 VDD VSS sg13g2_decap_8
XFILLER_44_203 VDD VSS sg13g2_decap_8
XFILLER_60_707 VDD VSS sg13g2_decap_8
XFILLER_13_623 VDD VSS sg13g2_decap_8
XFILLER_16_63 VDD VSS sg13g2_decap_8
XFILLER_40_420 VDD VSS sg13g2_decap_8
XFILLER_52_280 VDD VSS sg13g2_decap_8
XFILLER_25_483 VDD VSS sg13g2_decap_8
XFILLER_9_616 VDD VSS sg13g2_decap_8
XFILLER_12_133 VDD VSS sg13g2_decap_8
XFILLER_8_126 VDD VSS sg13g2_decap_8
XFILLER_40_497 VDD VSS sg13g2_decap_8
XFILLER_32_84 VDD VSS sg13g2_decap_8
XFILLER_4_343 VDD VSS sg13g2_decap_8
XFILLER_79_133 VDD VSS sg13g2_decap_8
XFILLER_95_637 VDD VSS sg13g2_decap_8
XFILLER_67_317 VDD VSS sg13g2_decap_8
XFILLER_0_560 VDD VSS sg13g2_decap_8
XFILLER_94_147 VDD VSS sg13g2_decap_8
XFILLER_48_553 VDD VSS sg13g2_decap_8
XFILLER_57_70 VDD VSS sg13g2_decap_8
XFILLER_63_501 VDD VSS sg13g2_decap_8
XFILLER_35_203 VDD VSS sg13g2_decap_8
XFILLER_63_578 VDD VSS sg13g2_decap_8
XFILLER_90_364 VDD VSS sg13g2_decap_8
XFILLER_51_707 VDD VSS sg13g2_decap_8
XFILLER_73_91 VDD VSS sg13g2_decap_8
XFILLER_31_420 VDD VSS sg13g2_decap_8
XFILLER_50_217 VDD VSS sg13g2_decap_8
XFILLER_16_483 VDD VSS sg13g2_decap_8
XFILLER_43_280 VDD VSS sg13g2_decap_8
XFILLER_31_497 VDD VSS sg13g2_decap_8
XFILLER_8_693 VDD VSS sg13g2_decap_8
XFILLER_86_637 VDD VSS sg13g2_decap_8
XFILLER_85_147 VDD VSS sg13g2_decap_8
XFILLER_39_553 VDD VSS sg13g2_decap_8
XFILLER_66_350 VDD VSS sg13g2_decap_8
XFILLER_26_203 VDD VSS sg13g2_decap_8
XFILLER_81_364 VDD VSS sg13g2_decap_8
XFILLER_54_567 VDD VSS sg13g2_decap_8
XFILLER_42_707 VDD VSS sg13g2_decap_8
XFILLER_53_28 VDD VSS sg13g2_decap_8
XFILLER_41_217 VDD VSS sg13g2_decap_8
XFILLER_22_420 VDD VSS sg13g2_decap_8
XFILLER_34_280 VDD VSS sg13g2_decap_8
XFILLER_10_637 VDD VSS sg13g2_decap_8
XFILLER_22_497 VDD VSS sg13g2_decap_8
XFILLER_78_14 VDD VSS sg13g2_decap_8
XFILLER_89_420 VDD VSS sg13g2_decap_8
XFILLER_77_604 VDD VSS sg13g2_decap_8
XFILLER_1_357 VDD VSS sg13g2_decap_8
XFILLER_89_497 VDD VSS sg13g2_decap_8
XFILLER_76_147 VDD VSS sg13g2_decap_8
XFILLER_94_35 VDD VSS sg13g2_decap_8
XFILLER_17_203 VDD VSS sg13g2_decap_8
XFILLER_57_350 VDD VSS sg13g2_decap_8
XFILLER_60_504 VDD VSS sg13g2_decap_8
XFILLER_27_84 VDD VSS sg13g2_decap_8
XFILLER_33_707 VDD VSS sg13g2_decap_8
XFILLER_45_567 VDD VSS sg13g2_decap_8
XFILLER_32_217 VDD VSS sg13g2_decap_8
XFILLER_13_420 VDD VSS sg13g2_decap_8
XFILLER_25_280 VDD VSS sg13g2_decap_8
XFILLER_9_413 VDD VSS sg13g2_decap_8
XFILLER_13_497 VDD VSS sg13g2_decap_8
XFILLER_40_294 VDD VSS sg13g2_decap_8
XFILLER_5_630 VDD VSS sg13g2_decap_8
Xvss_pads\[0\].vss_pad IOVDD IOVSS VDD VSS sg13g2_IOPadVss
XFILLER_4_140 VDD VSS sg13g2_decap_8
XFILLER_57_7 VDD VSS sg13g2_decap_8
XFILLER_4_77 VDD VSS sg13g2_decap_8
XFILLER_68_615 VDD VSS sg13g2_decap_8
XFILLER_95_434 VDD VSS sg13g2_decap_8
XFILLER_67_147 VDD VSS sg13g2_decap_8
XFILLER_68_91 VDD VSS sg13g2_decap_8
XFILLER_48_350 VDD VSS sg13g2_decap_8
XFILLER_76_692 VDD VSS sg13g2_decap_8
XFILLER_91_651 VDD VSS sg13g2_decap_8
XFILLER_63_364 VDD VSS sg13g2_decap_8
XFILLER_51_504 VDD VSS sg13g2_decap_8
XFILLER_24_707 VDD VSS sg13g2_decap_8
XFILLER_36_567 VDD VSS sg13g2_decap_8
XFILLER_90_161 VDD VSS sg13g2_decap_8
XFILLER_23_217 VDD VSS sg13g2_decap_8
XFILLER_16_280 VDD VSS sg13g2_decap_8
XFILLER_83_0 VDD VSS sg13g2_decap_8
XFILLER_31_294 VDD VSS sg13g2_decap_8
XFILLER_8_490 VDD VSS sg13g2_decap_8
XFILLER_59_637 VDD VSS sg13g2_decap_8
XFILLER_48_28 VDD VSS sg13g2_decap_8
XFILLER_86_434 VDD VSS sg13g2_decap_8
XFILLER_58_147 VDD VSS sg13g2_decap_8
XFILLER_39_350 VDD VSS sg13g2_decap_8
XFILLER_67_681 VDD VSS sg13g2_decap_8
XFILLER_82_651 VDD VSS sg13g2_decap_8
XFILLER_64_49 VDD VSS sg13g2_decap_8
XFILLER_54_364 VDD VSS sg13g2_decap_8
XFILLER_15_707 VDD VSS sg13g2_decap_8
XFILLER_27_567 VDD VSS sg13g2_decap_8
XFILLER_42_504 VDD VSS sg13g2_decap_8
XFILLER_81_161 VDD VSS sg13g2_decap_8
XFILLER_14_217 VDD VSS sg13g2_decap_8
XFILLER_50_581 VDD VSS sg13g2_decap_8
XFILLER_10_434 VDD VSS sg13g2_decap_8
XFILLER_13_42 VDD VSS sg13g2_decap_8
XFILLER_22_294 VDD VSS sg13g2_decap_8
XFILLER_6_427 VDD VSS sg13g2_decap_8
XFILLER_89_35 VDD VSS sg13g2_decap_8
XFILLER_2_644 VDD VSS sg13g2_decap_8
XFILLER_1_154 VDD VSS sg13g2_decap_8
XFILLER_89_294 VDD VSS sg13g2_decap_8
XFILLER_77_456 VDD VSS sg13g2_decap_4
XFILLER_49_147 VDD VSS sg13g2_decap_8
XFILLER_77_478 VDD VSS sg13g2_decap_8
XFILLER_92_448 VDD VSS sg13g2_decap_8
XFILLER_18_567 VDD VSS sg13g2_decap_8
XFILLER_33_504 VDD VSS sg13g2_decap_8
XFILLER_73_695 VDD VSS sg13g2_decap_8
XFILLER_72_161 VDD VSS sg13g2_decap_8
XFILLER_45_364 VDD VSS sg13g2_decap_8
XFILLER_60_301 VDD VSS sg13g2_decap_8
XFILLER_60_378 VDD VSS sg13g2_decap_8
XFILLER_13_294 VDD VSS sg13g2_decap_8
XFILLER_9_210 VDD VSS sg13g2_decap_8
XFILLER_41_581 VDD VSS sg13g2_decap_8
XFILLER_70_70 VDD VSS sg13g2_decap_8
XFILLER_9_287 VDD VSS sg13g2_decap_8
XFILLER_68_412 VDD VSS sg13g2_decap_8
XFILLER_95_231 VDD VSS sg13g2_decap_8
XFILLER_68_489 VDD VSS sg13g2_decap_8
XFILLER_83_448 VDD VSS sg13g2_decap_8
XFILLER_64_651 VDD VSS sg13g2_decap_8
XFILLER_63_161 VDD VSS sg13g2_decap_8
XFILLER_36_364 VDD VSS sg13g2_decap_8
XFILLER_51_301 VDD VSS sg13g2_decap_8
XFILLER_24_504 VDD VSS sg13g2_decap_8
XFILLER_51_378 VDD VSS sg13g2_decap_8
XFILLER_20_721 VDD VSS sg13g2_decap_8
XFILLER_32_581 VDD VSS sg13g2_decap_8
XFILLER_59_49 VDD VSS sg13g2_decap_8
XFILLER_87_721 VDD VSS sg13g2_decap_8
XFILLER_86_231 VDD VSS sg13g2_decap_8
XFILLER_59_434 VDD VSS sg13g2_decap_8
XFILLER_74_437 VDD VSS sg13g2_decap_8
XFILLER_74_448 VDD VSS sg13g2_decap_8
XFILLER_55_651 VDD VSS sg13g2_decap_8
XFILLER_70_610 VDD VSS sg13g2_decap_8
XFILLER_91_14 VDD VSS sg13g2_decap_8
XFILLER_27_364 VDD VSS sg13g2_decap_8
XFILLER_42_301 VDD VSS sg13g2_decap_8
XFILLER_54_161 VDD VSS sg13g2_decap_8
XFILLER_15_504 VDD VSS sg13g2_decap_8
XFILLER_70_687 VDD VSS sg13g2_decap_8
XFILLER_42_378 VDD VSS sg13g2_decap_8
XFILLER_30_518 VDD VSS sg13g2_decap_8
XFILLER_11_721 VDD VSS sg13g2_decap_8
XFILLER_24_63 VDD VSS sg13g2_decap_8
XFILLER_23_581 VDD VSS sg13g2_decap_8
XFILLER_7_714 VDD VSS sg13g2_decap_8
XFILLER_10_231 VDD VSS sg13g2_decap_8
XFILLER_6_224 VDD VSS sg13g2_decap_8
XFILLER_40_84 VDD VSS sg13g2_decap_8
XFILLER_2_441 VDD VSS sg13g2_decap_8
XFILLER_78_721 VDD VSS sg13g2_decap_8
XFILLER_77_253 VDD VSS sg13g2_decap_8
XFILLER_93_735 VDD VSS sg13g2_decap_8
XFILLER_65_448 VDD VSS sg13g2_decap_8
XFILLER_1_56 VDD VSS sg13g2_decap_8
XFILLER_92_245 VDD VSS sg13g2_decap_8
XFILLER_46_651 VDD VSS sg13g2_decap_8
XFILLER_65_70 VDD VSS sg13g2_decap_8
XFILLER_18_364 VDD VSS sg13g2_decap_8
XFILLER_33_301 VDD VSS sg13g2_decap_8
XFILLER_45_161 VDD VSS sg13g2_decap_8
XFILLER_73_492 VDD VSS sg13g2_decap_8
XFILLER_61_665 VDD VSS sg13g2_decap_8
XFILLER_33_378 VDD VSS sg13g2_decap_8
XFILLER_21_518 VDD VSS sg13g2_decap_8
XFILLER_60_175 VDD VSS sg13g2_decap_8
XFILLER_14_581 VDD VSS sg13g2_decap_8
XFILLER_81_91 VDD VSS sg13g2_decap_8
XFILLER_46_0 VDD VSS sg13g2_decap_8
XFILLER_88_518 VDD VSS sg13g2_decap_8
Xhold19 _64_/Y VDD VSS _79_/D sg13g2_dlygate4sd3_1
XFILLER_84_735 VDD VSS sg13g2_decap_8
XFILLER_68_286 VDD VSS sg13g2_decap_8
XFILLER_56_448 VDD VSS sg13g2_decap_8
XFILLER_83_245 VDD VSS sg13g2_decap_8
XFILLER_37_651 VDD VSS sg13g2_decap_8
XFILLER_71_429 VDD VSS sg13g2_decap_8
XFILLER_24_301 VDD VSS sg13g2_decap_8
XFILLER_36_161 VDD VSS sg13g2_decap_8
XFILLER_52_665 VDD VSS sg13g2_decap_8
XFILLER_12_518 VDD VSS sg13g2_decap_8
XFILLER_24_378 VDD VSS sg13g2_decap_8
XFILLER_61_28 VDD VSS sg13g2_decap_8
XFILLER_51_175 VDD VSS sg13g2_decap_8
XFILLER_20_595 VDD VSS sg13g2_decap_8
XFILLER_4_728 VDD VSS sg13g2_decap_8
XFILLER_10_21 VDD VSS sg13g2_decap_8
XFILLER_3_238 VDD VSS sg13g2_decap_8
XFILLER_79_518 VDD VSS sg13g2_decap_8
XFILLER_86_14 VDD VSS sg13g2_decap_8
XFILLER_10_98 VDD VSS sg13g2_decap_8
XFILLER_59_231 VDD VSS sg13g2_decap_8
XFILLER_87_595 VDD VSS sg13g2_decap_8
XFILLER_75_746 VDD VSS sg13g2_decap_8
XFILLER_19_63 VDD VSS sg13g2_decap_8
XFILLER_47_448 VDD VSS sg13g2_decap_8
XFILLER_28_651 VDD VSS sg13g2_decap_8
XFILLER_90_749 VDD VSS sg13g2_decap_8
XFILLER_15_301 VDD VSS sg13g2_decap_8
XFILLER_27_161 VDD VSS sg13g2_decap_8
XFILLER_35_84 VDD VSS sg13g2_decap_8
XFILLER_15_378 VDD VSS sg13g2_decap_8
XFILLER_43_665 VDD VSS sg13g2_decap_8
XFILLER_70_484 VDD VSS sg13g2_decap_8
XFILLER_30_315 VDD VSS sg13g2_decap_8
XFILLER_42_175 VDD VSS sg13g2_decap_8
XFILLER_7_511 VDD VSS sg13g2_decap_8
XFILLER_11_595 VDD VSS sg13g2_decap_8
XFILLER_7_588 VDD VSS sg13g2_decap_8
XFILLER_66_702 VDD VSS sg13g2_decap_8
XFILLER_93_532 VDD VSS sg13g2_decap_8
XFILLER_78_595 VDD VSS sg13g2_decap_8
XFILLER_65_245 VDD VSS sg13g2_decap_8
XFILLER_76_91 VDD VSS sg13g2_decap_8
XFILLER_38_448 VDD VSS sg13g2_decap_8
XFILLER_19_651 VDD VSS sg13g2_decap_8
XFILLER_18_161 VDD VSS sg13g2_decap_8
XFILLER_81_749 VDD VSS sg13g2_decap_8
XFILLER_80_259 VDD VSS sg13g2_decap_8
XFILLER_61_462 VDD VSS sg13g2_decap_8
XFILLER_34_665 VDD VSS sg13g2_decap_8
XFILLER_21_315 VDD VSS sg13g2_decap_8
XFILLER_33_175 VDD VSS sg13g2_decap_8
XFILLER_88_315 VDD VSS sg13g2_decap_8
XFILLER_69_573 VDD VSS sg13g2_decap_8
XFILLER_57_735 VDD VSS sg13g2_decap_8
XFILLER_56_28 VDD VSS sg13g2_decap_8
XFILLER_84_532 VDD VSS sg13g2_decap_8
XFILLER_72_705 VDD VSS sg13g2_decap_8
XFILLER_29_448 VDD VSS sg13g2_decap_8
XFILLER_56_245 VDD VSS sg13g2_decap_8
XFILLER_72_49 VDD VSS sg13g2_decap_8
XFILLER_52_462 VDD VSS sg13g2_decap_8
XFILLER_25_665 VDD VSS sg13g2_decap_8
XFILLER_40_602 VDD VSS sg13g2_decap_8
XFILLER_12_315 VDD VSS sg13g2_decap_8
XFILLER_24_175 VDD VSS sg13g2_decap_8
XFILLER_8_308 VDD VSS sg13g2_decap_8
XFILLER_40_679 VDD VSS sg13g2_decap_8
XFILLER_20_392 VDD VSS sg13g2_decap_8
XFILLER_4_525 VDD VSS sg13g2_decap_8
XFILLER_21_42 VDD VSS sg13g2_decap_8
XFILLER_79_315 VDD VSS sg13g2_decap_8
XFILLER_0_742 VDD VSS sg13g2_decap_8
XFILLER_94_329 VDD VSS sg13g2_decap_8
XFILLER_48_735 VDD VSS sg13g2_decap_8
XFILLER_75_543 VDD VSS sg13g2_decap_8
XFILLER_87_392 VDD VSS sg13g2_decap_8
XFILLER_47_245 VDD VSS sg13g2_decap_8
X_79__6 VDD VSS _79__6/L_HI sg13g2_tiehi
XFILLER_90_546 VDD VSS sg13g2_decap_8
XFILLER_62_259 VDD VSS sg13g2_decap_8
XFILLER_43_462 VDD VSS sg13g2_decap_8
XFILLER_16_665 VDD VSS sg13g2_decap_8
XFILLER_31_602 VDD VSS sg13g2_decap_8
XFILLER_70_270 VDD VSS sg13g2_decap_8
XFILLER_15_175 VDD VSS sg13g2_decap_8
XFILLER_30_112 VDD VSS sg13g2_decap_8
XFILLER_87_7 VDD VSS sg13g2_decap_8
XFILLER_31_679 VDD VSS sg13g2_decap_8
XFILLER_11_392 VDD VSS sg13g2_decap_8
XFILLER_30_189 VDD VSS sg13g2_decap_8
XFILLER_7_77 VDD VSS sg13g2_decap_8
XFILLER_7_385 VDD VSS sg13g2_decap_8
XFILLER_85_329 VDD VSS sg13g2_decap_8
XFILLER_39_735 VDD VSS sg13g2_decap_8
XFILLER_78_392 VDD VSS sg13g2_decap_8
XFILLER_38_245 VDD VSS sg13g2_decap_8
XFILLER_66_576 VDD VSS sg13g2_decap_8
XFILLER_81_546 VDD VSS sg13g2_decap_8
XFILLER_54_749 VDD VSS sg13g2_decap_8
XFILLER_53_259 VDD VSS sg13g2_decap_8
XFILLER_22_602 VDD VSS sg13g2_decap_8
XFILLER_21_112 VDD VSS sg13g2_decap_8
XFILLER_34_462 VDD VSS sg13g2_decap_8
XFILLER_22_679 VDD VSS sg13g2_decap_8
XFILLER_21_189 VDD VSS sg13g2_decap_8
XFILLER_89_602 VDD VSS sg13g2_decap_8
XFILLER_88_112 VDD VSS sg13g2_decap_8
XFILLER_1_539 VDD VSS sg13g2_decap_8
XFILLER_89_679 VDD VSS sg13g2_decap_8
XFILLER_88_189 VDD VSS sg13g2_decap_8
XFILLER_67_49 VDD VSS sg13g2_decap_8
XFILLER_57_532 VDD VSS sg13g2_decap_8
XFILLER_29_245 VDD VSS sg13g2_decap_8
XFILLER_72_502 VDD VSS sg13g2_decap_8
XFILLER_45_749 VDD VSS sg13g2_decap_8
XFILLER_72_579 VDD VSS sg13g2_decap_8
XFILLER_16_42 VDD VSS sg13g2_decap_8
XFILLER_44_259 VDD VSS sg13g2_decap_8
XFILLER_13_602 VDD VSS sg13g2_decap_8
XFILLER_25_462 VDD VSS sg13g2_decap_8
XFILLER_12_112 VDD VSS sg13g2_decap_8
XFILLER_13_679 VDD VSS sg13g2_decap_8
XFILLER_8_105 VDD VSS sg13g2_decap_8
XFILLER_40_476 VDD VSS sg13g2_decap_8
XFILLER_12_189 VDD VSS sg13g2_decap_8
XFILLER_32_63 VDD VSS sg13g2_decap_8
XFILLER_4_322 VDD VSS sg13g2_decap_8
XFILLER_79_112 VDD VSS sg13g2_decap_8
XFILLER_4_399 VDD VSS sg13g2_decap_8
XFILLER_95_616 VDD VSS sg13g2_decap_8
XFILLER_94_126 VDD VSS sg13g2_decap_8
XFILLER_79_189 VDD VSS sg13g2_decap_8
XFILLER_48_532 VDD VSS sg13g2_decap_8
XFILLER_75_395 VDD VSS sg13g2_decap_8
XFILLER_36_749 VDD VSS sg13g2_decap_8
XFILLER_63_557 VDD VSS sg13g2_decap_8
XFILLER_90_343 VDD VSS sg13g2_decap_8
XFILLER_35_259 VDD VSS sg13g2_decap_8
XFILLER_73_70 VDD VSS sg13g2_decap_8
XFILLER_16_462 VDD VSS sg13g2_decap_8
XFILLER_71_590 VDD VSS sg13g2_decap_8
XFILLER_31_476 VDD VSS sg13g2_decap_8
XFILLER_8_672 VDD VSS sg13g2_decap_8
XFILLER_7_182 VDD VSS sg13g2_decap_8
XFILLER_86_616 VDD VSS sg13g2_decap_8
XFILLER_58_329 VDD VSS sg13g2_decap_8
XFILLER_85_126 VDD VSS sg13g2_decap_8
XFILLER_39_532 VDD VSS sg13g2_decap_8
XFILLER_94_693 VDD VSS sg13g2_decap_8
XFILLER_54_546 VDD VSS sg13g2_decap_8
XFILLER_27_749 VDD VSS sg13g2_decap_8
XFILLER_81_343 VDD VSS sg13g2_decap_8
XFILLER_26_259 VDD VSS sg13g2_decap_8
XFILLER_10_616 VDD VSS sg13g2_decap_8
XFILLER_22_476 VDD VSS sg13g2_decap_8
XFILLER_6_609 VDD VSS sg13g2_decap_8
XFILLER_5_119 VDD VSS sg13g2_decap_8
XFILLER_1_336 VDD VSS sg13g2_decap_8
XFILLER_89_476 VDD VSS sg13g2_decap_8
XFILLER_49_329 VDD VSS sg13g2_decap_8
XFILLER_76_126 VDD VSS sg13g2_decap_8
XFILLER_94_14 VDD VSS sg13g2_decap_8
XFILLER_85_693 VDD VSS sg13g2_decap_8
XFILLER_27_63 VDD VSS sg13g2_decap_8
XFILLER_18_749 VDD VSS sg13g2_decap_8
XFILLER_45_546 VDD VSS sg13g2_decap_8
XFILLER_72_332 VDD VSS sg13g2_decap_4
XFILLER_17_259 VDD VSS sg13g2_decap_8
XFILLER_13_476 VDD VSS sg13g2_decap_8
XFILLER_43_84 VDD VSS sg13g2_decap_8
XFILLER_40_273 VDD VSS sg13g2_decap_8
XFILLER_9_469 VDD VSS sg13g2_decap_8
XFILLER_5_686 VDD VSS sg13g2_decap_8
XFILLER_4_196 VDD VSS sg13g2_decap_8
XFILLER_4_56 VDD VSS sg13g2_decap_8
XFILLER_95_413 VDD VSS sg13g2_decap_8
XFILLER_68_70 VDD VSS sg13g2_decap_8
XFILLER_67_126 VDD VSS sg13g2_decap_8
XFILLER_76_671 VDD VSS sg13g2_decap_8
XFILLER_91_630 VDD VSS sg13g2_decap_8
XFILLER_90_140 VDD VSS sg13g2_decap_8
XFILLER_63_343 VDD VSS sg13g2_decap_8
XFILLER_84_91 VDD VSS sg13g2_decap_8
XFILLER_36_546 VDD VSS sg13g2_decap_8
XFILLER_31_273 VDD VSS sg13g2_decap_8
XFILLER_76_0 VDD VSS sg13g2_decap_8
XFILLER_86_413 VDD VSS sg13g2_decap_8
XFILLER_59_616 VDD VSS sg13g2_decap_8
XFILLER_58_126 VDD VSS sg13g2_decap_8
XFILLER_67_660 VDD VSS sg13g2_decap_8
XFILLER_94_490 VDD VSS sg13g2_decap_8
XFILLER_82_630 VDD VSS sg13g2_decap_8
XFILLER_81_140 VDD VSS sg13g2_decap_8
XFILLER_64_28 VDD VSS sg13g2_decap_4
XFILLER_54_343 VDD VSS sg13g2_decap_8
XFILLER_27_546 VDD VSS sg13g2_decap_8
XFILLER_50_560 VDD VSS sg13g2_decap_8
XFILLER_80_49 VDD VSS sg13g2_decap_8
XFILLER_10_413 VDD VSS sg13g2_decap_8
XFILLER_13_21 VDD VSS sg13g2_decap_8
XFILLER_22_273 VDD VSS sg13g2_decap_8
XFILLER_6_406 VDD VSS sg13g2_decap_8
XFILLER_89_14 VDD VSS sg13g2_decap_8
XFILLER_13_98 VDD VSS sg13g2_decap_8
XFILLER_2_623 VDD VSS sg13g2_decap_8
XFILLER_1_133 VDD VSS sg13g2_decap_8
XFILLER_89_273 VDD VSS sg13g2_decap_8
XFILLER_77_435 VDD VSS sg13g2_decap_8
XFILLER_49_126 VDD VSS sg13g2_decap_8
XFILLER_65_619 VDD VSS sg13g2_decap_8
XFILLER_92_427 VDD VSS sg13g2_decap_8
XFILLER_58_693 VDD VSS sg13g2_decap_8
XFILLER_38_84 VDD VSS sg13g2_decap_8
XFILLER_85_490 VDD VSS sg13g2_decap_8
XFILLER_72_140 VDD VSS sg13g2_decap_8
XFILLER_45_343 VDD VSS sg13g2_decap_8
XFILLER_18_546 VDD VSS sg13g2_decap_8
XFILLER_73_674 VDD VSS sg13g2_decap_8
XFILLER_60_357 VDD VSS sg13g2_decap_8
XFILLER_41_560 VDD VSS sg13g2_decap_8
XFILLER_13_273 VDD VSS sg13g2_decap_8
XFILLER_9_266 VDD VSS sg13g2_decap_8
XFILLER_5_483 VDD VSS sg13g2_decap_8
XFILLER_79_91 VDD VSS sg13g2_decap_8
XFILLER_95_210 VDD VSS sg13g2_decap_8
XFILLER_68_468 VDD VSS sg13g2_decap_8
XFILLER_95_287 VDD VSS sg13g2_decap_8
XFILLER_83_427 VDD VSS sg13g2_decap_8
XFILLER_49_693 VDD VSS sg13g2_decap_8
XFILLER_64_630 VDD VSS sg13g2_decap_8
XFILLER_36_343 VDD VSS sg13g2_decap_8
XFILLER_63_140 VDD VSS sg13g2_decap_8
XFILLER_51_357 VDD VSS sg13g2_decap_8
XFILLER_20_700 VDD VSS sg13g2_decap_8
XFILLER_32_560 VDD VSS sg13g2_decap_8
XFILLER_59_28 VDD VSS sg13g2_decap_8
XFILLER_87_700 VDD VSS sg13g2_decap_8
XFILLER_59_413 VDD VSS sg13g2_decap_8
XFILLER_86_210 VDD VSS sg13g2_decap_8
XFILLER_86_287 VDD VSS sg13g2_decap_8
XFILLER_74_416 VDD VSS sg13g2_decap_8
XFILLER_55_630 VDD VSS sg13g2_decap_8
XFILLER_27_343 VDD VSS sg13g2_decap_8
XFILLER_54_140 VDD VSS sg13g2_decap_8
XFILLER_70_666 VDD VSS sg13g2_decap_8
XFILLER_11_700 VDD VSS sg13g2_decap_8
XFILLER_24_42 VDD VSS sg13g2_decap_8
XFILLER_42_357 VDD VSS sg13g2_decap_8
XFILLER_23_560 VDD VSS sg13g2_decap_8
XFILLER_10_210 VDD VSS sg13g2_decap_8
XFILLER_6_203 VDD VSS sg13g2_decap_8
XFILLER_10_287 VDD VSS sg13g2_decap_8
XFILLER_40_63 VDD VSS sg13g2_decap_8
XFILLER_2_420 VDD VSS sg13g2_decap_8
XFILLER_6_0 VDD VSS sg13g2_decap_8
XFILLER_78_700 VDD VSS sg13g2_decap_8
XFILLER_77_210 VDD VSS sg13g2_decap_8
XFILLER_2_497 VDD VSS sg13g2_decap_8
XFILLER_93_714 VDD VSS sg13g2_decap_8
XFILLER_92_224 VDD VSS sg13g2_decap_8
XFILLER_65_427 VDD VSS sg13g2_decap_8
XFILLER_1_35 VDD VSS sg13g2_decap_8
XFILLER_58_490 VDD VSS sg13g2_decap_8
XFILLER_46_630 VDD VSS sg13g2_decap_8
XFILLER_18_343 VDD VSS sg13g2_decap_8
XFILLER_73_471 VDD VSS sg13g2_decap_8
XFILLER_45_140 VDD VSS sg13g2_decap_8
XFILLER_61_644 VDD VSS sg13g2_decap_8
XFILLER_33_357 VDD VSS sg13g2_decap_8
XFILLER_60_154 VDD VSS sg13g2_decap_8
XFILLER_81_70 VDD VSS sg13g2_decap_8
XFILLER_14_560 VDD VSS sg13g2_decap_8
XFILLER_5_280 VDD VSS sg13g2_decap_8
XFILLER_69_755 VDD VSS sg13g2_fill_2
XFILLER_39_0 VDD VSS sg13g2_decap_8
XFILLER_84_714 VDD VSS sg13g2_decap_8
XFILLER_68_265 VDD VSS sg13g2_decap_8
XFILLER_83_224 VDD VSS sg13g2_decap_8
XFILLER_56_427 VDD VSS sg13g2_decap_8
XFILLER_49_490 VDD VSS sg13g2_decap_8
XFILLER_37_630 VDD VSS sg13g2_decap_8
XFILLER_36_140 VDD VSS sg13g2_decap_8
XFILLER_52_644 VDD VSS sg13g2_decap_8
XFILLER_24_357 VDD VSS sg13g2_decap_8
XFILLER_51_154 VDD VSS sg13g2_decap_8
XFILLER_20_574 VDD VSS sg13g2_decap_8
XFILLER_4_707 VDD VSS sg13g2_decap_8
XFILLER_3_217 VDD VSS sg13g2_decap_8
XFILLER_10_77 VDD VSS sg13g2_decap_8
XFILLER_59_210 VDD VSS sg13g2_decap_8
XFILLER_87_574 VDD VSS sg13g2_decap_8
XFILLER_75_725 VDD VSS sg13g2_decap_8
XFILLER_19_42 VDD VSS sg13g2_decap_8
XFILLER_47_427 VDD VSS sg13g2_decap_8
XFILLER_59_287 VDD VSS sg13g2_decap_8
XFILLER_74_257 VDD VSS sg13g2_decap_8
XFILLER_74_224 VDD VSS sg13g2_decap_8
XFILLER_74_235 VDD VSS sg13g2_fill_1
XFILLER_28_630 VDD VSS sg13g2_decap_8
XFILLER_90_728 VDD VSS sg13g2_decap_8
XFILLER_74_279 VDD VSS sg13g2_decap_8
XFILLER_27_140 VDD VSS sg13g2_decap_8
XFILLER_43_644 VDD VSS sg13g2_decap_8
XFILLER_35_63 VDD VSS sg13g2_decap_8
XFILLER_15_357 VDD VSS sg13g2_decap_8
XFILLER_42_154 VDD VSS sg13g2_decap_8
XFILLER_11_574 VDD VSS sg13g2_decap_8
XFILLER_7_567 VDD VSS sg13g2_decap_8
XFILLER_51_84 VDD VSS sg13g2_decap_8
XFILLER_32_7 VDD VSS sg13g2_decap_8
XFILLER_2_294 VDD VSS sg13g2_decap_8
XFILLER_93_511 VDD VSS sg13g2_decap_8
XFILLER_78_574 VDD VSS sg13g2_decap_8
XFILLER_76_70 VDD VSS sg13g2_decap_8
XFILLER_38_427 VDD VSS sg13g2_decap_8
XFILLER_65_224 VDD VSS sg13g2_decap_8
XFILLER_19_630 VDD VSS sg13g2_decap_8
XFILLER_93_588 VDD VSS sg13g2_decap_8
XFILLER_81_728 VDD VSS sg13g2_decap_8
XFILLER_18_140 VDD VSS sg13g2_decap_8
XFILLER_80_238 VDD VSS sg13g2_decap_8
XFILLER_34_644 VDD VSS sg13g2_decap_8
XFILLER_33_154 VDD VSS sg13g2_decap_8
XFILLER_61_441 VDD VSS sg13g2_decap_8
XFILLER_92_91 VDD VSS sg13g2_decap_8
XFILLER_69_552 VDD VSS sg13g2_decap_8
XFILLER_84_511 VDD VSS sg13g2_decap_8
XFILLER_57_714 VDD VSS sg13g2_decap_8
XFILLER_29_427 VDD VSS sg13g2_decap_8
XFILLER_56_224 VDD VSS sg13g2_decap_8
XFILLER_84_588 VDD VSS sg13g2_decap_8
XFILLER_71_249 VDD VSS sg13g2_decap_8
XFILLER_25_644 VDD VSS sg13g2_decap_8
XFILLER_72_28 VDD VSS sg13g2_decap_8
XFILLER_52_441 VDD VSS sg13g2_decap_8
XFILLER_24_154 VDD VSS sg13g2_decap_8
XFILLER_40_658 VDD VSS sg13g2_decap_8
XFILLER_21_21 VDD VSS sg13g2_decap_8
XFILLER_20_371 VDD VSS sg13g2_decap_8
XFILLER_4_504 VDD VSS sg13g2_decap_8
XFILLER_21_98 VDD VSS sg13g2_decap_8
XIO_BOND_vdd_pads\[0\].vdd_pad VDD bondpad_70x70_novias
XFILLER_0_721 VDD VSS sg13g2_decap_8
XFILLER_94_308 VDD VSS sg13g2_decap_8
XFILLER_75_522 VDD VSS sg13g2_decap_8
XFILLER_87_371 VDD VSS sg13g2_decap_8
XFILLER_48_714 VDD VSS sg13g2_decap_8
XFILLER_47_224 VDD VSS sg13g2_decap_8
XFILLER_90_525 VDD VSS sg13g2_decap_8
XFILLER_75_599 VDD VSS sg13g2_decap_8
XFILLER_63_739 VDD VSS sg13g2_decap_8
XFILLER_62_238 VDD VSS sg13g2_decap_8
XFILLER_46_84 VDD VSS sg13g2_decap_8
XFILLER_43_441 VDD VSS sg13g2_decap_8
XFILLER_16_644 VDD VSS sg13g2_decap_8
XFILLER_15_154 VDD VSS sg13g2_decap_8
XFILLER_31_658 VDD VSS sg13g2_decap_8
XFILLER_30_168 VDD VSS sg13g2_decap_8
XFILLER_11_371 VDD VSS sg13g2_decap_8
XFILLER_7_364 VDD VSS sg13g2_decap_8
XFILLER_7_56 VDD VSS sg13g2_decap_8
XFILLER_3_581 VDD VSS sg13g2_decap_8
XFILLER_85_308 VDD VSS sg13g2_decap_8
XFILLER_78_371 VDD VSS sg13g2_decap_8
XFILLER_87_91 VDD VSS sg13g2_decap_8
XFILLER_39_714 VDD VSS sg13g2_decap_8
XFILLER_66_555 VDD VSS sg13g2_decap_8
XFILLER_38_224 VDD VSS sg13g2_decap_8
XFILLER_54_728 VDD VSS sg13g2_decap_8
XFILLER_26_419 VDD VSS sg13g2_decap_8
XFILLER_81_525 VDD VSS sg13g2_decap_8
XFILLER_93_385 VDD VSS sg13g2_decap_8
XFILLER_53_238 VDD VSS sg13g2_decap_8
XFILLER_34_441 VDD VSS sg13g2_decap_8
XFILLER_22_658 VDD VSS sg13g2_decap_8
XFILLER_21_168 VDD VSS sg13g2_decap_8
XFILLER_1_518 VDD VSS sg13g2_decap_8
Xoutputs\[3\].output_pad _79_/Q IOVDD IOVSS output_PAD[3] VDD VSS sg13g2_IOPadOut30mA
XFILLER_89_658 VDD VSS sg13g2_decap_8
XFILLER_67_28 VDD VSS sg13g2_decap_8
XFILLER_88_168 VDD VSS sg13g2_decap_8
XFILLER_57_511 VDD VSS sg13g2_decap_8
XFILLER_29_224 VDD VSS sg13g2_decap_8
XFILLER_57_588 VDD VSS sg13g2_decap_8
XFILLER_45_728 VDD VSS sg13g2_decap_8
XFILLER_84_385 VDD VSS sg13g2_decap_8
XFILLER_83_49 VDD VSS sg13g2_decap_8
XFILLER_44_238 VDD VSS sg13g2_decap_8
XFILLER_72_558 VDD VSS sg13g2_decap_8
XFILLER_16_21 VDD VSS sg13g2_decap_8
XFILLER_25_441 VDD VSS sg13g2_decap_8
XFILLER_13_658 VDD VSS sg13g2_decap_8
XFILLER_16_98 VDD VSS sg13g2_decap_8
XFILLER_12_168 VDD VSS sg13g2_decap_8
XFILLER_40_455 VDD VSS sg13g2_decap_8
XFILLER_32_42 VDD VSS sg13g2_decap_8
XFILLER_4_301 VDD VSS sg13g2_decap_8
XFILLER_4_378 VDD VSS sg13g2_decap_8
XFILLER_79_168 VDD VSS sg13g2_decap_8
XFILLER_94_105 VDD VSS sg13g2_decap_8
XFILLER_48_511 VDD VSS sg13g2_decap_8
XFILLER_0_595 VDD VSS sg13g2_decap_8
XFILLER_75_341 VDD VSS sg13g2_decap_8
XFILLER_48_588 VDD VSS sg13g2_decap_8
XFILLER_36_728 VDD VSS sg13g2_decap_8
XFILLER_63_536 VDD VSS sg13g2_decap_8
XFILLER_90_322 VDD VSS sg13g2_decap_8
XFILLER_75_374 VDD VSS sg13g2_decap_8
XFILLER_35_238 VDD VSS sg13g2_decap_8
XFILLER_16_441 VDD VSS sg13g2_decap_8
XFILLER_90_399 VDD VSS sg13g2_decap_8
XFILLER_31_455 VDD VSS sg13g2_decap_8
XFILLER_8_651 VDD VSS sg13g2_decap_8
XFILLER_7_161 VDD VSS sg13g2_decap_8
XFILLER_85_105 VDD VSS sg13g2_decap_8
XFILLER_21_0 VDD VSS sg13g2_decap_8
XFILLER_58_308 VDD VSS sg13g2_decap_8
XFILLER_39_511 VDD VSS sg13g2_decap_8
XFILLER_94_672 VDD VSS sg13g2_decap_8
XFILLER_93_182 VDD VSS sg13g2_decap_8
XFILLER_81_322 VDD VSS sg13g2_decap_8
XFILLER_66_385 VDD VSS sg13g2_decap_8
XFILLER_54_525 VDD VSS sg13g2_decap_8
XFILLER_27_728 VDD VSS sg13g2_decap_8
XFILLER_39_588 VDD VSS sg13g2_decap_8
XFILLER_26_238 VDD VSS sg13g2_decap_8
XFILLER_81_399 VDD VSS sg13g2_decap_8
XFILLER_50_742 VDD VSS sg13g2_decap_8
XFILLER_22_455 VDD VSS sg13g2_decap_8
XFILLER_78_49 VDD VSS sg13g2_decap_8
XFILLER_1_315 VDD VSS sg13g2_decap_8
XFILLER_89_455 VDD VSS sg13g2_decap_8
XFILLER_77_639 VDD VSS sg13g2_decap_8
XFILLER_76_105 VDD VSS sg13g2_decap_8
XFILLER_49_308 VDD VSS sg13g2_decap_8
XFILLER_92_609 VDD VSS sg13g2_decap_8
XFILLER_85_672 VDD VSS sg13g2_decap_8
XFILLER_91_119 VDD VSS sg13g2_decap_8
XFILLER_84_182 VDD VSS sg13g2_decap_8
XFILLER_72_311 VDD VSS sg13g2_decap_8
XFILLER_27_42 VDD VSS sg13g2_decap_8
XFILLER_57_385 VDD VSS sg13g2_decap_8
XFILLER_18_728 VDD VSS sg13g2_decap_8
XFILLER_45_525 VDD VSS sg13g2_decap_8
XFILLER_17_238 VDD VSS sg13g2_decap_8
XFILLER_72_388 VDD VSS sg13g2_decap_8
XFILLER_60_539 VDD VSS sg13g2_decap_8
XFILLER_41_742 VDD VSS sg13g2_decap_8
XFILLER_13_455 VDD VSS sg13g2_decap_8
XFILLER_43_63 VDD VSS sg13g2_decap_8
XFILLER_40_252 VDD VSS sg13g2_decap_8
XFILLER_9_448 VDD VSS sg13g2_decap_8
XFILLER_5_665 VDD VSS sg13g2_decap_8
XFILLER_4_175 VDD VSS sg13g2_decap_8
XFILLER_4_35 VDD VSS sg13g2_decap_8
XFILLER_67_105 VDD VSS sg13g2_decap_8
XFILLER_83_609 VDD VSS sg13g2_decap_8
XFILLER_76_650 VDD VSS sg13g2_decap_8
XFILLER_95_469 VDD VSS sg13g2_decap_8
XFILLER_0_392 VDD VSS sg13g2_decap_8
XFILLER_82_119 VDD VSS sg13g2_decap_8
XFILLER_63_322 VDD VSS sg13g2_decap_8
XFILLER_48_385 VDD VSS sg13g2_decap_8
XFILLER_36_525 VDD VSS sg13g2_decap_8
XFILLER_75_193 VDD VSS sg13g2_decap_8
XFILLER_84_70 VDD VSS sg13g2_decap_8
XFILLER_91_686 VDD VSS sg13g2_decap_8
XFILLER_90_196 VDD VSS sg13g2_decap_8
XFILLER_63_399 VDD VSS sg13g2_decap_8
XFILLER_51_539 VDD VSS sg13g2_decap_8
XFILLER_32_742 VDD VSS sg13g2_decap_8
XFILLER_31_252 VDD VSS sg13g2_decap_8
XFILLER_69_0 VDD VSS sg13g2_decap_8
XFILLER_58_105 VDD VSS sg13g2_decap_8
XFILLER_74_609 VDD VSS sg13g2_decap_8
XFILLER_86_469 VDD VSS sg13g2_decap_8
XFILLER_73_119 VDD VSS sg13g2_decap_8
XFILLER_39_385 VDD VSS sg13g2_decap_8
XFILLER_27_525 VDD VSS sg13g2_decap_8
XFILLER_66_182 VDD VSS sg13g2_decap_8
XFILLER_54_322 VDD VSS sg13g2_decap_8
XFILLER_82_686 VDD VSS sg13g2_decap_8
XFILLER_81_196 VDD VSS sg13g2_decap_8
XFILLER_54_399 VDD VSS sg13g2_decap_8
XFILLER_23_742 VDD VSS sg13g2_decap_8
XFILLER_42_539 VDD VSS sg13g2_decap_8
XFILLER_80_28 VDD VSS sg13g2_decap_8
XFILLER_22_252 VDD VSS sg13g2_decap_8
XFILLER_10_469 VDD VSS sg13g2_decap_8
XFILLER_13_77 VDD VSS sg13g2_decap_8
XFILLER_2_602 VDD VSS sg13g2_decap_8
XFILLER_1_112 VDD VSS sg13g2_decap_8
XFILLER_89_252 VDD VSS sg13g2_decap_8
XFILLER_2_679 VDD VSS sg13g2_decap_8
XFILLER_49_105 VDD VSS sg13g2_decap_8
XFILLER_1_189 VDD VSS sg13g2_decap_8
XFILLER_92_406 VDD VSS sg13g2_decap_8
XFILLER_38_63 VDD VSS sg13g2_decap_8
XFILLER_64_119 VDD VSS sg13g2_decap_8
XFILLER_58_672 VDD VSS sg13g2_decap_8
XFILLER_18_525 VDD VSS sg13g2_decap_8
XFILLER_73_653 VDD VSS sg13g2_decap_8
XFILLER_45_322 VDD VSS sg13g2_decap_8
XFILLER_57_182 VDD VSS sg13g2_decap_8
XFILLER_72_196 VDD VSS sg13g2_decap_8
XFILLER_54_84 VDD VSS sg13g2_decap_8
XFILLER_45_399 VDD VSS sg13g2_decap_8
XFILLER_60_336 VDD VSS sg13g2_decap_8
XFILLER_14_742 VDD VSS sg13g2_decap_8
XFILLER_26_580 VDD VSS sg13g2_decap_8
XFILLER_33_539 VDD VSS sg13g2_decap_8
XFILLER_13_252 VDD VSS sg13g2_decap_8
XFILLER_9_245 VDD VSS sg13g2_decap_8
XFILLER_62_7 VDD VSS sg13g2_decap_8
XFILLER_5_462 VDD VSS sg13g2_decap_8
XFILLER_79_70 VDD VSS sg13g2_decap_8
XFILLER_68_447 VDD VSS sg13g2_fill_2
XFILLER_95_266 VDD VSS sg13g2_decap_8
XFILLER_83_406 VDD VSS sg13g2_decap_8
XFILLER_56_609 VDD VSS sg13g2_decap_8
XFILLER_95_91 VDD VSS sg13g2_decap_8
XFILLER_49_672 VDD VSS sg13g2_decap_8
XFILLER_55_119 VDD VSS sg13g2_decap_8
XFILLER_36_322 VDD VSS sg13g2_decap_8
XFILLER_48_182 VDD VSS sg13g2_decap_8
XFILLER_64_686 VDD VSS sg13g2_decap_8
XFILLER_91_483 VDD VSS sg13g2_decap_8
XFILLER_63_196 VDD VSS sg13g2_decap_8
XFILLER_36_399 VDD VSS sg13g2_decap_8
XFILLER_51_336 VDD VSS sg13g2_decap_8
XFILLER_24_539 VDD VSS sg13g2_decap_8
XFILLER_20_756 VDD VSS sg13g2_fill_1
XFILLER_87_756 VDD VSS sg13g2_fill_1
XFILLER_86_266 VDD VSS sg13g2_decap_8
XFILLER_75_28 VDD VSS sg13g2_fill_2
XFILLER_47_609 VDD VSS sg13g2_decap_8
XFILLER_59_469 VDD VSS sg13g2_decap_8
XFILLER_75_39 VDD VSS sg13g2_decap_8
XFILLER_46_119 VDD VSS sg13g2_decap_8
XFILLER_27_322 VDD VSS sg13g2_decap_8
XFILLER_39_182 VDD VSS sg13g2_decap_8
XFILLER_55_686 VDD VSS sg13g2_decap_8
XFILLER_82_483 VDD VSS sg13g2_decap_8
XFILLER_70_645 VDD VSS sg13g2_decap_8
XFILLER_91_49 VDD VSS sg13g2_decap_8
XFILLER_27_399 VDD VSS sg13g2_decap_8
XFILLER_42_336 VDD VSS sg13g2_decap_8
XFILLER_54_196 VDD VSS sg13g2_decap_8
XFILLER_15_539 VDD VSS sg13g2_decap_8
XFILLER_24_21 VDD VSS sg13g2_decap_8
XFILLER_11_756 VDD VSS sg13g2_fill_1
XFILLER_24_98 VDD VSS sg13g2_decap_8
XFILLER_7_749 VDD VSS sg13g2_decap_8
XFILLER_10_266 VDD VSS sg13g2_decap_8
XFILLER_6_259 VDD VSS sg13g2_decap_8
XFILLER_40_42 VDD VSS sg13g2_decap_8
XFILLER_2_476 VDD VSS sg13g2_decap_8
XFILLER_78_756 VDD VSS sg13g2_fill_1
XFILLER_1_14 VDD VSS sg13g2_decap_8
XFILLER_49_84 VDD VSS sg13g2_decap_8
XFILLER_38_609 VDD VSS sg13g2_decap_8
XFILLER_92_203 VDD VSS sg13g2_decap_8
XFILLER_77_288 VDD VSS sg13g2_decap_8
XFILLER_65_406 VDD VSS sg13g2_decap_8
XFILLER_37_119 VDD VSS sg13g2_decap_8
XFILLER_18_322 VDD VSS sg13g2_decap_8
XFILLER_46_686 VDD VSS sg13g2_decap_8
XFILLER_61_623 VDD VSS sg13g2_decap_8
XFILLER_18_399 VDD VSS sg13g2_decap_8
XFILLER_33_336 VDD VSS sg13g2_decap_8
XFILLER_45_196 VDD VSS sg13g2_decap_8
XFILLER_60_133 VDD VSS sg13g2_decap_8
XFILLER_69_734 VDD VSS sg13g2_decap_8
XFILLER_68_244 VDD VSS sg13g2_decap_8
XFILLER_29_609 VDD VSS sg13g2_decap_8
XFILLER_83_203 VDD VSS sg13g2_decap_8
Xoutputs\[8\].output_pad outputs\[8\].output_pad/c2p IOVDD IOVSS output_PAD[8] VDD
+ VSS sg13g2_IOPadOut30mA
XFILLER_28_119 VDD VSS sg13g2_decap_8
XFILLER_56_406 VDD VSS sg13g2_decap_8
X_79_ _79__6/L_HI VSS VDD _79_/D _79_/Q _79_/CLK sg13g2_dfrbpq_1
XFILLER_37_686 VDD VSS sg13g2_decap_8
XFILLER_64_483 VDD VSS sg13g2_decap_8
XFILLER_91_280 VDD VSS sg13g2_decap_8
XFILLER_52_623 VDD VSS sg13g2_decap_8
XFILLER_24_336 VDD VSS sg13g2_decap_8
XFILLER_36_196 VDD VSS sg13g2_decap_8
XFILLER_51_133 VDD VSS sg13g2_decap_8
XFILLER_20_553 VDD VSS sg13g2_decap_8
XFILLER_10_56 VDD VSS sg13g2_decap_8
XFILLER_87_553 VDD VSS sg13g2_decap_8
XFILLER_75_704 VDD VSS sg13g2_decap_8
XFILLER_86_49 VDD VSS sg13g2_decap_8
XFILLER_19_21 VDD VSS sg13g2_decap_8
XFILLER_74_203 VDD VSS sg13g2_decap_8
XFILLER_19_119 VDD VSS sg13g2_decap_8
XFILLER_47_406 VDD VSS sg13g2_decap_8
XFILLER_59_266 VDD VSS sg13g2_decap_8
XFILLER_19_98 VDD VSS sg13g2_decap_8
XFILLER_90_707 VDD VSS sg13g2_decap_8
XFILLER_82_280 VDD VSS sg13g2_decap_8
XFILLER_55_483 VDD VSS sg13g2_decap_8
XFILLER_35_42 VDD VSS sg13g2_decap_8
XFILLER_15_336 VDD VSS sg13g2_decap_8
XFILLER_28_686 VDD VSS sg13g2_decap_8
XFILLER_43_623 VDD VSS sg13g2_decap_8
XFILLER_70_453 VDD VSS sg13g2_fill_2
XFILLER_27_196 VDD VSS sg13g2_decap_8
XFILLER_42_133 VDD VSS sg13g2_decap_8
XFILLER_11_553 VDD VSS sg13g2_decap_8
XFILLER_51_63 VDD VSS sg13g2_decap_8
XFILLER_7_546 VDD VSS sg13g2_decap_8
XFILLER_2_273 VDD VSS sg13g2_decap_8
XFILLER_78_553 VDD VSS sg13g2_decap_8
XFILLER_25_7 VDD VSS sg13g2_decap_8
XFILLER_66_737 VDD VSS sg13g2_decap_8
XFILLER_65_203 VDD VSS sg13g2_decap_8
XFILLER_38_406 VDD VSS sg13g2_decap_8
XFILLER_93_567 VDD VSS sg13g2_decap_8
XFILLER_81_707 VDD VSS sg13g2_decap_8
XFILLER_80_217 VDD VSS sg13g2_decap_8
XFILLER_46_483 VDD VSS sg13g2_decap_8
XFILLER_61_420 VDD VSS sg13g2_decap_8
XFILLER_19_686 VDD VSS sg13g2_decap_8
XFILLER_34_623 VDD VSS sg13g2_decap_8
XFILLER_92_70 VDD VSS sg13g2_decap_8
XFILLER_18_196 VDD VSS sg13g2_decap_8
XFILLER_33_133 VDD VSS sg13g2_decap_8
XFILLER_61_497 VDD VSS sg13g2_decap_8
XFILLER_51_0 VDD VSS sg13g2_decap_8
XFILLER_69_531 VDD VSS sg13g2_decap_8
XFILLER_29_406 VDD VSS sg13g2_decap_8
XFILLER_56_203 VDD VSS sg13g2_decap_8
XFILLER_84_567 VDD VSS sg13g2_decap_8
XFILLER_71_228 VDD VSS sg13g2_decap_8
XFILLER_64_280 VDD VSS sg13g2_decap_8
XFILLER_52_420 VDD VSS sg13g2_decap_8
XFILLER_25_623 VDD VSS sg13g2_decap_8
XFILLER_37_483 VDD VSS sg13g2_decap_8
XFILLER_24_133 VDD VSS sg13g2_decap_8
XFILLER_52_497 VDD VSS sg13g2_decap_8
XFILLER_40_637 VDD VSS sg13g2_decap_8
XFILLER_20_350 VDD VSS sg13g2_decap_8
XFILLER_21_77 VDD VSS sg13g2_decap_8
XFILLER_0_700 VDD VSS sg13g2_decap_8
XFILLER_75_501 VDD VSS sg13g2_decap_8
XFILLER_87_350 VDD VSS sg13g2_decap_8
XFILLER_47_203 VDD VSS sg13g2_decap_8
XFILLER_90_504 VDD VSS sg13g2_decap_8
XFILLER_75_578 VDD VSS sg13g2_decap_8
XFILLER_63_718 VDD VSS sg13g2_decap_8
XFILLER_62_217 VDD VSS sg13g2_decap_8
XFILLER_46_63 VDD VSS sg13g2_decap_8
XFILLER_16_623 VDD VSS sg13g2_decap_8
XFILLER_28_483 VDD VSS sg13g2_decap_8
XFILLER_71_751 VDD VSS sg13g2_decap_4
XIO_CORNER_SOUTH_WEST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XFILLER_15_133 VDD VSS sg13g2_decap_8
XFILLER_43_420 VDD VSS sg13g2_decap_8
XFILLER_55_280 VDD VSS sg13g2_decap_8
XFILLER_31_637 VDD VSS sg13g2_decap_8
XFILLER_43_497 VDD VSS sg13g2_decap_8
XFILLER_62_84 VDD VSS sg13g2_decap_8
XFILLER_11_350 VDD VSS sg13g2_decap_8
XFILLER_30_147 VDD VSS sg13g2_decap_8
XFILLER_7_35 VDD VSS sg13g2_decap_8
XFILLER_7_343 VDD VSS sg13g2_decap_8
XFILLER_3_560 VDD VSS sg13g2_decap_8
XFILLER_87_70 VDD VSS sg13g2_decap_8
XFILLER_78_350 VDD VSS sg13g2_decap_8
XFILLER_38_203 VDD VSS sg13g2_decap_8
XFILLER_66_534 VDD VSS sg13g2_decap_8
XFILLER_81_504 VDD VSS sg13g2_decap_8
XFILLER_93_364 VDD VSS sg13g2_decap_8
XFILLER_54_707 VDD VSS sg13g2_decap_8
XFILLER_53_217 VDD VSS sg13g2_decap_8
XFILLER_19_483 VDD VSS sg13g2_decap_8
XFILLER_34_420 VDD VSS sg13g2_decap_8
XFILLER_46_280 VDD VSS sg13g2_decap_8
XFILLER_61_294 VDD VSS sg13g2_decap_8
XFILLER_22_637 VDD VSS sg13g2_decap_8
XFILLER_34_497 VDD VSS sg13g2_decap_8
XFILLER_21_147 VDD VSS sg13g2_decap_8
XFILLER_89_637 VDD VSS sg13g2_decap_8
XFILLER_88_147 VDD VSS sg13g2_decap_8
XFILLER_29_203 VDD VSS sg13g2_decap_8
XFILLER_69_394 VDD VSS sg13g2_decap_8
XFILLER_84_364 VDD VSS sg13g2_decap_8
XFILLER_57_567 VDD VSS sg13g2_decap_8
XFILLER_45_707 VDD VSS sg13g2_decap_8
XFILLER_72_537 VDD VSS sg13g2_decap_8
XFILLER_83_28 VDD VSS sg13g2_decap_8
XFILLER_44_217 VDD VSS sg13g2_decap_8
XFILLER_25_420 VDD VSS sg13g2_decap_8
XFILLER_37_280 VDD VSS sg13g2_decap_8
XFILLER_16_77 VDD VSS sg13g2_decap_8
XFILLER_80_581 VDD VSS sg13g2_decap_8
XFILLER_13_637 VDD VSS sg13g2_decap_8
XFILLER_40_434 VDD VSS sg13g2_decap_8
XFILLER_52_294 VDD VSS sg13g2_decap_8
XFILLER_25_497 VDD VSS sg13g2_decap_8
XFILLER_12_147 VDD VSS sg13g2_decap_8
XFILLER_32_21 VDD VSS sg13g2_decap_8
XFILLER_32_98 VDD VSS sg13g2_decap_8
X_81__9 VDD VSS _81__9/L_HI sg13g2_tiehi
XFILLER_4_357 VDD VSS sg13g2_decap_8
XFILLER_79_147 VDD VSS sg13g2_decap_8
XFILLER_0_574 VDD VSS sg13g2_decap_8
XFILLER_75_320 VDD VSS sg13g2_decap_8
XFILLER_48_567 VDD VSS sg13g2_decap_8
XFILLER_57_84 VDD VSS sg13g2_decap_8
XFILLER_36_707 VDD VSS sg13g2_decap_8
XFILLER_63_515 VDD VSS sg13g2_decap_8
XFILLER_90_301 VDD VSS sg13g2_decap_8
XFILLER_35_217 VDD VSS sg13g2_decap_8
XFILLER_16_420 VDD VSS sg13g2_decap_8
XFILLER_28_280 VDD VSS sg13g2_decap_8
XFILLER_90_378 VDD VSS sg13g2_decap_8
XFILLER_92_7 VDD VSS sg13g2_decap_8
XFILLER_31_434 VDD VSS sg13g2_decap_8
XFILLER_43_294 VDD VSS sg13g2_decap_8
XFILLER_16_497 VDD VSS sg13g2_decap_8
XFILLER_8_630 VDD VSS sg13g2_decap_8
XFILLER_7_140 VDD VSS sg13g2_decap_8
XFILLER_94_651 VDD VSS sg13g2_decap_8
XFILLER_54_504 VDD VSS sg13g2_decap_8
XFILLER_14_0 VDD VSS sg13g2_decap_8
XFILLER_27_707 VDD VSS sg13g2_decap_8
XFILLER_39_567 VDD VSS sg13g2_decap_8
XFILLER_93_161 VDD VSS sg13g2_decap_8
XFILLER_81_301 VDD VSS sg13g2_decap_8
XFILLER_66_364 VDD VSS sg13g2_decap_8
XFILLER_26_217 VDD VSS sg13g2_decap_8
XFILLER_19_280 VDD VSS sg13g2_decap_8
XFILLER_81_378 VDD VSS sg13g2_decap_8
XFILLER_62_581 VDD VSS sg13g2_decap_8
XFILLER_50_721 VDD VSS sg13g2_decap_8
XFILLER_22_434 VDD VSS sg13g2_decap_8
XFILLER_34_294 VDD VSS sg13g2_decap_8
XFILLER_78_28 VDD VSS sg13g2_decap_8
XFILLER_89_434 VDD VSS sg13g2_decap_8
XFILLER_77_618 VDD VSS sg13g2_decap_8
XFILLER_85_651 VDD VSS sg13g2_decap_8
XFILLER_94_49 VDD VSS sg13g2_decap_8
XFILLER_18_707 VDD VSS sg13g2_decap_8
XFILLER_84_161 VDD VSS sg13g2_decap_8
XFILLER_72_301 VDD VSS sg13g2_fill_1
XFILLER_27_21 VDD VSS sg13g2_decap_8
XFILLER_17_217 VDD VSS sg13g2_decap_8
XFILLER_57_364 VDD VSS sg13g2_decap_8
XFILLER_45_504 VDD VSS sg13g2_decap_8
XFILLER_72_367 VDD VSS sg13g2_decap_8
XFILLER_60_518 VDD VSS sg13g2_decap_8
XFILLER_27_98 VDD VSS sg13g2_decap_8
XFILLER_53_581 VDD VSS sg13g2_decap_8
XFILLER_13_434 VDD VSS sg13g2_decap_8
XFILLER_25_294 VDD VSS sg13g2_decap_8
XFILLER_41_721 VDD VSS sg13g2_decap_8
XFILLER_43_42 VDD VSS sg13g2_decap_8
XFILLER_40_231 VDD VSS sg13g2_decap_8
XFILLER_9_427 VDD VSS sg13g2_decap_8
XFILLER_5_644 VDD VSS sg13g2_decap_8
XFILLER_4_154 VDD VSS sg13g2_decap_8
XFILLER_4_14 VDD VSS sg13g2_decap_8
XFILLER_68_629 VDD VSS sg13g2_decap_8
XFILLER_95_448 VDD VSS sg13g2_decap_8
XFILLER_0_371 VDD VSS sg13g2_decap_8
XFILLER_75_172 VDD VSS sg13g2_decap_8
XFILLER_63_301 VDD VSS sg13g2_decap_8
XFILLER_48_364 VDD VSS sg13g2_decap_8
XFILLER_36_504 VDD VSS sg13g2_decap_8
XFILLER_91_665 VDD VSS sg13g2_decap_8
XFILLER_63_378 VDD VSS sg13g2_decap_8
XFILLER_51_518 VDD VSS sg13g2_decap_8
XFILLER_90_175 VDD VSS sg13g2_decap_8
XFILLER_32_721 VDD VSS sg13g2_decap_8
XFILLER_44_581 VDD VSS sg13g2_decap_8
XFILLER_16_294 VDD VSS sg13g2_decap_8
XFILLER_31_231 VDD VSS sg13g2_decap_8
XFILLER_86_448 VDD VSS sg13g2_decap_8
XFILLER_67_695 VDD VSS sg13g2_decap_8
XFILLER_66_161 VDD VSS sg13g2_decap_8
XFILLER_39_364 VDD VSS sg13g2_decap_8
XFILLER_54_301 VDD VSS sg13g2_decap_8
XFILLER_27_504 VDD VSS sg13g2_decap_8
XFILLER_82_665 VDD VSS sg13g2_decap_8
XFILLER_54_378 VDD VSS sg13g2_decap_8
XFILLER_42_518 VDD VSS sg13g2_decap_8
XFILLER_81_175 VDD VSS sg13g2_decap_8
XFILLER_23_721 VDD VSS sg13g2_decap_8
XFILLER_35_581 VDD VSS sg13g2_decap_8
XFILLER_22_231 VDD VSS sg13g2_decap_8
XFILLER_50_595 VDD VSS sg13g2_decap_8
XFILLER_10_448 VDD VSS sg13g2_decap_8
XFILLER_13_56 VDD VSS sg13g2_decap_8
XFILLER_89_49 VDD VSS sg13g2_decap_8
XFILLER_89_231 VDD VSS sg13g2_decap_8
XFILLER_2_658 VDD VSS sg13g2_decap_8
XFILLER_1_168 VDD VSS sg13g2_decap_8
XFILLER_58_651 VDD VSS sg13g2_decap_8
XFILLER_38_42 VDD VSS sg13g2_decap_8
XFILLER_45_301 VDD VSS sg13g2_decap_8
XFILLER_57_161 VDD VSS sg13g2_decap_8
XFILLER_18_504 VDD VSS sg13g2_decap_8
XFILLER_73_632 VDD VSS sg13g2_decap_8
XFILLER_45_378 VDD VSS sg13g2_decap_8
XFILLER_33_518 VDD VSS sg13g2_decap_8
XFILLER_72_175 VDD VSS sg13g2_decap_8
XFILLER_54_63 VDD VSS sg13g2_decap_8
XFILLER_60_315 VDD VSS sg13g2_decap_8
XFILLER_14_721 VDD VSS sg13g2_decap_8
XFILLER_13_231 VDD VSS sg13g2_decap_8
XFILLER_9_224 VDD VSS sg13g2_decap_8
XFILLER_41_595 VDD VSS sg13g2_decap_8
XFILLER_70_84 VDD VSS sg13g2_decap_8
XFILLER_5_441 VDD VSS sg13g2_decap_8
XFILLER_55_7 VDD VSS sg13g2_decap_8
XFILLER_68_426 VDD VSS sg13g2_decap_8
XFILLER_95_245 VDD VSS sg13g2_decap_8
XFILLER_49_651 VDD VSS sg13g2_decap_8
XFILLER_95_70 VDD VSS sg13g2_decap_8
XFILLER_36_301 VDD VSS sg13g2_decap_8
XFILLER_48_161 VDD VSS sg13g2_decap_8
XFILLER_64_665 VDD VSS sg13g2_decap_8
XFILLER_91_462 VDD VSS sg13g2_decap_8
XFILLER_36_378 VDD VSS sg13g2_decap_8
XFILLER_24_518 VDD VSS sg13g2_decap_8
XFILLER_63_175 VDD VSS sg13g2_decap_8
XFILLER_51_315 VDD VSS sg13g2_decap_8
XFILLER_17_581 VDD VSS sg13g2_decap_8
XFILLER_81_0 VDD VSS sg13g2_decap_8
XFILLER_20_735 VDD VSS sg13g2_decap_8
XFILLER_32_595 VDD VSS sg13g2_decap_8
XFILLER_87_735 VDD VSS sg13g2_decap_8
XFILLER_86_245 VDD VSS sg13g2_decap_8
XFILLER_59_448 VDD VSS sg13g2_decap_8
XFILLER_27_301 VDD VSS sg13g2_decap_8
XFILLER_39_161 VDD VSS sg13g2_decap_8
XFILLER_67_492 VDD VSS sg13g2_decap_8
XFILLER_82_462 VDD VSS sg13g2_decap_8
XFILLER_55_665 VDD VSS sg13g2_decap_8
XFILLER_27_378 VDD VSS sg13g2_decap_8
XFILLER_15_518 VDD VSS sg13g2_decap_8
XFILLER_70_624 VDD VSS sg13g2_decap_8
XFILLER_91_28 VDD VSS sg13g2_decap_8
XFILLER_42_315 VDD VSS sg13g2_decap_8
XFILLER_54_175 VDD VSS sg13g2_decap_8
XFILLER_11_735 VDD VSS sg13g2_decap_8
XFILLER_24_77 VDD VSS sg13g2_decap_8
XFILLER_50_392 VDD VSS sg13g2_decap_8
XFILLER_23_595 VDD VSS sg13g2_decap_8
XFILLER_7_728 VDD VSS sg13g2_decap_8
XFILLER_10_245 VDD VSS sg13g2_decap_8
XFILLER_6_238 VDD VSS sg13g2_decap_8
XFILLER_40_21 VDD VSS sg13g2_decap_8
XFILLER_40_98 VDD VSS sg13g2_decap_8
XFILLER_2_455 VDD VSS sg13g2_decap_8
XFILLER_78_735 VDD VSS sg13g2_decap_8
XFILLER_49_63 VDD VSS sg13g2_decap_8
XFILLER_77_267 VDD VSS sg13g2_decap_8
XFILLER_18_301 VDD VSS sg13g2_decap_8
XFILLER_93_749 VDD VSS sg13g2_decap_8
XFILLER_92_259 VDD VSS sg13g2_decap_8
XFILLER_73_451 VDD VSS sg13g2_fill_1
XFILLER_65_84 VDD VSS sg13g2_decap_8
XFILLER_61_602 VDD VSS sg13g2_decap_8
XFILLER_46_665 VDD VSS sg13g2_decap_8
XFILLER_18_378 VDD VSS sg13g2_decap_8
XFILLER_33_315 VDD VSS sg13g2_decap_8
XFILLER_45_175 VDD VSS sg13g2_decap_8
XFILLER_60_112 VDD VSS sg13g2_decap_8
XFILLER_61_679 VDD VSS sg13g2_decap_8
XFILLER_60_189 VDD VSS sg13g2_decap_8
XFILLER_41_392 VDD VSS sg13g2_decap_8
XFILLER_14_595 VDD VSS sg13g2_decap_8
XFILLER_69_713 VDD VSS sg13g2_decap_8
XFILLER_68_223 VDD VSS sg13g2_decap_8
XFILLER_84_749 VDD VSS sg13g2_decap_8
XFILLER_83_259 VDD VSS sg13g2_decap_8
X_78_ _78__8/L_HI VSS VDD _78_/D _78_/Q _79_/CLK sg13g2_dfrbpq_1
XFILLER_64_462 VDD VSS sg13g2_decap_8
XFILLER_52_602 VDD VSS sg13g2_decap_8
XFILLER_37_665 VDD VSS sg13g2_decap_8
XFILLER_24_315 VDD VSS sg13g2_decap_8
XFILLER_36_175 VDD VSS sg13g2_decap_8
XFILLER_51_112 VDD VSS sg13g2_decap_8
XFILLER_52_679 VDD VSS sg13g2_decap_8
XFILLER_51_189 VDD VSS sg13g2_decap_8
XFILLER_32_392 VDD VSS sg13g2_decap_8
XFILLER_20_532 VDD VSS sg13g2_decap_8
XFILLER_10_35 VDD VSS sg13g2_decap_8
XFILLER_86_28 VDD VSS sg13g2_decap_8
XFILLER_87_532 VDD VSS sg13g2_decap_8
XFILLER_59_245 VDD VSS sg13g2_decap_8
XFILLER_19_77 VDD VSS sg13g2_decap_8
XFILLER_55_462 VDD VSS sg13g2_decap_8
XFILLER_28_665 VDD VSS sg13g2_decap_8
XFILLER_43_602 VDD VSS sg13g2_decap_8
XFILLER_35_21 VDD VSS sg13g2_decap_8
XFILLER_15_315 VDD VSS sg13g2_decap_8
XFILLER_27_175 VDD VSS sg13g2_decap_8
XFILLER_42_112 VDD VSS sg13g2_decap_8
XFILLER_70_432 VDD VSS sg13g2_decap_8
XFILLER_35_98 VDD VSS sg13g2_decap_8
XFILLER_43_679 VDD VSS sg13g2_decap_8
XFILLER_70_498 VDD VSS sg13g2_decap_8
XFILLER_11_532 VDD VSS sg13g2_decap_8
XFILLER_23_392 VDD VSS sg13g2_decap_8
XFILLER_30_329 VDD VSS sg13g2_decap_8
XFILLER_42_189 VDD VSS sg13g2_decap_8
XFILLER_51_42 VDD VSS sg13g2_decap_8
XFILLER_7_525 VDD VSS sg13g2_decap_8
XFILLER_3_742 VDD VSS sg13g2_decap_8
XFILLER_2_252 VDD VSS sg13g2_decap_8
XFILLER_78_532 VDD VSS sg13g2_decap_8
XFILLER_66_716 VDD VSS sg13g2_decap_8
XFILLER_93_546 VDD VSS sg13g2_decap_8
XFILLER_18_7 VDD VSS sg13g2_decap_8
XFILLER_65_259 VDD VSS sg13g2_decap_8
XFILLER_19_665 VDD VSS sg13g2_decap_8
XFILLER_18_175 VDD VSS sg13g2_decap_8
XFILLER_46_462 VDD VSS sg13g2_decap_8
XFILLER_34_602 VDD VSS sg13g2_decap_8
XFILLER_33_112 VDD VSS sg13g2_decap_8
XFILLER_61_476 VDD VSS sg13g2_decap_8
XFILLER_34_679 VDD VSS sg13g2_decap_8
XFILLER_14_392 VDD VSS sg13g2_decap_8
XFILLER_21_329 VDD VSS sg13g2_decap_8
XFILLER_33_189 VDD VSS sg13g2_decap_8
XFILLER_44_0 VDD VSS sg13g2_decap_8
XFILLER_69_510 VDD VSS sg13g2_decap_8
XFILLER_88_329 VDD VSS sg13g2_decap_8
XFILLER_69_587 VDD VSS sg13g2_decap_8
XFILLER_84_546 VDD VSS sg13g2_decap_8
XFILLER_57_749 VDD VSS sg13g2_decap_8
XFILLER_72_719 VDD VSS sg13g2_decap_8
XFILLER_2_91 VDD VSS sg13g2_decap_8
XFILLER_56_259 VDD VSS sg13g2_decap_8
XFILLER_37_462 VDD VSS sg13g2_decap_8
XFILLER_25_602 VDD VSS sg13g2_decap_8
XFILLER_24_112 VDD VSS sg13g2_decap_8
XFILLER_52_476 VDD VSS sg13g2_decap_8
XFILLER_25_679 VDD VSS sg13g2_decap_8
XFILLER_40_616 VDD VSS sg13g2_decap_8
XFILLER_12_329 VDD VSS sg13g2_decap_8
XFILLER_24_189 VDD VSS sg13g2_decap_8
XFILLER_4_539 VDD VSS sg13g2_decap_8
XFILLER_21_56 VDD VSS sg13g2_decap_8
XFILLER_79_329 VDD VSS sg13g2_decap_8
XFILLER_48_749 VDD VSS sg13g2_decap_8
XFILLER_75_557 VDD VSS sg13g2_decap_8
XFILLER_46_42 VDD VSS sg13g2_decap_8
XFILLER_47_259 VDD VSS sg13g2_decap_8
XFILLER_28_462 VDD VSS sg13g2_decap_8
XFILLER_16_602 VDD VSS sg13g2_decap_8
XFILLER_71_730 VDD VSS sg13g2_decap_8
XFILLER_15_112 VDD VSS sg13g2_decap_8
XFILLER_43_476 VDD VSS sg13g2_decap_8
XFILLER_16_679 VDD VSS sg13g2_decap_8
XFILLER_31_616 VDD VSS sg13g2_decap_8
XFILLER_70_284 VDD VSS sg13g2_decap_8
XFILLER_62_63 VDD VSS sg13g2_decap_8
XFILLER_15_189 VDD VSS sg13g2_decap_8
XFILLER_30_126 VDD VSS sg13g2_decap_8
XFILLER_7_322 VDD VSS sg13g2_decap_8
XFILLER_7_14 VDD VSS sg13g2_decap_8
XFILLER_7_399 VDD VSS sg13g2_decap_8
XFILLER_66_513 VDD VSS sg13g2_decap_8
XFILLER_39_749 VDD VSS sg13g2_decap_8
XFILLER_93_343 VDD VSS sg13g2_decap_8
XFILLER_38_259 VDD VSS sg13g2_decap_8
XFILLER_19_462 VDD VSS sg13g2_decap_8
XFILLER_34_476 VDD VSS sg13g2_decap_8
XFILLER_22_616 VDD VSS sg13g2_decap_8
XFILLER_21_126 VDD VSS sg13g2_decap_8
XFILLER_61_273 VDD VSS sg13g2_decap_8
XFILLER_30_693 VDD VSS sg13g2_decap_8
XFILLER_89_616 VDD VSS sg13g2_decap_8
XFILLER_88_126 VDD VSS sg13g2_decap_8
XFILLER_69_373 VDD VSS sg13g2_decap_8
XFILLER_84_343 VDD VSS sg13g2_decap_8
XFILLER_57_546 VDD VSS sg13g2_decap_8
XFILLER_29_259 VDD VSS sg13g2_decap_8
XFILLER_72_516 VDD VSS sg13g2_decap_8
XFILLER_80_560 VDD VSS sg13g2_decap_8
XFILLER_13_616 VDD VSS sg13g2_decap_8
XFILLER_16_56 VDD VSS sg13g2_decap_8
XFILLER_25_476 VDD VSS sg13g2_decap_8
XFILLER_12_126 VDD VSS sg13g2_decap_8
XFILLER_40_413 VDD VSS sg13g2_decap_8
XFILLER_52_273 VDD VSS sg13g2_decap_8
XFILLER_9_609 VDD VSS sg13g2_decap_8
XFILLER_8_119 VDD VSS sg13g2_decap_8
XFILLER_32_77 VDD VSS sg13g2_decap_8
XFILLER_21_693 VDD VSS sg13g2_decap_8
XFILLER_4_336 VDD VSS sg13g2_decap_8
XFILLER_79_126 VDD VSS sg13g2_decap_8
XFILLER_0_553 VDD VSS sg13g2_decap_8
XFILLER_88_693 VDD VSS sg13g2_decap_8
XFILLER_48_546 VDD VSS sg13g2_decap_8
XFILLER_57_63 VDD VSS sg13g2_decap_8
XFILLER_90_357 VDD VSS sg13g2_decap_8
XFILLER_16_476 VDD VSS sg13g2_decap_8
XFILLER_73_84 VDD VSS sg13g2_decap_8
XFILLER_31_413 VDD VSS sg13g2_decap_8
XFILLER_43_273 VDD VSS sg13g2_decap_8
XFILLER_85_7 VDD VSS sg13g2_decap_8
XFILLER_12_693 VDD VSS sg13g2_decap_8
XFILLER_8_686 VDD VSS sg13g2_decap_8
XFILLER_7_196 VDD VSS sg13g2_decap_8
XFILLER_94_630 VDD VSS sg13g2_decap_8
XFILLER_79_693 VDD VSS sg13g2_decap_8
XFILLER_93_140 VDD VSS sg13g2_decap_8
XFILLER_66_343 VDD VSS sg13g2_decap_8
XFILLER_39_546 VDD VSS sg13g2_decap_8
XFILLER_62_560 VDD VSS sg13g2_decap_8
XFILLER_81_357 VDD VSS sg13g2_decap_8
XFILLER_50_700 VDD VSS sg13g2_decap_8
XFILLER_22_413 VDD VSS sg13g2_decap_8
XFILLER_34_273 VDD VSS sg13g2_decap_8
XFILLER_30_490 VDD VSS sg13g2_decap_8
XFILLER_89_413 VDD VSS sg13g2_decap_8
XFILLER_85_630 VDD VSS sg13g2_decap_8
XFILLER_94_28 VDD VSS sg13g2_decap_8
XFILLER_57_343 VDD VSS sg13g2_decap_8
XFILLER_84_140 VDD VSS sg13g2_decap_8
XFILLER_27_77 VDD VSS sg13g2_decap_8
XFILLER_26_741 VDD VSS sg13g2_decap_8
XFILLER_53_560 VDD VSS sg13g2_decap_8
XFILLER_41_700 VDD VSS sg13g2_decap_8
XFILLER_13_413 VDD VSS sg13g2_decap_8
XFILLER_43_21 VDD VSS sg13g2_decap_8
XFILLER_25_273 VDD VSS sg13g2_decap_8
XFILLER_40_210 VDD VSS sg13g2_decap_8
XFILLER_9_406 VDD VSS sg13g2_decap_8
XFILLER_43_98 VDD VSS sg13g2_decap_8
XFILLER_40_287 VDD VSS sg13g2_decap_8
XFILLER_21_490 VDD VSS sg13g2_decap_8
XFILLER_5_623 VDD VSS sg13g2_decap_8
XFILLER_4_133 VDD VSS sg13g2_decap_8
XFILLER_68_608 VDD VSS sg13g2_decap_8
XFILLER_95_427 VDD VSS sg13g2_decap_8
XFILLER_68_84 VDD VSS sg13g2_decap_8
XFILLER_0_350 VDD VSS sg13g2_decap_8
XFILLER_88_490 VDD VSS sg13g2_decap_8
XFILLER_48_343 VDD VSS sg13g2_decap_8
XFILLER_76_685 VDD VSS sg13g2_decap_8
XFILLER_75_151 VDD VSS sg13g2_decap_8
XFILLER_91_644 VDD VSS sg13g2_decap_8
XFILLER_90_154 VDD VSS sg13g2_decap_8
XFILLER_63_357 VDD VSS sg13g2_decap_8
XFILLER_32_700 VDD VSS sg13g2_decap_8
XFILLER_44_560 VDD VSS sg13g2_decap_8
XFILLER_16_273 VDD VSS sg13g2_decap_8
XFILLER_31_210 VDD VSS sg13g2_decap_8
XFILLER_12_490 VDD VSS sg13g2_decap_8
XFILLER_31_287 VDD VSS sg13g2_decap_8
XFILLER_8_483 VDD VSS sg13g2_decap_8
XFILLER_86_427 VDD VSS sg13g2_decap_8
XFILLER_79_490 VDD VSS sg13g2_decap_8
XFILLER_39_343 VDD VSS sg13g2_decap_8
XFILLER_67_674 VDD VSS sg13g2_decap_8
XFILLER_66_140 VDD VSS sg13g2_decap_8
XFILLER_82_644 VDD VSS sg13g2_decap_8
XFILLER_81_154 VDD VSS sg13g2_decap_8
XFILLER_54_357 VDD VSS sg13g2_decap_8
XFILLER_23_700 VDD VSS sg13g2_decap_8
XFILLER_22_210 VDD VSS sg13g2_decap_8
XFILLER_35_560 VDD VSS sg13g2_decap_8
XFILLER_50_574 VDD VSS sg13g2_decap_8
XFILLER_10_427 VDD VSS sg13g2_decap_8
XFILLER_13_35 VDD VSS sg13g2_decap_8
XFILLER_22_287 VDD VSS sg13g2_decap_8
XFILLER_89_28 VDD VSS sg13g2_decap_8
XFILLER_89_210 VDD VSS sg13g2_decap_8
XFILLER_2_637 VDD VSS sg13g2_decap_8
XFILLER_1_147 VDD VSS sg13g2_decap_8
XFILLER_89_287 VDD VSS sg13g2_decap_8
XFILLER_38_21 VDD VSS sg13g2_decap_8
XFILLER_77_449 VDD VSS sg13g2_decap_8
XFILLER_58_630 VDD VSS sg13g2_decap_8
XFILLER_73_611 VDD VSS sg13g2_decap_8
XFILLER_57_140 VDD VSS sg13g2_decap_8
XFILLER_38_98 VDD VSS sg13g2_decap_8
XFILLER_73_688 VDD VSS sg13g2_decap_8
XFILLER_72_154 VDD VSS sg13g2_decap_8
XFILLER_45_357 VDD VSS sg13g2_decap_8
XFILLER_54_42 VDD VSS sg13g2_decap_8
XFILLER_14_700 VDD VSS sg13g2_decap_8
XFILLER_13_210 VDD VSS sg13g2_decap_8
XFILLER_9_203 VDD VSS sg13g2_decap_8
XFILLER_41_574 VDD VSS sg13g2_decap_8
XFILLER_13_287 VDD VSS sg13g2_decap_8
XFILLER_70_63 VDD VSS sg13g2_decap_8
XFILLER_5_420 VDD VSS sg13g2_decap_8
XFILLER_5_497 VDD VSS sg13g2_decap_8
XFILLER_48_7 VDD VSS sg13g2_decap_8
XFILLER_68_405 VDD VSS sg13g2_decap_8
XFILLER_95_224 VDD VSS sg13g2_decap_8
XFILLER_49_630 VDD VSS sg13g2_decap_8
XFILLER_48_140 VDD VSS sg13g2_decap_8
XFILLER_64_644 VDD VSS sg13g2_decap_8
XFILLER_76_482 VDD VSS sg13g2_decap_8
XFILLER_91_441 VDD VSS sg13g2_decap_8
XFILLER_63_154 VDD VSS sg13g2_decap_8
XFILLER_36_357 VDD VSS sg13g2_decap_8
XFILLER_17_560 VDD VSS sg13g2_decap_8
XFILLER_20_714 VDD VSS sg13g2_decap_8
XFILLER_32_574 VDD VSS sg13g2_decap_8
XFILLER_74_0 VDD VSS sg13g2_decap_8
XFILLER_8_280 VDD VSS sg13g2_decap_8
XFILLER_5_91 VDD VSS sg13g2_decap_8
XFILLER_87_714 VDD VSS sg13g2_decap_8
XFILLER_59_427 VDD VSS sg13g2_decap_8
XFILLER_86_224 VDD VSS sg13g2_decap_8
XFILLER_39_140 VDD VSS sg13g2_decap_8
XFILLER_67_471 VDD VSS sg13g2_decap_8
XFILLER_55_644 VDD VSS sg13g2_decap_8
XFILLER_70_603 VDD VSS sg13g2_decap_8
XFILLER_82_441 VDD VSS sg13g2_decap_8
XFILLER_27_357 VDD VSS sg13g2_decap_8
XFILLER_54_154 VDD VSS sg13g2_decap_8
XFILLER_11_714 VDD VSS sg13g2_decap_8
XFILLER_24_56 VDD VSS sg13g2_decap_8
XFILLER_23_574 VDD VSS sg13g2_decap_8
XFILLER_7_707 VDD VSS sg13g2_decap_8
XFILLER_10_224 VDD VSS sg13g2_decap_8
XFILLER_50_371 VDD VSS sg13g2_decap_8
XFILLER_6_217 VDD VSS sg13g2_decap_8
XFILLER_40_77 VDD VSS sg13g2_decap_8
XFILLER_2_434 VDD VSS sg13g2_decap_8
XFILLER_78_714 VDD VSS sg13g2_decap_8
XFILLER_49_42 VDD VSS sg13g2_decap_8
XFILLER_77_224 VDD VSS sg13g2_fill_2
XFILLER_93_728 VDD VSS sg13g2_decap_8
XFILLER_92_238 VDD VSS sg13g2_decap_8
XFILLER_46_644 VDD VSS sg13g2_decap_8
XFILLER_1_49 VDD VSS sg13g2_decap_8
XFILLER_65_63 VDD VSS sg13g2_decap_8
XFILLER_18_357 VDD VSS sg13g2_decap_8
XFILLER_45_154 VDD VSS sg13g2_decap_8
XFILLER_73_485 VDD VSS sg13g2_decap_8
XFILLER_61_658 VDD VSS sg13g2_decap_8
XFILLER_60_168 VDD VSS sg13g2_decap_8
XFILLER_14_574 VDD VSS sg13g2_decap_8
XFILLER_81_84 VDD VSS sg13g2_decap_8
XFILLER_41_371 VDD VSS sg13g2_decap_8
XFILLER_5_294 VDD VSS sg13g2_decap_8
XFILLER_68_202 VDD VSS sg13g2_decap_8
XFILLER_84_728 VDD VSS sg13g2_decap_8
XFILLER_68_279 VDD VSS sg13g2_decap_8
XFILLER_83_238 VDD VSS sg13g2_decap_8
X_77_ _77__10/L_HI VSS VDD _77_/D _77_/Q _79_/CLK sg13g2_dfrbpq_1
XFILLER_64_441 VDD VSS sg13g2_decap_8
XFILLER_37_644 VDD VSS sg13g2_decap_8
XFILLER_36_154 VDD VSS sg13g2_decap_8
XFILLER_52_658 VDD VSS sg13g2_decap_8
XFILLER_51_168 VDD VSS sg13g2_decap_8
XFILLER_32_371 VDD VSS sg13g2_decap_8
XFILLER_20_511 VDD VSS sg13g2_decap_8
XFILLER_20_588 VDD VSS sg13g2_decap_8
XFILLER_10_14 VDD VSS sg13g2_decap_8
XFILLER_87_511 VDD VSS sg13g2_decap_8
XFILLER_59_224 VDD VSS sg13g2_decap_8
XFILLER_87_588 VDD VSS sg13g2_decap_8
XFILLER_19_56 VDD VSS sg13g2_decap_8
XFILLER_75_739 VDD VSS sg13g2_decap_8
XFILLER_55_441 VDD VSS sg13g2_decap_8
XFILLER_28_644 VDD VSS sg13g2_decap_8
XFILLER_70_411 VDD VSS sg13g2_decap_8
XFILLER_27_154 VDD VSS sg13g2_decap_8
XFILLER_43_658 VDD VSS sg13g2_decap_8
XFILLER_70_455 VDD VSS sg13g2_fill_1
XFILLER_35_77 VDD VSS sg13g2_decap_8
XFILLER_30_308 VDD VSS sg13g2_decap_8
XFILLER_42_168 VDD VSS sg13g2_decap_8
XFILLER_11_511 VDD VSS sg13g2_decap_8
XFILLER_51_21 VDD VSS sg13g2_decap_8
XFILLER_23_371 VDD VSS sg13g2_decap_8
XFILLER_7_504 VDD VSS sg13g2_decap_8
XFILLER_11_588 VDD VSS sg13g2_decap_8
XFILLER_51_98 VDD VSS sg13g2_decap_8
XFILLER_3_721 VDD VSS sg13g2_decap_8
XFILLER_4_0 VDD VSS sg13g2_decap_8
XFILLER_2_231 VDD VSS sg13g2_decap_8
XFILLER_78_511 VDD VSS sg13g2_decap_8
XFILLER_78_588 VDD VSS sg13g2_decap_8
XFILLER_93_525 VDD VSS sg13g2_decap_8
XFILLER_65_238 VDD VSS sg13g2_decap_8
XFILLER_76_84 VDD VSS sg13g2_decap_8
XFILLER_46_441 VDD VSS sg13g2_decap_8
XFILLER_19_644 VDD VSS sg13g2_decap_8
XFILLER_18_154 VDD VSS sg13g2_decap_8
XFILLER_34_658 VDD VSS sg13g2_decap_8
XFILLER_21_308 VDD VSS sg13g2_decap_8
XFILLER_33_168 VDD VSS sg13g2_decap_8
XFILLER_61_455 VDD VSS sg13g2_decap_8
XFILLER_14_371 VDD VSS sg13g2_decap_8
XFILLER_6_581 VDD VSS sg13g2_decap_8
XFILLER_88_308 VDD VSS sg13g2_decap_8
XFILLER_37_0 VDD VSS sg13g2_decap_8
XFILLER_69_566 VDD VSS sg13g2_decap_8
XFILLER_57_728 VDD VSS sg13g2_decap_8
XFILLER_84_525 VDD VSS sg13g2_decap_8
XFILLER_2_70 VDD VSS sg13g2_decap_8
XFILLER_56_238 VDD VSS sg13g2_decap_8
XFILLER_37_441 VDD VSS sg13g2_decap_8
XFILLER_80_742 VDD VSS sg13g2_decap_8
XFILLER_25_658 VDD VSS sg13g2_decap_8
XFILLER_12_308 VDD VSS sg13g2_decap_8
XFILLER_24_168 VDD VSS sg13g2_decap_8
XFILLER_52_455 VDD VSS sg13g2_decap_8
XFILLER_21_35 VDD VSS sg13g2_decap_8
XFILLER_20_385 VDD VSS sg13g2_decap_8
XFILLER_4_518 VDD VSS sg13g2_decap_8
XFILLER_79_308 VDD VSS sg13g2_decap_8
XFILLER_0_735 VDD VSS sg13g2_decap_8
XFILLER_48_728 VDD VSS sg13g2_decap_8
XFILLER_75_536 VDD VSS sg13g2_decap_8
XFILLER_87_385 VDD VSS sg13g2_decap_8
XFILLER_46_21 VDD VSS sg13g2_decap_8
XFILLER_28_441 VDD VSS sg13g2_decap_8
XFILLER_47_238 VDD VSS sg13g2_decap_8
XFILLER_90_539 VDD VSS sg13g2_decap_8
XFILLER_46_98 VDD VSS sg13g2_decap_8
XFILLER_16_658 VDD VSS sg13g2_decap_8
XFILLER_70_263 VDD VSS sg13g2_decap_8
XFILLER_15_168 VDD VSS sg13g2_decap_8
XFILLER_43_455 VDD VSS sg13g2_decap_8
XFILLER_62_42 VDD VSS sg13g2_decap_8
XFILLER_30_105 VDD VSS sg13g2_decap_8
XFILLER_7_301 VDD VSS sg13g2_decap_8
XFILLER_11_385 VDD VSS sg13g2_decap_8
XFILLER_7_378 VDD VSS sg13g2_decap_8
XFILLER_3_595 VDD VSS sg13g2_decap_8
XFILLER_30_7 VDD VSS sg13g2_decap_8
XFILLER_93_322 VDD VSS sg13g2_decap_8
XFILLER_78_385 VDD VSS sg13g2_decap_8
XFILLER_39_728 VDD VSS sg13g2_decap_8
XFILLER_66_569 VDD VSS sg13g2_decap_8
XFILLER_19_441 VDD VSS sg13g2_decap_8
XFILLER_38_238 VDD VSS sg13g2_decap_8
XFILLER_81_539 VDD VSS sg13g2_decap_8
XFILLER_62_742 VDD VSS sg13g2_decap_8
XFILLER_93_399 VDD VSS sg13g2_decap_8
XFILLER_34_455 VDD VSS sg13g2_decap_8
XFILLER_61_252 VDD VSS sg13g2_decap_8
XFILLER_21_105 VDD VSS sg13g2_decap_8
XFILLER_30_672 VDD VSS sg13g2_decap_8
XFILLER_88_105 VDD VSS sg13g2_decap_8
XFILLER_69_352 VDD VSS sg13g2_decap_8
XFILLER_84_322 VDD VSS sg13g2_decap_8
XFILLER_57_525 VDD VSS sg13g2_decap_8
XFILLER_29_238 VDD VSS sg13g2_decap_8
XFILLER_65_591 VDD VSS sg13g2_decap_8
XFILLER_84_399 VDD VSS sg13g2_decap_8
XFILLER_53_742 VDD VSS sg13g2_decap_8
XFILLER_16_35 VDD VSS sg13g2_decap_8
XFILLER_25_455 VDD VSS sg13g2_decap_8
XFILLER_52_252 VDD VSS sg13g2_decap_8
XFILLER_12_105 VDD VSS sg13g2_decap_8
XFILLER_40_469 VDD VSS sg13g2_decap_8
XFILLER_32_56 VDD VSS sg13g2_decap_8
XFILLER_21_672 VDD VSS sg13g2_decap_8
XFILLER_20_182 VDD VSS sg13g2_decap_8
XFILLER_4_315 VDD VSS sg13g2_decap_8
XFILLER_79_105 VDD VSS sg13g2_decap_8
XFILLER_95_609 VDD VSS sg13g2_decap_8
XFILLER_0_532 VDD VSS sg13g2_decap_8
XFILLER_88_672 VDD VSS sg13g2_decap_8
XFILLER_94_119 VDD VSS sg13g2_decap_8
XFILLER_48_525 VDD VSS sg13g2_decap_8
XFILLER_57_42 VDD VSS sg13g2_decap_8
XFILLER_87_182 VDD VSS sg13g2_decap_8
XFILLER_75_355 VDD VSS sg13g2_fill_1
XFILLER_75_388 VDD VSS sg13g2_decap_8
XFILLER_90_336 VDD VSS sg13g2_decap_8
XFILLER_44_742 VDD VSS sg13g2_decap_8
XFILLER_73_63 VDD VSS sg13g2_decap_8
XFILLER_16_455 VDD VSS sg13g2_decap_8
XFILLER_43_252 VDD VSS sg13g2_decap_8
XFILLER_71_583 VDD VSS sg13g2_decap_8
XFILLER_31_469 VDD VSS sg13g2_decap_8
XFILLER_12_672 VDD VSS sg13g2_decap_8
XFILLER_78_7 VDD VSS sg13g2_decap_8
XFILLER_8_665 VDD VSS sg13g2_decap_8
XFILLER_11_182 VDD VSS sg13g2_decap_8
XFILLER_7_175 VDD VSS sg13g2_decap_8
XFILLER_86_609 VDD VSS sg13g2_decap_8
XFILLER_3_392 VDD VSS sg13g2_decap_8
XFILLER_79_672 VDD VSS sg13g2_decap_8
XFILLER_85_119 VDD VSS sg13g2_decap_8
XFILLER_39_525 VDD VSS sg13g2_decap_8
XFILLER_78_182 VDD VSS sg13g2_decap_8
XFILLER_66_322 VDD VSS sg13g2_decap_8
XFILLER_94_686 VDD VSS sg13g2_decap_8
XIO_BOND_outputs\[1\].output_pad output_PAD[1] bondpad_70x70_novias
XFILLER_93_196 VDD VSS sg13g2_decap_8
XFILLER_81_336 VDD VSS sg13g2_decap_8
XFILLER_66_399 VDD VSS sg13g2_decap_8
XFILLER_54_539 VDD VSS sg13g2_decap_8
XFILLER_35_742 VDD VSS sg13g2_decap_8
XFILLER_34_252 VDD VSS sg13g2_decap_8
XFILLER_50_756 VDD VSS sg13g2_fill_1
XFILLER_10_609 VDD VSS sg13g2_decap_8
XFILLER_22_469 VDD VSS sg13g2_decap_8
XFILLER_8_91 VDD VSS sg13g2_decap_8
XFILLER_1_329 VDD VSS sg13g2_decap_8
XFILLER_89_469 VDD VSS sg13g2_decap_8
XFILLER_76_119 VDD VSS sg13g2_decap_8
XFILLER_69_182 VDD VSS sg13g2_decap_8
XFILLER_57_322 VDD VSS sg13g2_decap_8
XFILLER_85_686 VDD VSS sg13g2_decap_8
XFILLER_84_196 VDD VSS sg13g2_decap_8
XFILLER_72_325 VDD VSS sg13g2_decap_8
XFILLER_72_336 VDD VSS sg13g2_fill_1
XFILLER_27_56 VDD VSS sg13g2_decap_8
XFILLER_57_399 VDD VSS sg13g2_decap_8
XFILLER_26_720 VDD VSS sg13g2_decap_8
XFILLER_45_539 VDD VSS sg13g2_decap_8
XFILLER_25_252 VDD VSS sg13g2_decap_8
XFILLER_41_756 VDD VSS sg13g2_fill_1
XFILLER_13_469 VDD VSS sg13g2_decap_8
XFILLER_43_77 VDD VSS sg13g2_decap_8
XFILLER_40_266 VDD VSS sg13g2_decap_8
XFILLER_5_602 VDD VSS sg13g2_decap_8
XFILLER_4_112 VDD VSS sg13g2_decap_8
XFILLER_5_679 VDD VSS sg13g2_decap_8
XFILLER_4_189 VDD VSS sg13g2_decap_8
XFILLER_4_49 VDD VSS sg13g2_decap_8
XFILLER_95_406 VDD VSS sg13g2_decap_8
XFILLER_68_63 VDD VSS sg13g2_decap_8
XFILLER_67_119 VDD VSS sg13g2_decap_8
XFILLER_75_130 VDD VSS sg13g2_decap_8
XFILLER_48_322 VDD VSS sg13g2_decap_8
XFILLER_76_664 VDD VSS sg13g2_decap_8
XFILLER_91_623 VDD VSS sg13g2_decap_8
XFILLER_63_336 VDD VSS sg13g2_decap_8
XFILLER_48_399 VDD VSS sg13g2_decap_8
XFILLER_36_539 VDD VSS sg13g2_decap_8
XFILLER_90_133 VDD VSS sg13g2_decap_8
XFILLER_84_84 VDD VSS sg13g2_decap_8
XFILLER_17_742 VDD VSS sg13g2_decap_8
XFILLER_16_252 VDD VSS sg13g2_decap_8
XFILLER_32_756 VDD VSS sg13g2_fill_1
XFILLER_31_266 VDD VSS sg13g2_decap_8
XFILLER_8_462 VDD VSS sg13g2_decap_8
XFILLER_86_406 VDD VSS sg13g2_decap_8
XFILLER_59_609 VDD VSS sg13g2_decap_8
XFILLER_58_119 VDD VSS sg13g2_decap_8
XFILLER_67_653 VDD VSS sg13g2_decap_8
XFILLER_39_322 VDD VSS sg13g2_decap_8
XFILLER_94_483 VDD VSS sg13g2_decap_8
XFILLER_82_623 VDD VSS sg13g2_decap_8
XFILLER_66_196 VDD VSS sg13g2_decap_8
XFILLER_39_399 VDD VSS sg13g2_decap_8
XFILLER_54_336 VDD VSS sg13g2_decap_8
XFILLER_27_539 VDD VSS sg13g2_decap_8
XFILLER_81_133 VDD VSS sg13g2_decap_8
XFILLER_23_756 VDD VSS sg13g2_fill_1
XFILLER_50_553 VDD VSS sg13g2_decap_8
XFILLER_10_406 VDD VSS sg13g2_decap_8
XFILLER_13_14 VDD VSS sg13g2_decap_8
XFILLER_22_266 VDD VSS sg13g2_decap_8
XFILLER_2_616 VDD VSS sg13g2_decap_8
XFILLER_8_7 VDD VSS sg13g2_decap_8
XFILLER_1_126 VDD VSS sg13g2_decap_8
XFILLER_89_266 VDD VSS sg13g2_decap_8
XFILLER_77_428 VDD VSS sg13g2_decap_8
XFILLER_49_119 VDD VSS sg13g2_decap_8
XFILLER_58_686 VDD VSS sg13g2_decap_8
XFILLER_38_77 VDD VSS sg13g2_decap_8
XFILLER_85_483 VDD VSS sg13g2_decap_8
XFILLER_45_336 VDD VSS sg13g2_decap_8
XFILLER_57_196 VDD VSS sg13g2_decap_8
XFILLER_18_539 VDD VSS sg13g2_decap_8
XFILLER_73_667 VDD VSS sg13g2_decap_8
XFILLER_72_133 VDD VSS sg13g2_decap_8
XFILLER_54_21 VDD VSS sg13g2_decap_8
XFILLER_54_98 VDD VSS sg13g2_decap_8
XFILLER_14_756 VDD VSS sg13g2_fill_1
XFILLER_26_594 VDD VSS sg13g2_decap_8
XFILLER_13_266 VDD VSS sg13g2_decap_8
XFILLER_41_553 VDD VSS sg13g2_decap_8
XFILLER_70_42 VDD VSS sg13g2_decap_8
XFILLER_9_259 VDD VSS sg13g2_decap_8
XFILLER_5_476 VDD VSS sg13g2_decap_8
XFILLER_79_84 VDD VSS sg13g2_decap_8
XFILLER_95_203 VDD VSS sg13g2_decap_8
XFILLER_1_693 VDD VSS sg13g2_decap_8
XFILLER_64_623 VDD VSS sg13g2_decap_8
XFILLER_91_420 VDD VSS sg13g2_decap_8
XFILLER_49_686 VDD VSS sg13g2_decap_8
XFILLER_36_336 VDD VSS sg13g2_decap_8
XFILLER_63_133 VDD VSS sg13g2_decap_8
XFILLER_48_196 VDD VSS sg13g2_decap_8
XFILLER_91_497 VDD VSS sg13g2_decap_8
XFILLER_32_553 VDD VSS sg13g2_decap_8
XFILLER_67_0 VDD VSS sg13g2_decap_8
XFILLER_5_70 VDD VSS sg13g2_decap_8
XFILLER_86_203 VDD VSS sg13g2_decap_8
XFILLER_59_406 VDD VSS sg13g2_decap_8
XFILLER_74_409 VDD VSS sg13g2_decap_8
XFILLER_67_450 VDD VSS sg13g2_decap_8
XFILLER_94_280 VDD VSS sg13g2_decap_8
XFILLER_82_420 VDD VSS sg13g2_decap_8
XFILLER_55_623 VDD VSS sg13g2_decap_8
XFILLER_27_336 VDD VSS sg13g2_decap_8
XFILLER_39_196 VDD VSS sg13g2_decap_8
XFILLER_54_133 VDD VSS sg13g2_decap_8
XFILLER_82_497 VDD VSS sg13g2_decap_8
XFILLER_70_659 VDD VSS sg13g2_decap_8
XFILLER_24_35 VDD VSS sg13g2_decap_8
XFILLER_50_350 VDD VSS sg13g2_decap_8
XFILLER_23_553 VDD VSS sg13g2_decap_8
XFILLER_10_203 VDD VSS sg13g2_decap_8
XFILLER_40_56 VDD VSS sg13g2_decap_8
XFILLER_2_413 VDD VSS sg13g2_decap_8
XFILLER_49_21 VDD VSS sg13g2_decap_8
XFILLER_77_203 VDD VSS sg13g2_decap_8
XFILLER_49_98 VDD VSS sg13g2_decap_8
XFILLER_93_707 VDD VSS sg13g2_decap_8
XFILLER_1_28 VDD VSS sg13g2_decap_8
XFILLER_92_217 VDD VSS sg13g2_decap_8
XFILLER_85_280 VDD VSS sg13g2_decap_8
XFILLER_65_42 VDD VSS sg13g2_decap_8
XFILLER_58_483 VDD VSS sg13g2_decap_8
XFILLER_46_623 VDD VSS sg13g2_decap_8
XFILLER_73_442 VDD VSS sg13g2_decap_8
XFILLER_18_336 VDD VSS sg13g2_decap_8
XFILLER_45_133 VDD VSS sg13g2_decap_8
XFILLER_73_464 VDD VSS sg13g2_decap_8
XFILLER_61_637 VDD VSS sg13g2_decap_8
XFILLER_26_391 VDD VSS sg13g2_decap_8
XFILLER_81_63 VDD VSS sg13g2_decap_8
XFILLER_41_350 VDD VSS sg13g2_decap_8
XFILLER_60_147 VDD VSS sg13g2_decap_8
XFILLER_14_553 VDD VSS sg13g2_decap_8
XFILLER_60_7 VDD VSS sg13g2_decap_8
XFILLER_5_273 VDD VSS sg13g2_decap_8
XFILLER_69_748 VDD VSS sg13g2_decap_8
XFILLER_84_707 VDD VSS sg13g2_decap_8
XFILLER_68_258 VDD VSS sg13g2_decap_8
XFILLER_1_490 VDD VSS sg13g2_decap_8
XFILLER_83_217 VDD VSS sg13g2_decap_8
XFILLER_49_483 VDD VSS sg13g2_decap_8
XFILLER_37_623 VDD VSS sg13g2_decap_8
X_76_ _76__3/L_HI VSS VDD _76_/D _76_/Q _79_/CLK sg13g2_dfrbpq_1
XFILLER_64_420 VDD VSS sg13g2_decap_8
XFILLER_36_133 VDD VSS sg13g2_decap_8
XFILLER_64_497 VDD VSS sg13g2_decap_8
XFILLER_91_294 VDD VSS sg13g2_decap_8
XFILLER_52_637 VDD VSS sg13g2_decap_8
XFILLER_32_350 VDD VSS sg13g2_decap_8
XFILLER_51_147 VDD VSS sg13g2_decap_8
XFILLER_20_567 VDD VSS sg13g2_decap_8
XFILLER_59_203 VDD VSS sg13g2_decap_8
XFILLER_87_567 VDD VSS sg13g2_decap_8
XFILLER_75_718 VDD VSS sg13g2_decap_8
XFILLER_19_35 VDD VSS sg13g2_decap_8
XFILLER_74_217 VDD VSS sg13g2_decap_8
XFILLER_28_623 VDD VSS sg13g2_decap_8
XFILLER_27_133 VDD VSS sg13g2_decap_8
XFILLER_55_420 VDD VSS sg13g2_decap_8
XFILLER_82_294 VDD VSS sg13g2_decap_8
XFILLER_55_497 VDD VSS sg13g2_decap_8
XFILLER_35_56 VDD VSS sg13g2_decap_8
XFILLER_43_637 VDD VSS sg13g2_decap_8
XFILLER_70_478 VDD VSS sg13g2_fill_2
XFILLER_23_350 VDD VSS sg13g2_decap_8
XFILLER_42_147 VDD VSS sg13g2_decap_8
XFILLER_11_567 VDD VSS sg13g2_decap_8
XFILLER_51_77 VDD VSS sg13g2_decap_8
XFILLER_3_700 VDD VSS sg13g2_decap_8
XFILLER_2_210 VDD VSS sg13g2_decap_8
XFILLER_2_287 VDD VSS sg13g2_decap_8
XFILLER_93_504 VDD VSS sg13g2_decap_8
XFILLER_78_567 VDD VSS sg13g2_decap_8
XFILLER_65_217 VDD VSS sg13g2_decap_8
XFILLER_76_63 VDD VSS sg13g2_decap_8
XFILLER_19_623 VDD VSS sg13g2_decap_8
XFILLER_18_133 VDD VSS sg13g2_decap_8
XFILLER_46_420 VDD VSS sg13g2_decap_8
XFILLER_58_280 VDD VSS sg13g2_decap_8
XFILLER_73_261 VDD VSS sg13g2_decap_8
XFILLER_73_272 VDD VSS sg13g2_fill_2
XFILLER_46_497 VDD VSS sg13g2_decap_8
XFILLER_61_434 VDD VSS sg13g2_decap_8
XFILLER_34_637 VDD VSS sg13g2_decap_8
XFILLER_92_84 VDD VSS sg13g2_decap_8
XIO_BOND_outputs\[6\].output_pad output_PAD[6] bondpad_70x70_novias
XFILLER_14_350 VDD VSS sg13g2_decap_8
XFILLER_33_147 VDD VSS sg13g2_decap_8
XFILLER_6_560 VDD VSS sg13g2_decap_8
XFILLER_69_545 VDD VSS sg13g2_decap_8
XFILLER_84_504 VDD VSS sg13g2_decap_8
XFILLER_57_707 VDD VSS sg13g2_decap_8
XFILLER_56_217 VDD VSS sg13g2_decap_8
XFILLER_37_420 VDD VSS sg13g2_decap_8
XFILLER_49_280 VDD VSS sg13g2_decap_8
X_59_ _59_/A _66_/D _59_/Y VDD VSS sg13g2_nor2_1
XFILLER_92_581 VDD VSS sg13g2_decap_8
XFILLER_80_721 VDD VSS sg13g2_decap_8
XFILLER_64_294 VDD VSS sg13g2_decap_8
XFILLER_52_434 VDD VSS sg13g2_decap_8
XFILLER_25_637 VDD VSS sg13g2_decap_8
XFILLER_37_497 VDD VSS sg13g2_decap_8
XFILLER_24_147 VDD VSS sg13g2_decap_8
XFILLER_20_364 VDD VSS sg13g2_decap_8
XFILLER_21_14 VDD VSS sg13g2_decap_8
XFILLER_0_714 VDD VSS sg13g2_decap_8
XFILLER_87_364 VDD VSS sg13g2_decap_8
XFILLER_48_707 VDD VSS sg13g2_decap_8
XFILLER_75_515 VDD VSS sg13g2_decap_8
XFILLER_47_217 VDD VSS sg13g2_decap_8
XFILLER_28_420 VDD VSS sg13g2_decap_8
XFILLER_90_518 VDD VSS sg13g2_decap_8
XFILLER_46_77 VDD VSS sg13g2_decap_8
XFILLER_83_581 VDD VSS sg13g2_decap_8
XFILLER_43_434 VDD VSS sg13g2_decap_8
XFILLER_55_294 VDD VSS sg13g2_decap_8
XFILLER_16_637 VDD VSS sg13g2_decap_8
XFILLER_28_497 VDD VSS sg13g2_decap_8
XFILLER_70_242 VDD VSS sg13g2_decap_8
XFILLER_62_21 VDD VSS sg13g2_decap_8
XFILLER_15_147 VDD VSS sg13g2_decap_8
XFILLER_62_98 VDD VSS sg13g2_decap_8
XFILLER_11_364 VDD VSS sg13g2_decap_8
XFILLER_7_357 VDD VSS sg13g2_decap_8
XFILLER_7_49 VDD VSS sg13g2_decap_8
XFILLER_11_91 VDD VSS sg13g2_decap_8
XFILLER_3_574 VDD VSS sg13g2_decap_8
XFILLER_87_84 VDD VSS sg13g2_decap_8
XFILLER_23_7 VDD VSS sg13g2_decap_8
XFILLER_39_707 VDD VSS sg13g2_decap_8
XFILLER_93_301 VDD VSS sg13g2_decap_8
XFILLER_78_364 VDD VSS sg13g2_decap_8
XFILLER_38_217 VDD VSS sg13g2_decap_8
XFILLER_66_548 VDD VSS sg13g2_decap_8
XFILLER_19_420 VDD VSS sg13g2_decap_8
XFILLER_81_518 VDD VSS sg13g2_decap_8
XFILLER_93_378 VDD VSS sg13g2_decap_8
XFILLER_74_581 VDD VSS sg13g2_decap_8
XFILLER_62_721 VDD VSS sg13g2_decap_8
XFILLER_34_434 VDD VSS sg13g2_decap_8
XFILLER_46_294 VDD VSS sg13g2_decap_8
XFILLER_19_497 VDD VSS sg13g2_decap_8
XFILLER_61_231 VDD VSS sg13g2_decap_8
XFILLER_30_651 VDD VSS sg13g2_decap_8
XFILLER_69_331 VDD VSS sg13g2_decap_8
XFILLER_84_301 VDD VSS sg13g2_decap_8
XFILLER_57_504 VDD VSS sg13g2_decap_8
XFILLER_29_217 VDD VSS sg13g2_decap_8
XFILLER_84_378 VDD VSS sg13g2_decap_8
XFILLER_65_570 VDD VSS sg13g2_decap_8
XFILLER_53_721 VDD VSS sg13g2_decap_8
XFILLER_16_14 VDD VSS sg13g2_decap_8
XFILLER_25_434 VDD VSS sg13g2_decap_8
XFILLER_37_294 VDD VSS sg13g2_decap_8
XFILLER_52_231 VDD VSS sg13g2_decap_8
XFILLER_80_595 VDD VSS sg13g2_decap_8
XFILLER_40_448 VDD VSS sg13g2_decap_8
XFILLER_32_35 VDD VSS sg13g2_decap_8
XFILLER_21_651 VDD VSS sg13g2_decap_8
XFILLER_20_161 VDD VSS sg13g2_decap_8
XFILLER_0_511 VDD VSS sg13g2_decap_8
XFILLER_88_651 VDD VSS sg13g2_decap_8
XFILLER_87_161 VDD VSS sg13g2_decap_8
XFILLER_48_504 VDD VSS sg13g2_decap_8
XFILLER_0_588 VDD VSS sg13g2_decap_8
XFILLER_57_21 VDD VSS sg13g2_decap_8
XFILLER_75_334 VDD VSS sg13g2_decap_8
XFILLER_63_529 VDD VSS sg13g2_decap_8
XFILLER_75_367 VDD VSS sg13g2_decap_8
XFILLER_57_98 VDD VSS sg13g2_decap_8
XFILLER_90_315 VDD VSS sg13g2_decap_8
XFILLER_56_581 VDD VSS sg13g2_decap_8
XFILLER_44_721 VDD VSS sg13g2_decap_8
XFILLER_73_42 VDD VSS sg13g2_decap_8
XFILLER_16_434 VDD VSS sg13g2_decap_8
XFILLER_28_294 VDD VSS sg13g2_decap_8
XFILLER_43_231 VDD VSS sg13g2_decap_8
XFILLER_71_562 VDD VSS sg13g2_decap_8
XFILLER_31_448 VDD VSS sg13g2_decap_8
XFILLER_12_651 VDD VSS sg13g2_decap_8
XFILLER_8_644 VDD VSS sg13g2_decap_8
XFILLER_11_161 VDD VSS sg13g2_decap_8
XFILLER_7_154 VDD VSS sg13g2_decap_8
XFILLER_3_371 VDD VSS sg13g2_decap_8
XFILLER_79_651 VDD VSS sg13g2_decap_8
XFILLER_78_161 VDD VSS sg13g2_decap_8
XFILLER_66_301 VDD VSS sg13g2_decap_8
XFILLER_39_504 VDD VSS sg13g2_decap_8
XFILLER_94_665 VDD VSS sg13g2_decap_8
XFILLER_66_378 VDD VSS sg13g2_decap_8
XFILLER_54_518 VDD VSS sg13g2_decap_8
XFILLER_93_175 VDD VSS sg13g2_decap_8
XFILLER_81_315 VDD VSS sg13g2_decap_8
XFILLER_47_581 VDD VSS sg13g2_decap_8
XFILLER_35_721 VDD VSS sg13g2_decap_8
XFILLER_19_294 VDD VSS sg13g2_decap_8
XFILLER_34_231 VDD VSS sg13g2_decap_8
XFILLER_50_735 VDD VSS sg13g2_decap_8
XFILLER_62_595 VDD VSS sg13g2_decap_8
XFILLER_22_448 VDD VSS sg13g2_decap_8
XFILLER_8_70 VDD VSS sg13g2_decap_8
XFILLER_1_308 VDD VSS sg13g2_decap_8
XFILLER_89_448 VDD VSS sg13g2_decap_8
XFILLER_69_161 VDD VSS sg13g2_decap_8
XFILLER_57_301 VDD VSS sg13g2_decap_8
XFILLER_85_665 VDD VSS sg13g2_decap_8
XFILLER_27_35 VDD VSS sg13g2_decap_8
XFILLER_57_378 VDD VSS sg13g2_decap_8
XFILLER_45_518 VDD VSS sg13g2_decap_8
XFILLER_84_175 VDD VSS sg13g2_decap_8
XFILLER_38_581 VDD VSS sg13g2_decap_8
XFILLER_25_231 VDD VSS sg13g2_decap_8
XFILLER_80_392 VDD VSS sg13g2_decap_8
XFILLER_53_595 VDD VSS sg13g2_decap_8
XFILLER_13_448 VDD VSS sg13g2_decap_8
XFILLER_43_56 VDD VSS sg13g2_decap_8
XFILLER_41_735 VDD VSS sg13g2_decap_8
XFILLER_40_245 VDD VSS sg13g2_decap_8
XFILLER_5_658 VDD VSS sg13g2_decap_8
XFILLER_4_168 VDD VSS sg13g2_decap_8
XFILLER_4_28 VDD VSS sg13g2_decap_8
XFILLER_68_42 VDD VSS sg13g2_decap_8
XFILLER_48_301 VDD VSS sg13g2_decap_8
XFILLER_76_643 VDD VSS sg13g2_decap_8
XFILLER_0_385 VDD VSS sg13g2_decap_8
XFILLER_91_602 VDD VSS sg13g2_decap_8
XFILLER_48_378 VDD VSS sg13g2_decap_8
XFILLER_36_518 VDD VSS sg13g2_decap_8
XFILLER_90_112 VDD VSS sg13g2_decap_8
XFILLER_75_186 VDD VSS sg13g2_decap_8
XFILLER_63_315 VDD VSS sg13g2_decap_8
XFILLER_84_63 VDD VSS sg13g2_decap_8
XFILLER_17_721 VDD VSS sg13g2_decap_8
XFILLER_29_581 VDD VSS sg13g2_decap_8
XFILLER_91_679 VDD VSS sg13g2_decap_8
XFILLER_16_231 VDD VSS sg13g2_decap_8
XFILLER_90_189 VDD VSS sg13g2_decap_8
XFILLER_90_7 VDD VSS sg13g2_decap_8
XFILLER_32_735 VDD VSS sg13g2_decap_8
XFILLER_44_595 VDD VSS sg13g2_decap_8
XFILLER_31_245 VDD VSS sg13g2_decap_8
XFILLER_8_441 VDD VSS sg13g2_decap_8
XFILLER_39_301 VDD VSS sg13g2_decap_8
XFILLER_67_632 VDD VSS sg13g2_decap_8
XFILLER_82_602 VDD VSS sg13g2_decap_8
XFILLER_94_462 VDD VSS sg13g2_decap_8
XFILLER_12_0 VDD VSS sg13g2_decap_8
XFILLER_27_518 VDD VSS sg13g2_decap_8
XFILLER_81_112 VDD VSS sg13g2_decap_8
XFILLER_66_175 VDD VSS sg13g2_decap_8
XFILLER_39_378 VDD VSS sg13g2_decap_8
XFILLER_54_315 VDD VSS sg13g2_decap_8
XFILLER_82_679 VDD VSS sg13g2_decap_8
XFILLER_81_189 VDD VSS sg13g2_decap_8
XFILLER_62_392 VDD VSS sg13g2_decap_8
XFILLER_50_532 VDD VSS sg13g2_decap_8
XFILLER_23_735 VDD VSS sg13g2_decap_8
XFILLER_35_595 VDD VSS sg13g2_decap_8
XFILLER_22_245 VDD VSS sg13g2_decap_8
XFILLER_1_105 VDD VSS sg13g2_decap_8
XFILLER_89_245 VDD VSS sg13g2_decap_8
XFILLER_85_462 VDD VSS sg13g2_decap_8
XFILLER_58_665 VDD VSS sg13g2_decap_8
XFILLER_38_56 VDD VSS sg13g2_decap_8
XFILLER_72_112 VDD VSS sg13g2_decap_8
XFILLER_45_315 VDD VSS sg13g2_decap_8
XFILLER_57_175 VDD VSS sg13g2_decap_8
XFILLER_18_518 VDD VSS sg13g2_decap_8
XFILLER_73_646 VDD VSS sg13g2_decap_8
XFILLER_72_189 VDD VSS sg13g2_decap_8
XFILLER_60_329 VDD VSS sg13g2_decap_8
XFILLER_26_573 VDD VSS sg13g2_decap_8
XFILLER_54_77 VDD VSS sg13g2_decap_8
XFILLER_53_392 VDD VSS sg13g2_decap_8
XFILLER_14_735 VDD VSS sg13g2_decap_8
XFILLER_41_532 VDD VSS sg13g2_decap_8
XFILLER_13_245 VDD VSS sg13g2_decap_8
XFILLER_70_21 VDD VSS sg13g2_decap_8
XFILLER_9_238 VDD VSS sg13g2_decap_8
XFILLER_70_98 VDD VSS sg13g2_decap_8
XFILLER_5_455 VDD VSS sg13g2_decap_8
XFILLER_79_63 VDD VSS sg13g2_decap_8
XFILLER_1_672 VDD VSS sg13g2_decap_8
XFILLER_64_602 VDD VSS sg13g2_decap_8
XFILLER_95_259 VDD VSS sg13g2_decap_8
XFILLER_76_440 VDD VSS sg13g2_decap_8
XFILLER_95_84 VDD VSS sg13g2_decap_8
XFILLER_49_665 VDD VSS sg13g2_decap_8
XFILLER_0_182 VDD VSS sg13g2_decap_8
XFILLER_63_112 VDD VSS sg13g2_decap_8
XFILLER_36_315 VDD VSS sg13g2_decap_8
XFILLER_48_175 VDD VSS sg13g2_decap_8
XFILLER_64_679 VDD VSS sg13g2_decap_8
XFILLER_91_476 VDD VSS sg13g2_decap_8
XFILLER_51_329 VDD VSS sg13g2_decap_8
XFILLER_63_189 VDD VSS sg13g2_decap_8
XFILLER_44_392 VDD VSS sg13g2_decap_8
XFILLER_17_595 VDD VSS sg13g2_decap_8
XFILLER_32_532 VDD VSS sg13g2_decap_8
XFILLER_20_749 VDD VSS sg13g2_decap_8
XFILLER_87_749 VDD VSS sg13g2_decap_8
XFILLER_86_259 VDD VSS sg13g2_decap_8
XFILLER_55_602 VDD VSS sg13g2_decap_8
XFILLER_27_315 VDD VSS sg13g2_decap_8
XFILLER_39_175 VDD VSS sg13g2_decap_8
XFILLER_54_112 VDD VSS sg13g2_decap_8
XFILLER_82_476 VDD VSS sg13g2_decap_8
XFILLER_55_679 VDD VSS sg13g2_decap_8
XFILLER_70_638 VDD VSS sg13g2_decap_8
XFILLER_63_690 VDD VSS sg13g2_decap_8
XFILLER_24_14 VDD VSS sg13g2_decap_8
XFILLER_35_392 VDD VSS sg13g2_decap_8
XFILLER_42_329 VDD VSS sg13g2_decap_8
XFILLER_54_189 VDD VSS sg13g2_decap_8
XFILLER_23_532 VDD VSS sg13g2_decap_8
XFILLER_11_749 VDD VSS sg13g2_decap_8
XFILLER_10_259 VDD VSS sg13g2_decap_8
XFILLER_40_35 VDD VSS sg13g2_decap_8
XFILLER_2_469 VDD VSS sg13g2_decap_8
XFILLER_78_749 VDD VSS sg13g2_decap_8
XFILLER_49_77 VDD VSS sg13g2_decap_8
XFILLER_65_21 VDD VSS sg13g2_decap_8
XFILLER_46_602 VDD VSS sg13g2_decap_8
XFILLER_18_315 VDD VSS sg13g2_decap_8
XFILLER_58_462 VDD VSS sg13g2_decap_8
XFILLER_73_421 VDD VSS sg13g2_decap_8
XFILLER_45_112 VDD VSS sg13g2_decap_8
XFILLER_65_98 VDD VSS sg13g2_decap_8
XFILLER_61_616 VDD VSS sg13g2_decap_8
XFILLER_46_679 VDD VSS sg13g2_decap_8
XFILLER_26_370 VDD VSS sg13g2_decap_8
XFILLER_33_329 VDD VSS sg13g2_decap_8
XFILLER_45_189 VDD VSS sg13g2_decap_8
XFILLER_60_126 VDD VSS sg13g2_decap_8
XFILLER_14_532 VDD VSS sg13g2_decap_8
XFILLER_81_42 VDD VSS sg13g2_decap_8
XFILLER_14_91 VDD VSS sg13g2_decap_8
XFILLER_6_742 VDD VSS sg13g2_decap_8
XFILLER_5_252 VDD VSS sg13g2_decap_8
XFILLER_53_7 VDD VSS sg13g2_decap_8
XFILLER_69_727 VDD VSS sg13g2_decap_8
XFILLER_68_237 VDD VSS sg13g2_decap_8
XFILLER_49_462 VDD VSS sg13g2_decap_8
XFILLER_37_602 VDD VSS sg13g2_decap_8
XFILLER_76_292 VDD VSS sg13g2_decap_8
X_75_ _83_/D _75_/A _75_/B _75_/C VDD VSS sg13g2_and3_1
XFILLER_36_112 VDD VSS sg13g2_decap_8
XFILLER_64_476 VDD VSS sg13g2_decap_8
XFILLER_52_616 VDD VSS sg13g2_decap_8
XFILLER_37_679 VDD VSS sg13g2_decap_8
XFILLER_91_273 VDD VSS sg13g2_decap_8
XFILLER_24_329 VDD VSS sg13g2_decap_8
XFILLER_36_189 VDD VSS sg13g2_decap_8
XFILLER_51_126 VDD VSS sg13g2_decap_8
XFILLER_17_392 VDD VSS sg13g2_decap_8
XFILLER_60_693 VDD VSS sg13g2_decap_8
XFILLER_20_546 VDD VSS sg13g2_decap_8
XFILLER_10_49 VDD VSS sg13g2_decap_8
XFILLER_87_546 VDD VSS sg13g2_decap_8
XFILLER_19_14 VDD VSS sg13g2_decap_8
XFILLER_59_259 VDD VSS sg13g2_decap_8
XFILLER_28_602 VDD VSS sg13g2_decap_8
XFILLER_27_112 VDD VSS sg13g2_decap_8
XFILLER_55_476 VDD VSS sg13g2_decap_8
XFILLER_28_679 VDD VSS sg13g2_decap_8
XFILLER_43_616 VDD VSS sg13g2_decap_8
XFILLER_82_273 VDD VSS sg13g2_decap_8
XFILLER_35_35 VDD VSS sg13g2_decap_8
XFILLER_15_329 VDD VSS sg13g2_decap_8
XFILLER_27_189 VDD VSS sg13g2_decap_8
XFILLER_42_126 VDD VSS sg13g2_decap_8
XFILLER_70_446 VDD VSS sg13g2_decap_8
XFILLER_51_693 VDD VSS sg13g2_decap_8
XFILLER_11_546 VDD VSS sg13g2_decap_8
XFILLER_7_539 VDD VSS sg13g2_decap_8
XFILLER_51_56 VDD VSS sg13g2_decap_8
XFILLER_3_756 VDD VSS sg13g2_fill_1
XFILLER_78_546 VDD VSS sg13g2_decap_8
XFILLER_2_266 VDD VSS sg13g2_decap_8
XFILLER_76_42 VDD VSS sg13g2_decap_8
XFILLER_19_602 VDD VSS sg13g2_decap_8
XFILLER_18_112 VDD VSS sg13g2_decap_8
XFILLER_46_476 VDD VSS sg13g2_decap_8
XFILLER_19_679 VDD VSS sg13g2_decap_8
XFILLER_34_616 VDD VSS sg13g2_decap_8
XFILLER_92_63 VDD VSS sg13g2_decap_8
XFILLER_18_189 VDD VSS sg13g2_decap_8
XFILLER_33_126 VDD VSS sg13g2_decap_8
XFILLER_61_413 VDD VSS sg13g2_decap_8
XFILLER_42_693 VDD VSS sg13g2_decap_8
XFILLER_69_524 VDD VSS sg13g2_decap_8
XFILLER_77_590 VDD VSS sg13g2_decap_8
XFILLER_65_752 VDD VSS sg13g2_decap_4
XFILLER_92_560 VDD VSS sg13g2_decap_8
XFILLER_80_700 VDD VSS sg13g2_decap_8
X_58_ _61_/A _58_/B _58_/C _58_/Y VDD VSS sg13g2_nor3_1
XFILLER_37_476 VDD VSS sg13g2_decap_8
XFILLER_25_616 VDD VSS sg13g2_decap_8
XFILLER_64_273 VDD VSS sg13g2_decap_8
XFILLER_24_126 VDD VSS sg13g2_decap_8
XFILLER_52_413 VDD VSS sg13g2_decap_8
XFILLER_60_490 VDD VSS sg13g2_decap_8
XFILLER_33_693 VDD VSS sg13g2_decap_8
XFILLER_20_343 VDD VSS sg13g2_decap_8
XFILLER_87_343 VDD VSS sg13g2_decap_8
XFILLER_83_560 VDD VSS sg13g2_decap_8
XFILLER_46_56 VDD VSS sg13g2_decap_8
XFILLER_28_476 VDD VSS sg13g2_decap_8
XFILLER_16_616 VDD VSS sg13g2_decap_8
XFILLER_71_744 VDD VSS sg13g2_decap_8
XFILLER_15_126 VDD VSS sg13g2_decap_8
XFILLER_43_413 VDD VSS sg13g2_decap_8
XFILLER_55_273 VDD VSS sg13g2_decap_8
XFILLER_71_755 VDD VSS sg13g2_fill_2
XFILLER_70_221 VDD VSS sg13g2_decap_8
XFILLER_62_77 VDD VSS sg13g2_decap_8
XFILLER_51_490 VDD VSS sg13g2_decap_8
XFILLER_24_693 VDD VSS sg13g2_decap_8
XFILLER_11_343 VDD VSS sg13g2_decap_8
XFILLER_7_28 VDD VSS sg13g2_decap_8
XFILLER_7_336 VDD VSS sg13g2_decap_8
XFILLER_3_553 VDD VSS sg13g2_decap_8
XFILLER_11_70 VDD VSS sg13g2_decap_8
XFILLER_78_343 VDD VSS sg13g2_decap_8
XFILLER_87_63 VDD VSS sg13g2_decap_8
XFILLER_66_527 VDD VSS sg13g2_decap_8
XFILLER_16_7 VDD VSS sg13g2_decap_8
XFILLER_74_560 VDD VSS sg13g2_decap_8
XFILLER_62_700 VDD VSS sg13g2_decap_8
XFILLER_93_357 VDD VSS sg13g2_decap_8
XFILLER_19_476 VDD VSS sg13g2_decap_8
XFILLER_34_413 VDD VSS sg13g2_decap_8
XFILLER_46_273 VDD VSS sg13g2_decap_8
XFILLER_61_210 VDD VSS sg13g2_decap_8
XFILLER_61_287 VDD VSS sg13g2_decap_8
XFILLER_15_693 VDD VSS sg13g2_decap_8
XFILLER_30_630 VDD VSS sg13g2_decap_8
XFILLER_42_490 VDD VSS sg13g2_decap_8
XFILLER_42_0 VDD VSS sg13g2_decap_8
XFILLER_69_310 VDD VSS sg13g2_decap_8
XFILLER_69_387 VDD VSS sg13g2_decap_8
XFILLER_84_357 VDD VSS sg13g2_decap_8
XFILLER_53_700 VDD VSS sg13g2_decap_8
XFILLER_25_413 VDD VSS sg13g2_decap_8
XFILLER_37_273 VDD VSS sg13g2_decap_8
XFILLER_52_210 VDD VSS sg13g2_decap_8
XFILLER_80_574 VDD VSS sg13g2_decap_8
XFILLER_40_427 VDD VSS sg13g2_decap_8
XFILLER_52_287 VDD VSS sg13g2_decap_8
XFILLER_21_630 VDD VSS sg13g2_decap_8
XFILLER_33_490 VDD VSS sg13g2_decap_8
XFILLER_32_14 VDD VSS sg13g2_decap_8
XFILLER_20_140 VDD VSS sg13g2_decap_8
XFILLER_88_630 VDD VSS sg13g2_decap_8
XFILLER_87_140 VDD VSS sg13g2_decap_8
XFILLER_0_567 VDD VSS sg13g2_decap_8
XFILLER_57_77 VDD VSS sg13g2_decap_8
XFILLER_63_508 VDD VSS sg13g2_decap_8
XFILLER_44_700 VDD VSS sg13g2_decap_8
XFILLER_73_21 VDD VSS sg13g2_decap_8
XFILLER_56_560 VDD VSS sg13g2_decap_8
XFILLER_16_413 VDD VSS sg13g2_decap_8
XFILLER_28_273 VDD VSS sg13g2_decap_8
XFILLER_43_210 VDD VSS sg13g2_decap_8
XFILLER_71_541 VDD VSS sg13g2_decap_8
XFILLER_73_98 VDD VSS sg13g2_decap_8
XFILLER_12_630 VDD VSS sg13g2_decap_8
XFILLER_31_427 VDD VSS sg13g2_decap_8
XFILLER_43_287 VDD VSS sg13g2_decap_8
XFILLER_24_490 VDD VSS sg13g2_decap_8
XFILLER_11_140 VDD VSS sg13g2_decap_8
XFILLER_8_623 VDD VSS sg13g2_decap_8
XFILLER_7_133 VDD VSS sg13g2_decap_8
XFILLER_22_91 VDD VSS sg13g2_decap_8
XFILLER_3_350 VDD VSS sg13g2_decap_8
XFILLER_79_630 VDD VSS sg13g2_decap_8
XFILLER_78_140 VDD VSS sg13g2_decap_8
XFILLER_94_644 VDD VSS sg13g2_decap_8
XFILLER_93_154 VDD VSS sg13g2_decap_8
XFILLER_66_357 VDD VSS sg13g2_decap_8
XFILLER_47_560 VDD VSS sg13g2_decap_8
XFILLER_19_273 VDD VSS sg13g2_decap_8
XFILLER_35_700 VDD VSS sg13g2_decap_8
XFILLER_34_210 VDD VSS sg13g2_decap_8
XFILLER_62_574 VDD VSS sg13g2_decap_8
XFILLER_50_714 VDD VSS sg13g2_decap_8
XFILLER_22_427 VDD VSS sg13g2_decap_8
XFILLER_34_287 VDD VSS sg13g2_decap_8
XFILLER_15_490 VDD VSS sg13g2_decap_8
XFILLER_89_427 VDD VSS sg13g2_decap_8
XFILLER_69_140 VDD VSS sg13g2_decap_8
XFILLER_85_644 VDD VSS sg13g2_decap_8
XFILLER_84_154 VDD VSS sg13g2_decap_8
XFILLER_27_14 VDD VSS sg13g2_decap_8
XFILLER_57_357 VDD VSS sg13g2_decap_8
XFILLER_38_560 VDD VSS sg13g2_decap_8
XFILLER_25_210 VDD VSS sg13g2_decap_8
XFILLER_26_755 VDD VSS sg13g2_fill_2
XFILLER_53_574 VDD VSS sg13g2_decap_8
XFILLER_41_714 VDD VSS sg13g2_decap_8
XFILLER_80_371 VDD VSS sg13g2_decap_8
XFILLER_13_427 VDD VSS sg13g2_decap_8
XFILLER_43_35 VDD VSS sg13g2_decap_8
XFILLER_25_287 VDD VSS sg13g2_decap_8
XFILLER_40_224 VDD VSS sg13g2_decap_8
XFILLER_5_637 VDD VSS sg13g2_decap_8
XFILLER_4_147 VDD VSS sg13g2_decap_8
XFILLER_68_21 VDD VSS sg13g2_decap_8
XFILLER_0_364 VDD VSS sg13g2_decap_8
XFILLER_76_622 VDD VSS sg13g2_decap_8
XFILLER_68_98 VDD VSS sg13g2_decap_8
XFILLER_48_357 VDD VSS sg13g2_decap_8
XFILLER_76_699 VDD VSS sg13g2_decap_8
XFILLER_75_165 VDD VSS sg13g2_decap_8
XFILLER_84_42 VDD VSS sg13g2_decap_8
XFILLER_17_700 VDD VSS sg13g2_decap_8
XFILLER_29_560 VDD VSS sg13g2_decap_8
XFILLER_91_658 VDD VSS sg13g2_decap_8
XFILLER_16_210 VDD VSS sg13g2_decap_8
XFILLER_90_168 VDD VSS sg13g2_decap_8
XFILLER_17_91 VDD VSS sg13g2_decap_8
XFILLER_32_714 VDD VSS sg13g2_decap_8
XFILLER_44_574 VDD VSS sg13g2_decap_8
XFILLER_16_287 VDD VSS sg13g2_decap_8
XFILLER_31_224 VDD VSS sg13g2_decap_8
XFILLER_83_7 VDD VSS sg13g2_decap_8
XFILLER_8_420 VDD VSS sg13g2_decap_8
XFILLER_8_497 VDD VSS sg13g2_decap_8
XFILLER_67_611 VDD VSS sg13g2_decap_8
XFILLER_94_441 VDD VSS sg13g2_decap_8
XFILLER_66_154 VDD VSS sg13g2_decap_8
XFILLER_39_357 VDD VSS sg13g2_decap_8
XFILLER_67_688 VDD VSS sg13g2_decap_8
XFILLER_82_658 VDD VSS sg13g2_decap_8
XFILLER_81_168 VDD VSS sg13g2_decap_8
XFILLER_23_714 VDD VSS sg13g2_decap_8
XFILLER_35_574 VDD VSS sg13g2_decap_8
XFILLER_62_371 VDD VSS sg13g2_decap_8
XFILLER_50_511 VDD VSS sg13g2_decap_8
XFILLER_22_224 VDD VSS sg13g2_decap_8
XFILLER_50_588 VDD VSS sg13g2_decap_8
XFILLER_13_49 VDD VSS sg13g2_decap_8
XFILLER_89_224 VDD VSS sg13g2_decap_8
XFILLER_38_35 VDD VSS sg13g2_decap_8
XFILLER_85_441 VDD VSS sg13g2_decap_8
XFILLER_58_644 VDD VSS sg13g2_decap_8
XFILLER_73_625 VDD VSS sg13g2_decap_8
XFILLER_57_154 VDD VSS sg13g2_decap_8
XFILLER_72_168 VDD VSS sg13g2_decap_8
XFILLER_54_56 VDD VSS sg13g2_decap_8
XFILLER_60_308 VDD VSS sg13g2_decap_8
XFILLER_14_714 VDD VSS sg13g2_decap_8
XFILLER_26_552 VDD VSS sg13g2_decap_8
XFILLER_13_224 VDD VSS sg13g2_decap_8
XFILLER_53_371 VDD VSS sg13g2_decap_8
XFILLER_41_511 VDD VSS sg13g2_decap_8
XFILLER_9_217 VDD VSS sg13g2_decap_8
XFILLER_41_588 VDD VSS sg13g2_decap_8
XFILLER_70_77 VDD VSS sg13g2_decap_8
XFILLER_5_434 VDD VSS sg13g2_decap_8
XFILLER_79_42 VDD VSS sg13g2_decap_8
XFILLER_68_419 VDD VSS sg13g2_decap_8
XFILLER_1_651 VDD VSS sg13g2_decap_8
XFILLER_95_238 VDD VSS sg13g2_decap_8
XFILLER_0_161 VDD VSS sg13g2_decap_8
XFILLER_95_63 VDD VSS sg13g2_decap_8
XFILLER_49_644 VDD VSS sg13g2_decap_8
XFILLER_48_154 VDD VSS sg13g2_decap_8
XFILLER_76_496 VDD VSS sg13g2_decap_8
XFILLER_64_658 VDD VSS sg13g2_decap_8
XFILLER_91_455 VDD VSS sg13g2_decap_8
XFILLER_63_168 VDD VSS sg13g2_decap_8
XFILLER_51_308 VDD VSS sg13g2_decap_8
XFILLER_17_574 VDD VSS sg13g2_decap_8
XFILLER_72_691 VDD VSS sg13g2_decap_8
XFILLER_44_371 VDD VSS sg13g2_decap_8
XFILLER_32_511 VDD VSS sg13g2_decap_8
XFILLER_20_728 VDD VSS sg13g2_decap_8
XFILLER_32_588 VDD VSS sg13g2_decap_8
XFILLER_8_294 VDD VSS sg13g2_decap_8
XFILLER_87_728 VDD VSS sg13g2_decap_8
XFILLER_86_238 VDD VSS sg13g2_decap_8
XFILLER_67_485 VDD VSS sg13g2_decap_8
XFILLER_39_154 VDD VSS sg13g2_decap_8
XFILLER_55_658 VDD VSS sg13g2_decap_8
XFILLER_70_617 VDD VSS sg13g2_decap_8
XFILLER_82_455 VDD VSS sg13g2_decap_8
XFILLER_42_308 VDD VSS sg13g2_decap_8
XFILLER_54_168 VDD VSS sg13g2_decap_8
XFILLER_35_371 VDD VSS sg13g2_decap_8
XFILLER_23_511 VDD VSS sg13g2_decap_8
XFILLER_11_728 VDD VSS sg13g2_decap_8
XFILLER_50_385 VDD VSS sg13g2_decap_8
XFILLER_23_588 VDD VSS sg13g2_decap_8
XFILLER_10_238 VDD VSS sg13g2_decap_8
XFILLER_40_14 VDD VSS sg13g2_decap_8
XFILLER_2_448 VDD VSS sg13g2_decap_8
XFILLER_78_728 VDD VSS sg13g2_decap_8
XFILLER_49_56 VDD VSS sg13g2_decap_8
XFILLER_58_441 VDD VSS sg13g2_decap_8
XFILLER_46_658 VDD VSS sg13g2_decap_8
XFILLER_65_77 VDD VSS sg13g2_decap_8
XFILLER_33_308 VDD VSS sg13g2_decap_8
XFILLER_45_168 VDD VSS sg13g2_decap_8
XFILLER_73_499 VDD VSS sg13g2_decap_8
XFILLER_60_105 VDD VSS sg13g2_decap_8
XFILLER_14_511 VDD VSS sg13g2_decap_8
XFILLER_81_21 VDD VSS sg13g2_decap_8
XFILLER_41_385 VDD VSS sg13g2_decap_8
XFILLER_14_588 VDD VSS sg13g2_decap_8
XFILLER_81_98 VDD VSS sg13g2_decap_8
XFILLER_14_70 VDD VSS sg13g2_decap_8
XFILLER_6_721 VDD VSS sg13g2_decap_8
XFILLER_5_231 VDD VSS sg13g2_decap_8
XFILLER_30_91 VDD VSS sg13g2_decap_8
XFILLER_46_7 VDD VSS sg13g2_decap_8
XFILLER_69_706 VDD VSS sg13g2_decap_8
XFILLER_68_216 VDD VSS sg13g2_decap_8
XFILLER_49_441 VDD VSS sg13g2_decap_8
X_74_ _74_/A _74_/B _74_/C _74_/D _75_/C VDD VSS sg13g2_or4_1
XFILLER_92_742 VDD VSS sg13g2_decap_8
XFILLER_76_271 VDD VSS sg13g2_decap_8
XFILLER_37_658 VDD VSS sg13g2_decap_8
XFILLER_91_252 VDD VSS sg13g2_decap_8
XFILLER_64_455 VDD VSS sg13g2_decap_8
XFILLER_24_308 VDD VSS sg13g2_decap_8
XFILLER_36_168 VDD VSS sg13g2_decap_8
XFILLER_51_105 VDD VSS sg13g2_decap_8
XFILLER_17_371 VDD VSS sg13g2_decap_8
XFILLER_60_672 VDD VSS sg13g2_decap_8
XFILLER_32_385 VDD VSS sg13g2_decap_8
XFILLER_20_525 VDD VSS sg13g2_decap_8
XFILLER_72_0 VDD VSS sg13g2_decap_8
XFILLER_9_581 VDD VSS sg13g2_decap_8
XFILLER_10_28 VDD VSS sg13g2_decap_8
XFILLER_87_525 VDD VSS sg13g2_decap_8
XFILLER_59_238 VDD VSS sg13g2_decap_8
XFILLER_83_742 VDD VSS sg13g2_decap_8
XFILLER_67_282 VDD VSS sg13g2_decap_8
XFILLER_28_658 VDD VSS sg13g2_decap_8
XFILLER_82_252 VDD VSS sg13g2_decap_8
XFILLER_35_14 VDD VSS sg13g2_decap_8
XFILLER_15_308 VDD VSS sg13g2_decap_8
XFILLER_27_168 VDD VSS sg13g2_decap_8
XFILLER_55_455 VDD VSS sg13g2_decap_8
XFILLER_70_425 VDD VSS sg13g2_decap_8
XFILLER_42_105 VDD VSS sg13g2_decap_8
XFILLER_51_672 VDD VSS sg13g2_decap_8
XFILLER_11_525 VDD VSS sg13g2_decap_8
XFILLER_51_35 VDD VSS sg13g2_decap_8
XFILLER_23_385 VDD VSS sg13g2_decap_8
XFILLER_50_182 VDD VSS sg13g2_decap_8
XFILLER_7_518 VDD VSS sg13g2_decap_8
XFILLER_3_735 VDD VSS sg13g2_decap_8
XFILLER_2_245 VDD VSS sg13g2_decap_8
XFILLER_78_525 VDD VSS sg13g2_decap_8
XFILLER_66_709 VDD VSS sg13g2_decap_8
XFILLER_76_21 VDD VSS sg13g2_decap_8
XFILLER_93_539 VDD VSS sg13g2_decap_8
XFILLER_74_742 VDD VSS sg13g2_decap_8
XFILLER_76_98 VDD VSS sg13g2_decap_8
XFILLER_19_658 VDD VSS sg13g2_decap_8
XFILLER_18_168 VDD VSS sg13g2_decap_8
XFILLER_46_455 VDD VSS sg13g2_decap_8
XFILLER_92_42 VDD VSS sg13g2_decap_8
XFILLER_33_105 VDD VSS sg13g2_decap_8
XFILLER_61_469 VDD VSS sg13g2_decap_8
XFILLER_42_672 VDD VSS sg13g2_decap_8
XFILLER_25_91 VDD VSS sg13g2_decap_8
XFILLER_14_385 VDD VSS sg13g2_decap_8
XFILLER_41_182 VDD VSS sg13g2_decap_8
XFILLER_6_595 VDD VSS sg13g2_decap_8
XFILLER_69_503 VDD VSS sg13g2_decap_8
XFILLER_84_539 VDD VSS sg13g2_decap_8
XFILLER_65_731 VDD VSS sg13g2_decap_8
XFILLER_2_84 VDD VSS sg13g2_decap_8
X_57_ _57_/A _57_/B _60_/D _66_/D VDD VSS sg13g2_nor3_1
XFILLER_64_252 VDD VSS sg13g2_decap_8
XFILLER_37_455 VDD VSS sg13g2_decap_8
XFILLER_24_105 VDD VSS sg13g2_decap_8
XFILLER_80_756 VDD VSS sg13g2_fill_1
XFILLER_52_469 VDD VSS sg13g2_decap_8
XFILLER_40_609 VDD VSS sg13g2_decap_8
XFILLER_33_672 VDD VSS sg13g2_decap_8
XFILLER_20_322 VDD VSS sg13g2_decap_8
XFILLER_32_182 VDD VSS sg13g2_decap_8
XFILLER_20_399 VDD VSS sg13g2_decap_8
XFILLER_21_49 VDD VSS sg13g2_decap_8
XFILLER_87_322 VDD VSS sg13g2_decap_8
XFILLER_0_749 VDD VSS sg13g2_decap_4
XFILLER_68_580 VDD VSS sg13g2_decap_8
XFILLER_87_399 VDD VSS sg13g2_decap_8
XFILLER_56_742 VDD VSS sg13g2_decap_8
XFILLER_46_35 VDD VSS sg13g2_decap_8
XFILLER_28_455 VDD VSS sg13g2_decap_8
XFILLER_55_252 VDD VSS sg13g2_decap_8
XFILLER_71_723 VDD VSS sg13g2_decap_8
XFILLER_70_211 VDD VSS sg13g2_fill_1
XFILLER_15_105 VDD VSS sg13g2_decap_8
XFILLER_31_609 VDD VSS sg13g2_decap_8
XFILLER_70_277 VDD VSS sg13g2_decap_8
XFILLER_30_119 VDD VSS sg13g2_decap_8
XFILLER_43_469 VDD VSS sg13g2_decap_8
XFILLER_24_672 VDD VSS sg13g2_decap_8
XFILLER_70_299 VDD VSS sg13g2_decap_8
XFILLER_62_56 VDD VSS sg13g2_decap_8
XFILLER_11_322 VDD VSS sg13g2_decap_8
XFILLER_23_182 VDD VSS sg13g2_decap_8
XFILLER_7_315 VDD VSS sg13g2_decap_8
XFILLER_11_399 VDD VSS sg13g2_decap_8
XFILLER_3_532 VDD VSS sg13g2_decap_8
XFILLER_2_0 VDD VSS sg13g2_decap_8
XFILLER_87_42 VDD VSS sg13g2_decap_8
XFILLER_78_322 VDD VSS sg13g2_decap_8
XFILLER_66_506 VDD VSS sg13g2_decap_8
XFILLER_93_336 VDD VSS sg13g2_decap_8
XFILLER_78_399 VDD VSS sg13g2_decap_8
XFILLER_47_742 VDD VSS sg13g2_decap_8
XFILLER_19_455 VDD VSS sg13g2_decap_8
XFILLER_46_252 VDD VSS sg13g2_decap_8
XFILLER_62_756 VDD VSS sg13g2_fill_1
XFILLER_34_469 VDD VSS sg13g2_decap_8
XFILLER_61_266 VDD VSS sg13g2_decap_8
XFILLER_15_672 VDD VSS sg13g2_decap_8
XFILLER_22_609 VDD VSS sg13g2_decap_8
XFILLER_14_182 VDD VSS sg13g2_decap_8
XFILLER_21_119 VDD VSS sg13g2_decap_8
XFILLER_30_686 VDD VSS sg13g2_decap_8
XFILLER_89_609 VDD VSS sg13g2_decap_8
XFILLER_6_392 VDD VSS sg13g2_decap_8
XFILLER_88_119 VDD VSS sg13g2_decap_8
XFILLER_35_0 VDD VSS sg13g2_decap_8
XFILLER_69_366 VDD VSS sg13g2_decap_8
XFILLER_84_336 VDD VSS sg13g2_decap_8
XFILLER_57_539 VDD VSS sg13g2_decap_8
XFILLER_72_509 VDD VSS sg13g2_decap_8
XFILLER_38_742 VDD VSS sg13g2_decap_8
XFILLER_37_252 VDD VSS sg13g2_decap_8
XFILLER_80_553 VDD VSS sg13g2_decap_8
XFILLER_53_756 VDD VSS sg13g2_fill_1
XFILLER_16_49 VDD VSS sg13g2_decap_8
XFILLER_13_609 VDD VSS sg13g2_decap_8
XFILLER_25_469 VDD VSS sg13g2_decap_8
XFILLER_40_406 VDD VSS sg13g2_decap_8
XFILLER_52_266 VDD VSS sg13g2_decap_8
XFILLER_12_119 VDD VSS sg13g2_decap_8
XFILLER_21_686 VDD VSS sg13g2_decap_8
XFILLER_20_196 VDD VSS sg13g2_decap_8
XFILLER_4_329 VDD VSS sg13g2_decap_8
XFILLER_79_119 VDD VSS sg13g2_decap_8
XFILLER_0_546 VDD VSS sg13g2_decap_8
XFILLER_88_686 VDD VSS sg13g2_decap_8
XFILLER_87_196 VDD VSS sg13g2_decap_8
XFILLER_48_539 VDD VSS sg13g2_decap_8
XFILLER_57_56 VDD VSS sg13g2_decap_8
XFILLER_29_742 VDD VSS sg13g2_decap_8
XFILLER_28_252 VDD VSS sg13g2_decap_8
XFILLER_71_520 VDD VSS sg13g2_decap_8
XFILLER_44_756 VDD VSS sg13g2_fill_1
XFILLER_73_77 VDD VSS sg13g2_decap_8
XFILLER_16_469 VDD VSS sg13g2_decap_8
XFILLER_31_406 VDD VSS sg13g2_decap_8
XFILLER_43_266 VDD VSS sg13g2_decap_8
XFILLER_71_597 VDD VSS sg13g2_decap_8
XFILLER_8_602 VDD VSS sg13g2_decap_8
XFILLER_12_686 VDD VSS sg13g2_decap_8
XFILLER_7_112 VDD VSS sg13g2_decap_8
XFILLER_8_679 VDD VSS sg13g2_decap_8
XFILLER_11_196 VDD VSS sg13g2_decap_8
XFILLER_22_70 VDD VSS sg13g2_decap_8
XFILLER_7_189 VDD VSS sg13g2_decap_8
XFILLER_79_686 VDD VSS sg13g2_decap_8
XFILLER_94_623 VDD VSS sg13g2_decap_8
XFILLER_78_196 VDD VSS sg13g2_decap_8
XFILLER_66_336 VDD VSS sg13g2_decap_8
XFILLER_39_539 VDD VSS sg13g2_decap_8
XFILLER_93_133 VDD VSS sg13g2_decap_8
XFILLER_19_252 VDD VSS sg13g2_decap_8
XFILLER_35_756 VDD VSS sg13g2_fill_1
XFILLER_62_553 VDD VSS sg13g2_decap_8
XFILLER_22_406 VDD VSS sg13g2_decap_8
XFILLER_34_266 VDD VSS sg13g2_decap_8
XFILLER_30_483 VDD VSS sg13g2_decap_8
XFILLER_89_406 VDD VSS sg13g2_decap_8
XFILLER_85_623 VDD VSS sg13g2_decap_8
XFILLER_57_336 VDD VSS sg13g2_decap_8
XFILLER_84_133 VDD VSS sg13g2_decap_8
XFILLER_69_196 VDD VSS sg13g2_decap_8
XFILLER_26_734 VDD VSS sg13g2_decap_8
XFILLER_80_350 VDD VSS sg13g2_decap_8
XFILLER_53_553 VDD VSS sg13g2_decap_8
XFILLER_13_406 VDD VSS sg13g2_decap_8
XFILLER_43_14 VDD VSS sg13g2_decap_8
XFILLER_25_266 VDD VSS sg13g2_decap_8
XFILLER_40_203 VDD VSS sg13g2_decap_8
XFILLER_21_483 VDD VSS sg13g2_decap_8
XFILLER_5_616 VDD VSS sg13g2_decap_8
XFILLER_4_126 VDD VSS sg13g2_decap_8
XFILLER_76_601 VDD VSS sg13g2_decap_8
XFILLER_68_77 VDD VSS sg13g2_decap_8
XFILLER_0_343 VDD VSS sg13g2_decap_8
XFILLER_88_483 VDD VSS sg13g2_decap_8
XFILLER_76_678 VDD VSS sg13g2_decap_8
XFILLER_75_144 VDD VSS sg13g2_decap_8
XFILLER_84_21 VDD VSS sg13g2_decap_8
XFILLER_48_336 VDD VSS sg13g2_decap_8
XFILLER_91_637 VDD VSS sg13g2_decap_8
XFILLER_90_147 VDD VSS sg13g2_decap_8
XFILLER_84_98 VDD VSS sg13g2_decap_8
XFILLER_17_756 VDD VSS sg13g2_fill_1
XFILLER_71_361 VDD VSS sg13g2_fill_1
XFILLER_17_70 VDD VSS sg13g2_decap_8
XFILLER_16_266 VDD VSS sg13g2_decap_8
XFILLER_44_553 VDD VSS sg13g2_decap_8
XFILLER_71_394 VDD VSS sg13g2_fill_2
XFILLER_31_203 VDD VSS sg13g2_decap_8
XFILLER_76_7 VDD VSS sg13g2_decap_8
XFILLER_12_483 VDD VSS sg13g2_decap_8
XFILLER_33_91 VDD VSS sg13g2_decap_8
XFILLER_8_476 VDD VSS sg13g2_decap_8
XFILLER_4_693 VDD VSS sg13g2_decap_8
XFILLER_79_483 VDD VSS sg13g2_decap_8
XFILLER_94_420 VDD VSS sg13g2_decap_8
XFILLER_67_667 VDD VSS sg13g2_decap_8
XFILLER_66_133 VDD VSS sg13g2_decap_8
XFILLER_39_336 VDD VSS sg13g2_decap_8
XFILLER_82_637 VDD VSS sg13g2_decap_8
XFILLER_94_497 VDD VSS sg13g2_decap_8
XFILLER_81_147 VDD VSS sg13g2_decap_8
XFILLER_62_350 VDD VSS sg13g2_decap_8
XFILLER_35_553 VDD VSS sg13g2_decap_8
XFILLER_22_203 VDD VSS sg13g2_decap_8
XFILLER_50_567 VDD VSS sg13g2_decap_8
XFILLER_13_28 VDD VSS sg13g2_decap_8
XFILLER_30_280 VDD VSS sg13g2_decap_8
XFILLER_89_203 VDD VSS sg13g2_decap_8
XFILLER_85_420 VDD VSS sg13g2_decap_8
XFILLER_58_623 VDD VSS sg13g2_decap_8
XFILLER_38_14 VDD VSS sg13g2_decap_8
XFILLER_57_133 VDD VSS sg13g2_decap_8
XFILLER_73_604 VDD VSS sg13g2_decap_8
XFILLER_85_497 VDD VSS sg13g2_decap_8
XFILLER_26_531 VDD VSS sg13g2_decap_8
XFILLER_72_147 VDD VSS sg13g2_decap_8
XFILLER_54_35 VDD VSS sg13g2_decap_8
XFILLER_53_350 VDD VSS sg13g2_decap_8
XFILLER_13_203 VDD VSS sg13g2_decap_8
XFILLER_41_567 VDD VSS sg13g2_decap_8
XFILLER_70_56 VDD VSS sg13g2_decap_8
XFILLER_21_280 VDD VSS sg13g2_decap_8
XFILLER_5_413 VDD VSS sg13g2_decap_8
XFILLER_79_21 VDD VSS sg13g2_decap_8
XFILLER_79_98 VDD VSS sg13g2_decap_8
XFILLER_1_630 VDD VSS sg13g2_decap_8
XFILLER_95_217 VDD VSS sg13g2_decap_8
XFILLER_49_623 VDD VSS sg13g2_decap_8
XFILLER_0_140 VDD VSS sg13g2_decap_8
XFILLER_88_280 VDD VSS sg13g2_decap_8
XFILLER_95_42 VDD VSS sg13g2_decap_8
XFILLER_48_133 VDD VSS sg13g2_decap_8
XFILLER_64_637 VDD VSS sg13g2_decap_8
XFILLER_91_434 VDD VSS sg13g2_decap_8
XFILLER_28_91 VDD VSS sg13g2_decap_8
XFILLER_63_147 VDD VSS sg13g2_decap_8
XFILLER_44_350 VDD VSS sg13g2_decap_8
XFILLER_17_553 VDD VSS sg13g2_decap_8
XFILLER_72_670 VDD VSS sg13g2_decap_8
XFILLER_20_707 VDD VSS sg13g2_decap_8
XFILLER_32_567 VDD VSS sg13g2_decap_8
XFILLER_12_280 VDD VSS sg13g2_decap_8
XFILLER_8_273 VDD VSS sg13g2_decap_8
XFILLER_87_707 VDD VSS sg13g2_decap_8
XFILLER_4_490 VDD VSS sg13g2_decap_8
XFILLER_5_84 VDD VSS sg13g2_decap_8
XFILLER_86_217 VDD VSS sg13g2_decap_8
XFILLER_79_280 VDD VSS sg13g2_decap_8
XFILLER_39_133 VDD VSS sg13g2_decap_8
XFILLER_67_464 VDD VSS sg13g2_decap_8
XFILLER_94_294 VDD VSS sg13g2_decap_8
XFILLER_82_434 VDD VSS sg13g2_decap_8
XFILLER_55_637 VDD VSS sg13g2_decap_8
XFILLER_35_350 VDD VSS sg13g2_decap_8
XFILLER_54_147 VDD VSS sg13g2_decap_8
XFILLER_11_707 VDD VSS sg13g2_decap_8
XFILLER_24_49 VDD VSS sg13g2_decap_8
XFILLER_50_364 VDD VSS sg13g2_decap_8
XFILLER_23_567 VDD VSS sg13g2_decap_8
XFILLER_10_217 VDD VSS sg13g2_decap_8
XFILLER_2_427 VDD VSS sg13g2_decap_8
XFILLER_6_7 VDD VSS sg13g2_decap_8
XFILLER_78_707 VDD VSS sg13g2_decap_8
XFILLER_49_35 VDD VSS sg13g2_decap_8
XFILLER_77_217 VDD VSS sg13g2_decap_8
XFILLER_58_420 VDD VSS sg13g2_decap_8
XFILLER_73_401 VDD VSS sg13g2_decap_8
XFILLER_85_294 VDD VSS sg13g2_decap_8
XFILLER_65_56 VDD VSS sg13g2_decap_8
XFILLER_58_497 VDD VSS sg13g2_decap_8
XFILLER_46_637 VDD VSS sg13g2_decap_8
XFILLER_73_478 VDD VSS sg13g2_decap_8
XFILLER_45_147 VDD VSS sg13g2_decap_8
XFILLER_81_77 VDD VSS sg13g2_decap_8
XFILLER_41_364 VDD VSS sg13g2_decap_8
XFILLER_14_567 VDD VSS sg13g2_decap_8
XFILLER_6_700 VDD VSS sg13g2_decap_8
XFILLER_5_210 VDD VSS sg13g2_decap_8
XFILLER_5_287 VDD VSS sg13g2_decap_8
XFILLER_30_70 VDD VSS sg13g2_decap_8
XFILLER_39_7 VDD VSS sg13g2_decap_8
XFILLER_77_751 VDD VSS sg13g2_decap_4
XFILLER_49_420 VDD VSS sg13g2_decap_8
XFILLER_76_250 VDD VSS sg13g2_decap_8
X_73_ _74_/A VDD _75_/B VSS _74_/B _69_/B sg13g2_o21ai_1
XFILLER_92_721 VDD VSS sg13g2_decap_8
XFILLER_64_434 VDD VSS sg13g2_decap_8
XFILLER_49_497 VDD VSS sg13g2_decap_8
XFILLER_37_637 VDD VSS sg13g2_decap_8
XFILLER_91_231 VDD VSS sg13g2_decap_8
XFILLER_36_147 VDD VSS sg13g2_decap_8
XFILLER_17_350 VDD VSS sg13g2_decap_8
XFILLER_60_651 VDD VSS sg13g2_decap_8
XFILLER_32_364 VDD VSS sg13g2_decap_8
XFILLER_20_504 VDD VSS sg13g2_decap_8
XFILLER_9_560 VDD VSS sg13g2_decap_8
XFILLER_65_0 VDD VSS sg13g2_decap_8
Xrst_n_pad IOVDD IOVSS hold11/A rst_n_PAD VDD VSS sg13g2_IOPadIn
XFILLER_87_504 VDD VSS sg13g2_decap_8
XFILLER_59_217 VDD VSS sg13g2_decap_8
XFILLER_67_261 VDD VSS sg13g2_decap_8
XFILLER_19_49 VDD VSS sg13g2_decap_8
XFILLER_95_581 VDD VSS sg13g2_decap_8
XFILLER_83_721 VDD VSS sg13g2_decap_8
XFILLER_55_434 VDD VSS sg13g2_decap_8
XFILLER_28_637 VDD VSS sg13g2_decap_8
XFILLER_82_231 VDD VSS sg13g2_decap_8
XFILLER_27_147 VDD VSS sg13g2_decap_8
XFILLER_70_404 VDD VSS sg13g2_decap_8
XFILLER_51_651 VDD VSS sg13g2_decap_8
XFILLER_11_504 VDD VSS sg13g2_decap_8
XFILLER_23_364 VDD VSS sg13g2_decap_8
XFILLER_51_14 VDD VSS sg13g2_decap_8
XFILLER_50_161 VDD VSS sg13g2_decap_8
XFILLER_3_714 VDD VSS sg13g2_decap_8
XFILLER_2_224 VDD VSS sg13g2_decap_8
XFILLER_78_504 VDD VSS sg13g2_decap_8
XFILLER_93_518 VDD VSS sg13g2_decap_8
XFILLER_86_581 VDD VSS sg13g2_decap_8
XFILLER_74_721 VDD VSS sg13g2_decap_8
XFILLER_76_77 VDD VSS sg13g2_decap_8
XFILLER_46_434 VDD VSS sg13g2_decap_8
XFILLER_58_294 VDD VSS sg13g2_decap_8
XFILLER_19_637 VDD VSS sg13g2_decap_8
XFILLER_73_231 VDD VSS sg13g2_decap_8
XFILLER_92_21 VDD VSS sg13g2_decap_8
XFILLER_18_147 VDD VSS sg13g2_decap_8
XFILLER_73_297 VDD VSS sg13g2_decap_8
XFILLER_61_448 VDD VSS sg13g2_decap_8
XFILLER_92_98 VDD VSS sg13g2_decap_8
XFILLER_25_70 VDD VSS sg13g2_decap_8
XFILLER_14_364 VDD VSS sg13g2_decap_8
XFILLER_42_651 VDD VSS sg13g2_decap_8
XFILLER_41_161 VDD VSS sg13g2_decap_8
XFILLER_10_581 VDD VSS sg13g2_decap_8
XFILLER_41_91 VDD VSS sg13g2_decap_8
XFILLER_6_574 VDD VSS sg13g2_decap_8
XFILLER_69_559 VDD VSS sg13g2_decap_8
XFILLER_84_518 VDD VSS sg13g2_decap_8
XFILLER_65_710 VDD VSS sg13g2_decap_8
XFILLER_2_63 VDD VSS sg13g2_decap_8
XFILLER_37_434 VDD VSS sg13g2_decap_8
X_56_ _60_/D _77_/Q _76_/Q VDD VSS sg13g2_nand2_1
XFILLER_64_231 VDD VSS sg13g2_decap_8
XFILLER_49_294 VDD VSS sg13g2_decap_8
XFILLER_92_595 VDD VSS sg13g2_decap_8
XFILLER_80_735 VDD VSS sg13g2_decap_8
XFILLER_52_448 VDD VSS sg13g2_decap_8
XFILLER_33_651 VDD VSS sg13g2_decap_8
XFILLER_20_301 VDD VSS sg13g2_decap_8
XFILLER_32_161 VDD VSS sg13g2_decap_8
XFILLER_21_28 VDD VSS sg13g2_decap_8
XFILLER_20_378 VDD VSS sg13g2_decap_8
XFILLER_87_301 VDD VSS sg13g2_decap_8
XFILLER_0_728 VDD VSS sg13g2_decap_8
XFILLER_87_378 VDD VSS sg13g2_decap_8
XFILLER_75_529 VDD VSS sg13g2_decap_8
XFILLER_56_721 VDD VSS sg13g2_decap_8
XFILLER_46_14 VDD VSS sg13g2_decap_8
XFILLER_28_434 VDD VSS sg13g2_decap_8
XFILLER_55_231 VDD VSS sg13g2_decap_8
XFILLER_83_595 VDD VSS sg13g2_decap_8
XFILLER_71_702 VDD VSS sg13g2_decap_8
XFILLER_43_448 VDD VSS sg13g2_decap_8
XFILLER_70_256 VDD VSS sg13g2_decap_8
XFILLER_62_35 VDD VSS sg13g2_decap_8
XFILLER_24_651 VDD VSS sg13g2_decap_8
XFILLER_11_301 VDD VSS sg13g2_decap_8
XFILLER_23_161 VDD VSS sg13g2_decap_8
XFILLER_11_378 VDD VSS sg13g2_decap_8
XFILLER_3_511 VDD VSS sg13g2_decap_8
XFILLER_78_301 VDD VSS sg13g2_decap_8
XFILLER_87_21 VDD VSS sg13g2_decap_8
XFILLER_3_588 VDD VSS sg13g2_decap_8
XFILLER_78_378 VDD VSS sg13g2_decap_8
XFILLER_87_98 VDD VSS sg13g2_decap_8
XFILLER_93_315 VDD VSS sg13g2_decap_8
XFILLER_59_581 VDD VSS sg13g2_decap_8
XFILLER_47_721 VDD VSS sg13g2_decap_8
XFILLER_19_434 VDD VSS sg13g2_decap_8
XFILLER_46_231 VDD VSS sg13g2_decap_8
XFILLER_74_595 VDD VSS sg13g2_decap_8
XFILLER_62_735 VDD VSS sg13g2_decap_8
XFILLER_36_91 VDD VSS sg13g2_decap_8
XFILLER_34_448 VDD VSS sg13g2_decap_8
XFILLER_61_245 VDD VSS sg13g2_decap_8
XFILLER_15_651 VDD VSS sg13g2_decap_8
XFILLER_14_161 VDD VSS sg13g2_decap_8
XFILLER_30_665 VDD VSS sg13g2_decap_8
XFILLER_6_371 VDD VSS sg13g2_decap_8
XFILLER_69_345 VDD VSS sg13g2_decap_8
XFILLER_57_518 VDD VSS sg13g2_decap_8
XFILLER_28_0 VDD VSS sg13g2_decap_8
XFILLER_84_315 VDD VSS sg13g2_decap_8
XFILLER_38_721 VDD VSS sg13g2_decap_8
XFILLER_37_231 VDD VSS sg13g2_decap_8
XFILLER_65_584 VDD VSS sg13g2_decap_8
XFILLER_80_532 VDD VSS sg13g2_decap_8
XFILLER_92_392 VDD VSS sg13g2_decap_8
XFILLER_53_735 VDD VSS sg13g2_decap_8
XFILLER_16_28 VDD VSS sg13g2_decap_8
XFILLER_25_448 VDD VSS sg13g2_decap_8
XFILLER_52_245 VDD VSS sg13g2_decap_8
XFILLER_21_665 VDD VSS sg13g2_decap_8
XFILLER_32_49 VDD VSS sg13g2_decap_8
XFILLER_20_175 VDD VSS sg13g2_decap_8
XFILLER_4_308 VDD VSS sg13g2_decap_8
XFILLER_0_525 VDD VSS sg13g2_decap_8
XFILLER_88_665 VDD VSS sg13g2_decap_8
XFILLER_48_518 VDD VSS sg13g2_decap_8
XFILLER_57_35 VDD VSS sg13g2_decap_8
XFILLER_87_175 VDD VSS sg13g2_decap_8
XFILLER_29_721 VDD VSS sg13g2_decap_8
XFILLER_75_348 VDD VSS sg13g2_decap_8
XFILLER_28_231 VDD VSS sg13g2_decap_8
XFILLER_90_329 VDD VSS sg13g2_decap_8
XFILLER_83_392 VDD VSS sg13g2_decap_8
XFILLER_73_56 VDD VSS sg13g2_decap_8
XFILLER_56_595 VDD VSS sg13g2_decap_8
XFILLER_16_448 VDD VSS sg13g2_decap_8
XFILLER_44_735 VDD VSS sg13g2_decap_8
XFILLER_71_576 VDD VSS sg13g2_decap_8
XFILLER_43_245 VDD VSS sg13g2_decap_8
XFILLER_12_665 VDD VSS sg13g2_decap_8
XFILLER_8_658 VDD VSS sg13g2_decap_8
XFILLER_11_175 VDD VSS sg13g2_decap_8
XFILLER_7_168 VDD VSS sg13g2_decap_8
XFILLER_3_385 VDD VSS sg13g2_decap_8
XFILLER_94_602 VDD VSS sg13g2_decap_8
XFILLER_79_665 VDD VSS sg13g2_decap_8
XFILLER_93_112 VDD VSS sg13g2_decap_8
XFILLER_78_175 VDD VSS sg13g2_decap_8
XFILLER_66_315 VDD VSS sg13g2_decap_8
XFILLER_21_7 VDD VSS sg13g2_decap_8
XFILLER_39_518 VDD VSS sg13g2_decap_8
XFILLER_94_679 VDD VSS sg13g2_decap_8
XFILLER_19_231 VDD VSS sg13g2_decap_8
XFILLER_93_189 VDD VSS sg13g2_decap_8
XFILLER_81_329 VDD VSS sg13g2_decap_8
XFILLER_62_532 VDD VSS sg13g2_decap_8
XFILLER_47_595 VDD VSS sg13g2_decap_8
XFILLER_35_735 VDD VSS sg13g2_decap_8
XFILLER_34_245 VDD VSS sg13g2_decap_8
XFILLER_50_749 VDD VSS sg13g2_decap_8
XFILLER_30_462 VDD VSS sg13g2_decap_8
XFILLER_8_84 VDD VSS sg13g2_decap_8
XFILLER_85_602 VDD VSS sg13g2_decap_8
XFILLER_84_112 VDD VSS sg13g2_decap_8
XFILLER_69_175 VDD VSS sg13g2_decap_8
XFILLER_57_315 VDD VSS sg13g2_decap_8
XFILLER_85_679 VDD VSS sg13g2_decap_8
XFILLER_72_318 VDD VSS sg13g2_decap_8
XFILLER_27_49 VDD VSS sg13g2_decap_8
XFILLER_26_713 VDD VSS sg13g2_decap_8
XFILLER_84_189 VDD VSS sg13g2_decap_8
XFILLER_65_392 VDD VSS sg13g2_decap_8
XFILLER_53_532 VDD VSS sg13g2_decap_8
XFILLER_38_595 VDD VSS sg13g2_decap_8
XFILLER_25_245 VDD VSS sg13g2_decap_8
XFILLER_41_749 VDD VSS sg13g2_decap_8
XFILLER_40_259 VDD VSS sg13g2_decap_8
XFILLER_21_462 VDD VSS sg13g2_decap_8
XFILLER_4_105 VDD VSS sg13g2_decap_8
XFILLER_68_56 VDD VSS sg13g2_decap_8
XFILLER_0_322 VDD VSS sg13g2_decap_8
XFILLER_88_462 VDD VSS sg13g2_decap_8
XFILLER_48_315 VDD VSS sg13g2_decap_8
XFILLER_76_657 VDD VSS sg13g2_decap_8
XFILLER_75_123 VDD VSS sg13g2_decap_8
XFILLER_0_399 VDD VSS sg13g2_decap_8
XFILLER_91_616 VDD VSS sg13g2_decap_8
XFILLER_90_126 VDD VSS sg13g2_decap_8
XFILLER_63_329 VDD VSS sg13g2_decap_8
XFILLER_84_77 VDD VSS sg13g2_decap_8
XFILLER_56_392 VDD VSS sg13g2_decap_8
XFILLER_17_735 VDD VSS sg13g2_decap_8
XFILLER_29_595 VDD VSS sg13g2_decap_8
XFILLER_44_532 VDD VSS sg13g2_decap_8
XFILLER_16_245 VDD VSS sg13g2_decap_8
XFILLER_32_749 VDD VSS sg13g2_decap_8
XFILLER_31_259 VDD VSS sg13g2_decap_8
XFILLER_12_462 VDD VSS sg13g2_decap_8
XFILLER_33_70 VDD VSS sg13g2_decap_8
XFILLER_8_455 VDD VSS sg13g2_decap_8
XFILLER_69_7 VDD VSS sg13g2_decap_8
XFILLER_4_672 VDD VSS sg13g2_decap_8
XFILLER_3_182 VDD VSS sg13g2_decap_8
XFILLER_79_462 VDD VSS sg13g2_decap_8
XFILLER_39_315 VDD VSS sg13g2_decap_8
XFILLER_67_646 VDD VSS sg13g2_decap_8
XFILLER_66_112 VDD VSS sg13g2_decap_8
XFILLER_82_616 VDD VSS sg13g2_decap_8
XFILLER_94_476 VDD VSS sg13g2_decap_8
XFILLER_75_690 VDD VSS sg13g2_decap_8
XFILLER_81_126 VDD VSS sg13g2_decap_8
XFILLER_66_189 VDD VSS sg13g2_decap_8
XFILLER_47_392 VDD VSS sg13g2_decap_8
XFILLER_54_329 VDD VSS sg13g2_decap_8
XFILLER_35_532 VDD VSS sg13g2_decap_8
Xoutputs\[4\].output_pad _80_/Q IOVDD IOVSS output_PAD[4] VDD VSS sg13g2_IOPadOut30mA
XFILLER_90_693 VDD VSS sg13g2_decap_8
XFILLER_23_749 VDD VSS sg13g2_decap_8
XFILLER_95_0 VDD VSS sg13g2_decap_8
XFILLER_50_546 VDD VSS sg13g2_decap_8
XFILLER_22_259 VDD VSS sg13g2_decap_8
XFILLER_2_609 VDD VSS sg13g2_decap_8
XFILLER_1_119 VDD VSS sg13g2_decap_8
XFILLER_89_259 VDD VSS sg13g2_decap_8
XFILLER_58_602 VDD VSS sg13g2_decap_8
XFILLER_57_112 VDD VSS sg13g2_decap_8
XFILLER_85_476 VDD VSS sg13g2_decap_8
XFILLER_58_679 VDD VSS sg13g2_decap_8
XFILLER_72_126 VDD VSS sg13g2_decap_8
XFILLER_54_14 VDD VSS sg13g2_decap_8
XFILLER_45_329 VDD VSS sg13g2_decap_8
XFILLER_57_189 VDD VSS sg13g2_decap_8
XFILLER_26_510 VDD VSS sg13g2_decap_8
XFILLER_38_392 VDD VSS sg13g2_decap_8
XFILLER_81_693 VDD VSS sg13g2_decap_8
XFILLER_26_587 VDD VSS sg13g2_decap_8
XFILLER_14_749 VDD VSS sg13g2_decap_8
XFILLER_41_546 VDD VSS sg13g2_decap_8
XFILLER_70_35 VDD VSS sg13g2_decap_8
XFILLER_13_259 VDD VSS sg13g2_decap_8
XFILLER_5_469 VDD VSS sg13g2_decap_8
XFILLER_79_77 VDD VSS sg13g2_decap_8
XFILLER_95_21 VDD VSS sg13g2_decap_8
XFILLER_49_602 VDD VSS sg13g2_decap_8
XFILLER_1_686 VDD VSS sg13g2_decap_8
XFILLER_0_196 VDD VSS sg13g2_decap_8
XFILLER_48_112 VDD VSS sg13g2_decap_8
XFILLER_64_616 VDD VSS sg13g2_decap_8
XFILLER_76_454 VDD VSS sg13g2_fill_1
XFILLER_95_98 VDD VSS sg13g2_decap_8
XFILLER_49_679 VDD VSS sg13g2_decap_8
XFILLER_91_413 VDD VSS sg13g2_decap_8
XFILLER_63_126 VDD VSS sg13g2_decap_8
XFILLER_28_70 VDD VSS sg13g2_decap_8
XFILLER_36_329 VDD VSS sg13g2_decap_8
XFILLER_48_189 VDD VSS sg13g2_decap_8
XFILLER_29_392 VDD VSS sg13g2_decap_8
XFILLER_17_532 VDD VSS sg13g2_decap_8
XFILLER_32_546 VDD VSS sg13g2_decap_8
XFILLER_44_91 VDD VSS sg13g2_decap_8
XFILLER_9_742 VDD VSS sg13g2_decap_8
XFILLER_8_252 VDD VSS sg13g2_decap_8
XFILLER_5_63 VDD VSS sg13g2_decap_8
XFILLER_67_443 VDD VSS sg13g2_decap_8
XFILLER_39_112 VDD VSS sg13g2_decap_8
XFILLER_55_616 VDD VSS sg13g2_decap_8
XFILLER_10_0 VDD VSS sg13g2_decap_8
XFILLER_94_273 VDD VSS sg13g2_decap_8
XFILLER_82_413 VDD VSS sg13g2_decap_8
XFILLER_27_329 VDD VSS sg13g2_decap_8
XFILLER_39_189 VDD VSS sg13g2_decap_8
XFILLER_54_126 VDD VSS sg13g2_decap_8
XFILLER_90_490 VDD VSS sg13g2_decap_8
XFILLER_24_28 VDD VSS sg13g2_decap_8
XFILLER_50_343 VDD VSS sg13g2_decap_8
XFILLER_23_546 VDD VSS sg13g2_decap_8
XFILLER_40_49 VDD VSS sg13g2_decap_8
XFILLER_2_406 VDD VSS sg13g2_decap_8
XFILLER_49_14 VDD VSS sg13g2_decap_8
XFILLER_46_616 VDD VSS sg13g2_decap_8
XFILLER_58_476 VDD VSS sg13g2_decap_8
XFILLER_85_273 VDD VSS sg13g2_decap_8
XFILLER_73_435 VDD VSS sg13g2_decap_8
XFILLER_65_35 VDD VSS sg13g2_decap_8
XFILLER_18_329 VDD VSS sg13g2_decap_8
XFILLER_45_126 VDD VSS sg13g2_decap_8
XFILLER_73_457 VDD VSS sg13g2_decap_8
XFILLER_81_490 VDD VSS sg13g2_decap_8
XFILLER_54_693 VDD VSS sg13g2_decap_8
XFILLER_26_384 VDD VSS sg13g2_decap_8
XFILLER_14_546 VDD VSS sg13g2_decap_8
XFILLER_81_56 VDD VSS sg13g2_decap_8
XFILLER_41_343 VDD VSS sg13g2_decap_8
XFILLER_6_756 VDD VSS sg13g2_fill_1
XFILLER_5_266 VDD VSS sg13g2_decap_8
XFILLER_77_730 VDD VSS sg13g2_decap_8
XFILLER_1_483 VDD VSS sg13g2_decap_8
XFILLER_92_700 VDD VSS sg13g2_decap_8
X_72_ VSS VDD _74_/B _69_/B _72_/Y _72_/B1 sg13g2_a21oi_1
XFILLER_39_91 VDD VSS sg13g2_decap_8
XFILLER_49_476 VDD VSS sg13g2_decap_8
XFILLER_37_616 VDD VSS sg13g2_decap_8
XFILLER_91_210 VDD VSS sg13g2_decap_8
XFILLER_64_413 VDD VSS sg13g2_decap_8
XFILLER_36_126 VDD VSS sg13g2_decap_8
XFILLER_91_287 VDD VSS sg13g2_decap_8
XFILLER_60_630 VDD VSS sg13g2_decap_8
XFILLER_45_693 VDD VSS sg13g2_decap_8
XFILLER_32_343 VDD VSS sg13g2_decap_8
XFILLER_58_0 VDD VSS sg13g2_decap_8
XFILLER_68_741 VDD VSS sg13g2_decap_8
XFILLER_19_28 VDD VSS sg13g2_decap_8
XFILLER_95_560 VDD VSS sg13g2_decap_8
XFILLER_83_700 VDD VSS sg13g2_decap_8
XFILLER_67_240 VDD VSS sg13g2_decap_8
XFILLER_28_616 VDD VSS sg13g2_decap_8
XFILLER_82_210 VDD VSS sg13g2_decap_8
XFILLER_27_126 VDD VSS sg13g2_decap_8
XFILLER_55_413 VDD VSS sg13g2_decap_8
XFILLER_82_287 VDD VSS sg13g2_decap_8
XFILLER_35_49 VDD VSS sg13g2_decap_8
XFILLER_51_630 VDD VSS sg13g2_decap_8
XFILLER_36_693 VDD VSS sg13g2_decap_8
XFILLER_23_343 VDD VSS sg13g2_decap_8
XFILLER_50_140 VDD VSS sg13g2_decap_8
XFILLER_2_203 VDD VSS sg13g2_decap_8
XFILLER_86_560 VDD VSS sg13g2_decap_8
XFILLER_74_700 VDD VSS sg13g2_decap_8
XFILLER_76_56 VDD VSS sg13g2_decap_8
XFILLER_73_210 VDD VSS sg13g2_decap_8
XFILLER_46_413 VDD VSS sg13g2_decap_8
XFILLER_58_273 VDD VSS sg13g2_decap_8
XFILLER_19_616 VDD VSS sg13g2_decap_8
XFILLER_18_126 VDD VSS sg13g2_decap_8
XFILLER_61_427 VDD VSS sg13g2_decap_8
XFILLER_92_77 VDD VSS sg13g2_decap_8
XFILLER_54_490 VDD VSS sg13g2_decap_8
XFILLER_27_693 VDD VSS sg13g2_decap_8
XFILLER_42_630 VDD VSS sg13g2_decap_8
XFILLER_14_343 VDD VSS sg13g2_decap_8
XFILLER_41_140 VDD VSS sg13g2_decap_8
XFILLER_10_560 VDD VSS sg13g2_decap_8
XFILLER_6_553 VDD VSS sg13g2_decap_8
XFILLER_41_70 VDD VSS sg13g2_decap_8
XFILLER_51_7 VDD VSS sg13g2_decap_8
XFILLER_69_538 VDD VSS sg13g2_decap_8
XFILLER_2_42 VDD VSS sg13g2_decap_8
XFILLER_1_280 VDD VSS sg13g2_decap_8
XFILLER_64_210 VDD VSS sg13g2_decap_8
XFILLER_37_413 VDD VSS sg13g2_decap_8
XFILLER_49_273 VDD VSS sg13g2_decap_8
X_55_ VSS VDD _76_/Q _55_/A2 _58_/B _77_/Q sg13g2_a21oi_1
XFILLER_92_574 VDD VSS sg13g2_decap_8
XFILLER_80_714 VDD VSS sg13g2_decap_8
XFILLER_64_287 VDD VSS sg13g2_decap_8
XFILLER_52_427 VDD VSS sg13g2_decap_8
XFILLER_18_693 VDD VSS sg13g2_decap_8
XFILLER_33_630 VDD VSS sg13g2_decap_8
XFILLER_45_490 VDD VSS sg13g2_decap_8
XFILLER_32_140 VDD VSS sg13g2_decap_8
XFILLER_20_357 VDD VSS sg13g2_decap_8
XFILLER_0_707 VDD VSS sg13g2_decap_8
XFILLER_75_508 VDD VSS sg13g2_decap_8
XFILLER_87_357 VDD VSS sg13g2_decap_8
XFILLER_56_700 VDD VSS sg13g2_decap_8
XFILLER_28_413 VDD VSS sg13g2_decap_8
XFILLER_55_210 VDD VSS sg13g2_decap_8
XFILLER_83_574 VDD VSS sg13g2_decap_8
XFILLER_70_202 VDD VSS sg13g2_decap_8
XFILLER_70_235 VDD VSS sg13g2_decap_8
XFILLER_43_427 VDD VSS sg13g2_decap_8
XFILLER_55_287 VDD VSS sg13g2_decap_8
XFILLER_24_630 VDD VSS sg13g2_decap_8
XFILLER_36_490 VDD VSS sg13g2_decap_8
XFILLER_62_14 VDD VSS sg13g2_decap_8
XFILLER_23_140 VDD VSS sg13g2_decap_8
XFILLER_11_357 VDD VSS sg13g2_decap_8
XFILLER_11_84 VDD VSS sg13g2_decap_8
XFILLER_3_567 VDD VSS sg13g2_decap_8
XFILLER_87_77 VDD VSS sg13g2_decap_8
XFILLER_78_357 VDD VSS sg13g2_decap_8
XFILLER_59_560 VDD VSS sg13g2_decap_8
XFILLER_47_700 VDD VSS sg13g2_decap_8
XFILLER_19_413 VDD VSS sg13g2_decap_8
XFILLER_46_210 VDD VSS sg13g2_decap_8
XFILLER_74_574 VDD VSS sg13g2_decap_8
XFILLER_62_714 VDD VSS sg13g2_decap_8
XFILLER_36_70 VDD VSS sg13g2_decap_8
XFILLER_34_427 VDD VSS sg13g2_decap_8
XFILLER_46_287 VDD VSS sg13g2_decap_8
XFILLER_61_224 VDD VSS sg13g2_decap_8
XFILLER_15_630 VDD VSS sg13g2_decap_8
XFILLER_27_490 VDD VSS sg13g2_decap_8
XFILLER_14_140 VDD VSS sg13g2_decap_8
Xoutputs\[9\].output_pad outputs\[9\].output_pad/c2p IOVDD IOVSS output_PAD[9] VDD
+ VSS sg13g2_IOPadOut30mA
XFILLER_30_644 VDD VSS sg13g2_decap_8
XFILLER_52_91 VDD VSS sg13g2_decap_8
XFILLER_6_350 VDD VSS sg13g2_decap_8
XFILLER_69_324 VDD VSS sg13g2_decap_8
XFILLER_38_700 VDD VSS sg13g2_decap_8
XFILLER_37_210 VDD VSS sg13g2_decap_8
XFILLER_65_563 VDD VSS sg13g2_decap_8
XFILLER_53_714 VDD VSS sg13g2_decap_8
XFILLER_80_511 VDD VSS sg13g2_decap_8
XFILLER_92_371 VDD VSS sg13g2_decap_8
XFILLER_25_427 VDD VSS sg13g2_decap_8
XFILLER_37_287 VDD VSS sg13g2_decap_8
XFILLER_52_224 VDD VSS sg13g2_decap_8
XFILLER_18_490 VDD VSS sg13g2_decap_8
XFILLER_80_588 VDD VSS sg13g2_decap_8
XFILLER_32_28 VDD VSS sg13g2_decap_8
XFILLER_21_644 VDD VSS sg13g2_decap_8
XFILLER_20_154 VDD VSS sg13g2_decap_8
XFILLER_0_504 VDD VSS sg13g2_decap_8
XFILLER_88_644 VDD VSS sg13g2_decap_8
XFILLER_87_154 VDD VSS sg13g2_decap_8
XFILLER_57_14 VDD VSS sg13g2_decap_8
XFILLER_75_327 VDD VSS sg13g2_decap_8
XFILLER_29_700 VDD VSS sg13g2_decap_8
XFILLER_28_210 VDD VSS sg13g2_decap_8
XFILLER_90_308 VDD VSS sg13g2_decap_8
XFILLER_56_574 VDD VSS sg13g2_decap_8
XFILLER_44_714 VDD VSS sg13g2_decap_8
XFILLER_83_371 VDD VSS sg13g2_decap_8
XFILLER_73_35 VDD VSS sg13g2_decap_8
XFILLER_16_427 VDD VSS sg13g2_decap_8
XFILLER_28_287 VDD VSS sg13g2_decap_8
XFILLER_43_224 VDD VSS sg13g2_decap_8
XFILLER_71_555 VDD VSS sg13g2_decap_8
XFILLER_12_644 VDD VSS sg13g2_decap_8
XFILLER_8_637 VDD VSS sg13g2_decap_8
XFILLER_11_154 VDD VSS sg13g2_decap_8
XFILLER_7_147 VDD VSS sg13g2_decap_8
XFILLER_3_364 VDD VSS sg13g2_decap_8
XFILLER_79_644 VDD VSS sg13g2_decap_8
XFILLER_78_154 VDD VSS sg13g2_decap_8
XFILLER_94_658 VDD VSS sg13g2_decap_8
XFILLER_14_7 VDD VSS sg13g2_decap_8
XFILLER_19_210 VDD VSS sg13g2_decap_8
XFILLER_93_168 VDD VSS sg13g2_decap_8
XFILLER_81_308 VDD VSS sg13g2_decap_8
XFILLER_47_574 VDD VSS sg13g2_decap_8
XFILLER_47_91 VDD VSS sg13g2_decap_8
XFILLER_35_714 VDD VSS sg13g2_decap_8
XFILLER_62_511 VDD VSS sg13g2_decap_8
XFILLER_19_287 VDD VSS sg13g2_decap_8
XFILLER_34_224 VDD VSS sg13g2_decap_8
XFILLER_62_588 VDD VSS sg13g2_decap_8
XFILLER_50_728 VDD VSS sg13g2_decap_8
XFILLER_30_441 VDD VSS sg13g2_decap_8
XFILLER_8_63 VDD VSS sg13g2_decap_8
XFILLER_40_0 VDD VSS sg13g2_decap_8
XFILLER_69_154 VDD VSS sg13g2_decap_8
XFILLER_85_658 VDD VSS sg13g2_decap_8
XFILLER_84_168 VDD VSS sg13g2_decap_8
XFILLER_27_28 VDD VSS sg13g2_decap_8
XFILLER_38_574 VDD VSS sg13g2_decap_8
XFILLER_65_371 VDD VSS sg13g2_decap_8
XFILLER_53_511 VDD VSS sg13g2_decap_8
XFILLER_25_224 VDD VSS sg13g2_decap_8
XFILLER_80_385 VDD VSS sg13g2_decap_8
XFILLER_53_588 VDD VSS sg13g2_decap_8
XFILLER_41_728 VDD VSS sg13g2_decap_8
XFILLER_43_49 VDD VSS sg13g2_decap_8
XFILLER_40_238 VDD VSS sg13g2_decap_8
XFILLER_21_441 VDD VSS sg13g2_decap_8
XFILLER_68_35 VDD VSS sg13g2_decap_8
XFILLER_0_301 VDD VSS sg13g2_decap_8
XFILLER_88_441 VDD VSS sg13g2_decap_8
XFILLER_75_102 VDD VSS sg13g2_decap_8
XFILLER_0_378 VDD VSS sg13g2_decap_8
XFILLER_76_636 VDD VSS sg13g2_decap_8
XFILLER_75_179 VDD VSS sg13g2_decap_8
XFILLER_63_308 VDD VSS sg13g2_decap_8
XFILLER_84_56 VDD VSS sg13g2_decap_8
XFILLER_17_714 VDD VSS sg13g2_decap_8
XFILLER_90_105 VDD VSS sg13g2_decap_8
XFILLER_16_224 VDD VSS sg13g2_decap_8
XFILLER_56_371 VDD VSS sg13g2_decap_8
XFILLER_29_574 VDD VSS sg13g2_decap_8
XFILLER_44_511 VDD VSS sg13g2_decap_8
XFILLER_71_352 VDD VSS sg13g2_decap_8
XFILLER_32_728 VDD VSS sg13g2_decap_8
XFILLER_44_588 VDD VSS sg13g2_decap_8
XFILLER_71_396 VDD VSS sg13g2_fill_1
XFILLER_31_238 VDD VSS sg13g2_decap_8
XFILLER_12_441 VDD VSS sg13g2_decap_8
XFILLER_8_434 VDD VSS sg13g2_decap_8
XFILLER_4_651 VDD VSS sg13g2_decap_8
XFILLER_3_161 VDD VSS sg13g2_decap_8
XFILLER_79_441 VDD VSS sg13g2_decap_8
XFILLER_67_625 VDD VSS sg13g2_decap_8
XFILLER_94_455 VDD VSS sg13g2_decap_8
XFILLER_66_168 VDD VSS sg13g2_decap_8
XFILLER_54_308 VDD VSS sg13g2_decap_8
XFILLER_81_105 VDD VSS sg13g2_decap_8
XFILLER_47_371 VDD VSS sg13g2_decap_8
XFILLER_35_511 VDD VSS sg13g2_decap_8
XFILLER_90_672 VDD VSS sg13g2_decap_8
XFILLER_62_385 VDD VSS sg13g2_decap_8
XFILLER_50_525 VDD VSS sg13g2_decap_8
XFILLER_23_728 VDD VSS sg13g2_decap_8
XFILLER_35_588 VDD VSS sg13g2_decap_8
XFILLER_22_238 VDD VSS sg13g2_decap_8
XFILLER_88_0 VDD VSS sg13g2_decap_8
XFILLER_89_238 VDD VSS sg13g2_decap_8
XFILLER_58_658 VDD VSS sg13g2_decap_8
XFILLER_38_49 VDD VSS sg13g2_decap_8
XFILLER_85_455 VDD VSS sg13g2_decap_8
XFILLER_45_308 VDD VSS sg13g2_decap_8
XFILLER_57_168 VDD VSS sg13g2_decap_8
XFILLER_73_639 VDD VSS sg13g2_decap_8
XFILLER_72_105 VDD VSS sg13g2_decap_8
XFILLER_38_371 VDD VSS sg13g2_decap_8
XFILLER_81_672 VDD VSS sg13g2_decap_8
XFILLER_14_728 VDD VSS sg13g2_decap_8
XFILLER_26_566 VDD VSS sg13g2_decap_8
XFILLER_41_525 VDD VSS sg13g2_decap_8
XFILLER_80_182 VDD VSS sg13g2_decap_8
XFILLER_13_238 VDD VSS sg13g2_decap_8
XFILLER_53_385 VDD VSS sg13g2_decap_8
XFILLER_70_14 VDD VSS sg13g2_decap_8
XFILLER_5_448 VDD VSS sg13g2_decap_8
XFILLER_79_56 VDD VSS sg13g2_decap_8
XFILLER_1_665 VDD VSS sg13g2_decap_8
XFILLER_76_433 VDD VSS sg13g2_decap_8
XFILLER_49_658 VDD VSS sg13g2_decap_8
XFILLER_0_175 VDD VSS sg13g2_decap_8
XFILLER_95_77 VDD VSS sg13g2_decap_8
XFILLER_36_308 VDD VSS sg13g2_decap_8
XFILLER_48_168 VDD VSS sg13g2_decap_8
XFILLER_63_105 VDD VSS sg13g2_decap_8
XFILLER_29_371 VDD VSS sg13g2_decap_8
XFILLER_17_511 VDD VSS sg13g2_decap_8
XFILLER_91_469 VDD VSS sg13g2_decap_8
XFILLER_17_588 VDD VSS sg13g2_decap_8
XFILLER_71_182 VDD VSS sg13g2_decap_8
XFILLER_44_70 VDD VSS sg13g2_decap_8
XFILLER_44_385 VDD VSS sg13g2_decap_8
XFILLER_32_525 VDD VSS sg13g2_decap_8
XFILLER_81_7 VDD VSS sg13g2_decap_8
XFILLER_9_721 VDD VSS sg13g2_decap_8
XFILLER_8_231 VDD VSS sg13g2_decap_8
XFILLER_60_91 VDD VSS sg13g2_decap_8
XFILLER_5_42 VDD VSS sg13g2_decap_8
XFILLER_95_742 VDD VSS sg13g2_decap_8
XFILLER_67_422 VDD VSS sg13g2_decap_8
XFILLER_94_252 VDD VSS sg13g2_decap_8
XFILLER_27_308 VDD VSS sg13g2_decap_8
XFILLER_39_168 VDD VSS sg13g2_decap_8
XFILLER_67_499 VDD VSS sg13g2_decap_8
XFILLER_54_105 VDD VSS sg13g2_decap_8
XFILLER_82_469 VDD VSS sg13g2_decap_8
XFILLER_63_683 VDD VSS sg13g2_decap_8
XFILLER_62_182 VDD VSS sg13g2_decap_8
XFILLER_35_385 VDD VSS sg13g2_decap_8
XFILLER_50_322 VDD VSS sg13g2_decap_8
XFILLER_23_525 VDD VSS sg13g2_decap_8
XFILLER_50_399 VDD VSS sg13g2_decap_8
XFILLER_40_28 VDD VSS sg13g2_decap_8
XFILLER_86_742 VDD VSS sg13g2_decap_8
XFILLER_85_252 VDD VSS sg13g2_decap_8
XFILLER_65_14 VDD VSS sg13g2_decap_8
XFILLER_18_308 VDD VSS sg13g2_decap_8
XFILLER_58_455 VDD VSS sg13g2_decap_8
XFILLER_73_414 VDD VSS sg13g2_decap_8
XFILLER_45_105 VDD VSS sg13g2_decap_8
XFILLER_61_609 VDD VSS sg13g2_decap_8
XFILLER_54_672 VDD VSS sg13g2_decap_8
XFILLER_26_363 VDD VSS sg13g2_decap_8
XFILLER_60_119 VDD VSS sg13g2_decap_8
XFILLER_81_35 VDD VSS sg13g2_decap_8
XFILLER_41_322 VDD VSS sg13g2_decap_8
XFILLER_53_182 VDD VSS sg13g2_decap_8
XFILLER_14_525 VDD VSS sg13g2_decap_8
XFILLER_41_399 VDD VSS sg13g2_decap_8
XFILLER_10_742 VDD VSS sg13g2_decap_8
XFILLER_14_84 VDD VSS sg13g2_decap_8
XFILLER_6_735 VDD VSS sg13g2_decap_8
XFILLER_5_245 VDD VSS sg13g2_decap_8
XFILLER_1_462 VDD VSS sg13g2_decap_8
X_71_ _75_/A VDD _71_/Y VSS _74_/B _69_/B sg13g2_o21ai_1
XFILLER_39_70 VDD VSS sg13g2_decap_8
XFILLER_49_455 VDD VSS sg13g2_decap_8
XFILLER_76_285 VDD VSS sg13g2_decap_8
XFILLER_36_105 VDD VSS sg13g2_decap_8
XFILLER_92_756 VDD VSS sg13g2_fill_1
XFILLER_64_469 VDD VSS sg13g2_decap_8
XFILLER_52_609 VDD VSS sg13g2_decap_8
XFILLER_91_266 VDD VSS sg13g2_decap_8
XFILLER_51_119 VDD VSS sg13g2_decap_8
XFILLER_45_672 VDD VSS sg13g2_decap_8
XFILLER_55_91 VDD VSS sg13g2_decap_8
XFILLER_17_385 VDD VSS sg13g2_decap_8
XFILLER_32_322 VDD VSS sg13g2_decap_8
XFILLER_44_182 VDD VSS sg13g2_decap_8
XFILLER_60_686 VDD VSS sg13g2_decap_8
XFILLER_32_399 VDD VSS sg13g2_decap_8
XFILLER_20_539 VDD VSS sg13g2_decap_8
XFILLER_9_595 VDD VSS sg13g2_decap_8
XFILLER_87_539 VDD VSS sg13g2_decap_8
XFILLER_68_720 VDD VSS sg13g2_decap_8
XFILLER_27_105 VDD VSS sg13g2_decap_8
XFILLER_83_756 VDD VSS sg13g2_fill_1
XFILLER_67_296 VDD VSS sg13g2_decap_8
XFILLER_82_266 VDD VSS sg13g2_decap_8
XFILLER_35_28 VDD VSS sg13g2_decap_8
XFILLER_55_469 VDD VSS sg13g2_decap_8
XFILLER_36_672 VDD VSS sg13g2_decap_8
XFILLER_43_609 VDD VSS sg13g2_decap_8
XFILLER_70_439 VDD VSS sg13g2_decap_8
XFILLER_63_480 VDD VSS sg13g2_decap_8
XFILLER_23_322 VDD VSS sg13g2_decap_8
XFILLER_35_182 VDD VSS sg13g2_decap_8
XFILLER_42_119 VDD VSS sg13g2_decap_8
XFILLER_51_686 VDD VSS sg13g2_decap_8
XFILLER_11_539 VDD VSS sg13g2_decap_8
XFILLER_23_399 VDD VSS sg13g2_decap_8
XFILLER_51_49 VDD VSS sg13g2_decap_8
XFILLER_50_196 VDD VSS sg13g2_decap_8
XFILLER_3_749 VDD VSS sg13g2_decap_8
XFILLER_2_259 VDD VSS sg13g2_decap_8
XFILLER_78_539 VDD VSS sg13g2_decap_8
XFILLER_76_35 VDD VSS sg13g2_decap_8
XFILLER_59_742 VDD VSS sg13g2_decap_8
XFILLER_18_105 VDD VSS sg13g2_decap_8
XFILLER_58_252 VDD VSS sg13g2_decap_8
XFILLER_74_756 VDD VSS sg13g2_fill_1
XFILLER_46_469 VDD VSS sg13g2_decap_8
XFILLER_61_406 VDD VSS sg13g2_decap_8
XFILLER_27_672 VDD VSS sg13g2_decap_8
XFILLER_34_609 VDD VSS sg13g2_decap_8
XFILLER_92_56 VDD VSS sg13g2_decap_8
XFILLER_14_322 VDD VSS sg13g2_decap_8
XFILLER_26_182 VDD VSS sg13g2_decap_8
XFILLER_33_119 VDD VSS sg13g2_decap_8
XFILLER_14_399 VDD VSS sg13g2_decap_8
XFILLER_42_686 VDD VSS sg13g2_decap_8
XFILLER_41_196 VDD VSS sg13g2_decap_8
XFILLER_6_532 VDD VSS sg13g2_decap_8
XFILLER_44_7 VDD VSS sg13g2_decap_8
XFILLER_69_517 VDD VSS sg13g2_decap_8
Xoutputs\[9\].output_pad_2 VDD VSS outputs\[9\].output_pad/c2p sg13g2_tielo
XFILLER_2_21 VDD VSS sg13g2_decap_8
XFILLER_77_583 VDD VSS sg13g2_decap_8
XFILLER_49_252 VDD VSS sg13g2_decap_8
XFILLER_65_756 VDD VSS sg13g2_fill_1
XFILLER_65_745 VDD VSS sg13g2_decap_8
X_54_ VSS VDD _76_/Q _55_/A2 _54_/Y _53_/Y sg13g2_a21oi_1
XFILLER_2_98 VDD VSS sg13g2_decap_8
XFILLER_92_553 VDD VSS sg13g2_decap_8
XFILLER_64_266 VDD VSS sg13g2_decap_8
XFILLER_37_469 VDD VSS sg13g2_decap_8
XFILLER_52_406 VDD VSS sg13g2_decap_8
XFILLER_18_672 VDD VSS sg13g2_decap_8
XFILLER_25_609 VDD VSS sg13g2_decap_8
XFILLER_17_182 VDD VSS sg13g2_decap_8
XFILLER_24_119 VDD VSS sg13g2_decap_8
XFILLER_60_483 VDD VSS sg13g2_decap_8
XFILLER_33_686 VDD VSS sg13g2_decap_8
XFILLER_20_336 VDD VSS sg13g2_decap_8
XFILLER_32_196 VDD VSS sg13g2_decap_8
XFILLER_70_0 VDD VSS sg13g2_decap_8
XFILLER_9_392 VDD VSS sg13g2_decap_8
XFILLER_87_336 VDD VSS sg13g2_decap_8
XFILLER_68_594 VDD VSS sg13g2_decap_8
XFILLER_56_756 VDD VSS sg13g2_fill_1
XFILLER_46_49 VDD VSS sg13g2_decap_8
XFILLER_83_553 VDD VSS sg13g2_decap_8
XFILLER_28_469 VDD VSS sg13g2_decap_8
XFILLER_43_406 VDD VSS sg13g2_decap_8
XFILLER_55_266 VDD VSS sg13g2_decap_8
XFILLER_16_609 VDD VSS sg13g2_decap_8
XFILLER_71_737 VDD VSS sg13g2_decap_8
XFILLER_15_119 VDD VSS sg13g2_decap_8
XFILLER_51_483 VDD VSS sg13g2_decap_8
XFILLER_24_686 VDD VSS sg13g2_decap_8
XFILLER_11_336 VDD VSS sg13g2_decap_8
XFILLER_23_196 VDD VSS sg13g2_decap_8
XFILLER_7_329 VDD VSS sg13g2_decap_8
XFILLER_3_546 VDD VSS sg13g2_decap_8
XFILLER_11_63 VDD VSS sg13g2_decap_8
XFILLER_78_336 VDD VSS sg13g2_decap_8
XFILLER_87_56 VDD VSS sg13g2_decap_8
XFILLER_47_756 VDD VSS sg13g2_fill_1
XFILLER_74_553 VDD VSS sg13g2_decap_8
XFILLER_19_469 VDD VSS sg13g2_decap_8
XFILLER_34_406 VDD VSS sg13g2_decap_8
XFILLER_46_266 VDD VSS sg13g2_decap_8
XFILLER_61_203 VDD VSS sg13g2_decap_8
XFILLER_15_686 VDD VSS sg13g2_decap_8
XFILLER_30_623 VDD VSS sg13g2_decap_8
XFILLER_14_196 VDD VSS sg13g2_decap_8
XFILLER_42_483 VDD VSS sg13g2_decap_8
XFILLER_52_70 VDD VSS sg13g2_decap_8
XFILLER_69_303 VDD VSS sg13g2_decap_8
XFILLER_65_542 VDD VSS sg13g2_decap_8
XFILLER_38_756 VDD VSS sg13g2_fill_1
XFILLER_92_350 VDD VSS sg13g2_decap_8
XFILLER_25_406 VDD VSS sg13g2_decap_8
XFILLER_37_266 VDD VSS sg13g2_decap_8
XFILLER_52_203 VDD VSS sg13g2_decap_8
XFILLER_80_567 VDD VSS sg13g2_decap_8
XFILLER_60_280 VDD VSS sg13g2_decap_8
XFILLER_21_623 VDD VSS sg13g2_decap_8
XFILLER_33_483 VDD VSS sg13g2_decap_8
XFILLER_20_133 VDD VSS sg13g2_decap_8
XFILLER_88_623 VDD VSS sg13g2_decap_8
XFILLER_87_133 VDD VSS sg13g2_decap_8
XFILLER_68_391 VDD VSS sg13g2_decap_8
XFILLER_29_756 VDD VSS sg13g2_fill_1
XFILLER_83_350 VDD VSS sg13g2_decap_8
XFILLER_56_553 VDD VSS sg13g2_decap_8
XFILLER_16_406 VDD VSS sg13g2_decap_8
XFILLER_28_266 VDD VSS sg13g2_decap_8
XFILLER_71_534 VDD VSS sg13g2_decap_8
XFILLER_73_14 VDD VSS sg13g2_decap_8
XFILLER_43_203 VDD VSS sg13g2_decap_8
XFILLER_12_623 VDD VSS sg13g2_decap_8
XFILLER_51_280 VDD VSS sg13g2_decap_8
XFILLER_24_483 VDD VSS sg13g2_decap_8
XFILLER_8_616 VDD VSS sg13g2_decap_8
XFILLER_11_133 VDD VSS sg13g2_decap_8
XFILLER_7_126 VDD VSS sg13g2_decap_8
XFILLER_22_84 VDD VSS sg13g2_decap_8
XFILLER_3_343 VDD VSS sg13g2_decap_8
XFILLER_79_623 VDD VSS sg13g2_decap_8
XFILLER_0_0 VDD VSS sg13g2_decap_8
XFILLER_78_133 VDD VSS sg13g2_decap_8
XFILLER_94_637 VDD VSS sg13g2_decap_8
XFILLER_93_147 VDD VSS sg13g2_decap_8
XFILLER_47_553 VDD VSS sg13g2_decap_8
XFILLER_47_70 VDD VSS sg13g2_decap_8
XFILLER_19_266 VDD VSS sg13g2_decap_8
XFILLER_34_203 VDD VSS sg13g2_decap_8
XFILLER_62_567 VDD VSS sg13g2_decap_8
XFILLER_50_707 VDD VSS sg13g2_decap_8
XFILLER_63_91 VDD VSS sg13g2_decap_8
XFILLER_30_420 VDD VSS sg13g2_decap_8
XFILLER_42_280 VDD VSS sg13g2_decap_8
XFILLER_15_483 VDD VSS sg13g2_decap_8
XFILLER_8_42 VDD VSS sg13g2_decap_8
XFILLER_30_497 VDD VSS sg13g2_decap_8
XFILLER_7_693 VDD VSS sg13g2_decap_8
XFILLER_69_133 VDD VSS sg13g2_decap_8
XFILLER_33_0 VDD VSS sg13g2_decap_8
XFILLER_85_637 VDD VSS sg13g2_decap_8
XFILLER_84_147 VDD VSS sg13g2_decap_8
XFILLER_65_350 VDD VSS sg13g2_decap_8
XFILLER_38_553 VDD VSS sg13g2_decap_8
XFILLER_25_203 VDD VSS sg13g2_decap_8
XFILLER_26_748 VDD VSS sg13g2_decap_8
XFILLER_53_567 VDD VSS sg13g2_decap_8
XFILLER_41_707 VDD VSS sg13g2_decap_8
XFILLER_80_364 VDD VSS sg13g2_decap_8
XFILLER_43_28 VDD VSS sg13g2_decap_8
XFILLER_40_217 VDD VSS sg13g2_decap_8
XFILLER_21_420 VDD VSS sg13g2_decap_8
XFILLER_33_280 VDD VSS sg13g2_decap_8
XFILLER_21_497 VDD VSS sg13g2_decap_8
XFILLER_68_14 VDD VSS sg13g2_decap_8
XFILLER_88_420 VDD VSS sg13g2_decap_8
XFILLER_76_615 VDD VSS sg13g2_decap_8
XFILLER_0_357 VDD VSS sg13g2_decap_8
XFILLER_88_497 VDD VSS sg13g2_decap_8
XFILLER_75_158 VDD VSS sg13g2_decap_8
XFILLER_84_35 VDD VSS sg13g2_decap_8
XFILLER_56_350 VDD VSS sg13g2_decap_8
XFILLER_29_553 VDD VSS sg13g2_decap_8
XFILLER_16_203 VDD VSS sg13g2_decap_8
XFILLER_71_331 VDD VSS sg13g2_decap_8
XFILLER_32_707 VDD VSS sg13g2_decap_8
XFILLER_17_84 VDD VSS sg13g2_decap_8
XFILLER_31_217 VDD VSS sg13g2_decap_8
XFILLER_44_567 VDD VSS sg13g2_decap_8
XFILLER_12_420 VDD VSS sg13g2_decap_8
XFILLER_24_280 VDD VSS sg13g2_decap_8
XFILLER_8_413 VDD VSS sg13g2_decap_8
XFILLER_12_497 VDD VSS sg13g2_decap_8
X_82__5 VDD VSS _82__5/L_HI sg13g2_tiehi
XFILLER_4_630 VDD VSS sg13g2_decap_8
XFILLER_3_140 VDD VSS sg13g2_decap_8
XFILLER_79_420 VDD VSS sg13g2_decap_8
XFILLER_67_604 VDD VSS sg13g2_decap_8
XFILLER_79_497 VDD VSS sg13g2_decap_8
XFILLER_94_434 VDD VSS sg13g2_decap_8
XFILLER_58_91 VDD VSS sg13g2_decap_8
XFILLER_66_147 VDD VSS sg13g2_decap_8
XFILLER_47_350 VDD VSS sg13g2_decap_8
XFILLER_90_651 VDD VSS sg13g2_decap_8
XFILLER_62_364 VDD VSS sg13g2_decap_8
XFILLER_50_504 VDD VSS sg13g2_decap_8
XFILLER_23_707 VDD VSS sg13g2_decap_8
XFILLER_35_567 VDD VSS sg13g2_decap_8
XFILLER_15_280 VDD VSS sg13g2_decap_8
XFILLER_22_217 VDD VSS sg13g2_decap_8
XFILLER_30_294 VDD VSS sg13g2_decap_8
XFILLER_7_490 VDD VSS sg13g2_decap_8
XFILLER_89_217 VDD VSS sg13g2_decap_8
XFILLER_85_434 VDD VSS sg13g2_decap_8
XFILLER_58_637 VDD VSS sg13g2_decap_8
XFILLER_38_28 VDD VSS sg13g2_decap_8
XFILLER_73_618 VDD VSS sg13g2_decap_8
XFILLER_57_147 VDD VSS sg13g2_decap_8
XFILLER_66_681 VDD VSS sg13g2_decap_8
XFILLER_38_350 VDD VSS sg13g2_decap_8
XFILLER_81_651 VDD VSS sg13g2_decap_8
XFILLER_26_545 VDD VSS sg13g2_decap_8
XFILLER_80_161 VDD VSS sg13g2_decap_8
XFILLER_54_49 VDD VSS sg13g2_decap_8
XFILLER_53_364 VDD VSS sg13g2_decap_8
XFILLER_14_707 VDD VSS sg13g2_decap_8
XFILLER_41_504 VDD VSS sg13g2_decap_8
XFILLER_13_217 VDD VSS sg13g2_decap_8
XFILLER_21_294 VDD VSS sg13g2_decap_8
XFILLER_5_427 VDD VSS sg13g2_decap_8
XFILLER_79_35 VDD VSS sg13g2_decap_8
XFILLER_1_644 VDD VSS sg13g2_decap_8
XFILLER_0_154 VDD VSS sg13g2_decap_8
XFILLER_88_294 VDD VSS sg13g2_decap_8
XFILLER_76_412 VDD VSS sg13g2_decap_8
XFILLER_95_56 VDD VSS sg13g2_decap_8
XFILLER_49_637 VDD VSS sg13g2_decap_8
XFILLER_48_147 VDD VSS sg13g2_decap_8
XFILLER_76_489 VDD VSS sg13g2_decap_8
XFILLER_29_350 VDD VSS sg13g2_decap_8
XFILLER_91_448 VDD VSS sg13g2_decap_8
XFILLER_72_684 VDD VSS sg13g2_decap_8
XFILLER_44_364 VDD VSS sg13g2_decap_8
XFILLER_17_567 VDD VSS sg13g2_decap_8
XFILLER_32_504 VDD VSS sg13g2_decap_8
XFILLER_71_161 VDD VSS sg13g2_decap_8
XFILLER_9_700 VDD VSS sg13g2_decap_8
XFILLER_8_210 VDD VSS sg13g2_decap_8
XFILLER_40_581 VDD VSS sg13g2_decap_8
XFILLER_74_7 VDD VSS sg13g2_decap_8
XFILLER_12_294 VDD VSS sg13g2_decap_8
XFILLER_8_287 VDD VSS sg13g2_decap_8
XFILLER_60_70 VDD VSS sg13g2_decap_8
XFILLER_5_21 VDD VSS sg13g2_decap_8
XFILLER_5_98 VDD VSS sg13g2_decap_8
XFILLER_67_401 VDD VSS sg13g2_decap_8
XFILLER_95_721 VDD VSS sg13g2_decap_8
XFILLER_79_294 VDD VSS sg13g2_decap_8
XFILLER_94_231 VDD VSS sg13g2_decap_8
XFILLER_39_147 VDD VSS sg13g2_decap_8
XFILLER_67_478 VDD VSS sg13g2_decap_8
XFILLER_82_448 VDD VSS sg13g2_decap_8
XFILLER_63_662 VDD VSS sg13g2_decap_8
XFILLER_35_364 VDD VSS sg13g2_decap_8
XFILLER_23_504 VDD VSS sg13g2_decap_8
XFILLER_62_161 VDD VSS sg13g2_decap_8
XFILLER_50_301 VDD VSS sg13g2_decap_8
XFILLER_50_378 VDD VSS sg13g2_decap_8
XFILLER_31_581 VDD VSS sg13g2_decap_8
XFILLER_49_49 VDD VSS sg13g2_decap_8
XFILLER_86_721 VDD VSS sg13g2_decap_8
XFILLER_58_434 VDD VSS sg13g2_decap_8
XFILLER_85_231 VDD VSS sg13g2_decap_8
XFILLER_54_651 VDD VSS sg13g2_decap_8
XFILLER_26_342 VDD VSS sg13g2_decap_8
XFILLER_14_504 VDD VSS sg13g2_decap_8
XFILLER_81_14 VDD VSS sg13g2_decap_8
XFILLER_41_301 VDD VSS sg13g2_decap_8
XFILLER_53_161 VDD VSS sg13g2_decap_8
XFILLER_14_63 VDD VSS sg13g2_decap_8
XFILLER_41_378 VDD VSS sg13g2_decap_8
XFILLER_10_721 VDD VSS sg13g2_decap_8
XFILLER_22_581 VDD VSS sg13g2_decap_8
XFILLER_6_714 VDD VSS sg13g2_decap_8
XFILLER_5_224 VDD VSS sg13g2_decap_8
XFILLER_30_84 VDD VSS sg13g2_decap_8
XFILLER_68_209 VDD VSS sg13g2_decap_8
XFILLER_1_441 VDD VSS sg13g2_decap_8
XFILLER_89_581 VDD VSS sg13g2_decap_8
X_70_ VSS VDD _74_/C _74_/D _70_/Y _69_/Y sg13g2_a21oi_1
XFILLER_49_434 VDD VSS sg13g2_decap_8
XFILLER_92_735 VDD VSS sg13g2_decap_8
XFILLER_76_264 VDD VSS sg13g2_decap_8
XFILLER_91_245 VDD VSS sg13g2_decap_8
XFILLER_64_448 VDD VSS sg13g2_decap_8
XFILLER_55_70 VDD VSS sg13g2_decap_8
XFILLER_17_364 VDD VSS sg13g2_decap_8
XFILLER_45_651 VDD VSS sg13g2_decap_8
XFILLER_72_481 VDD VSS sg13g2_decap_8
XFILLER_32_301 VDD VSS sg13g2_decap_8
XFILLER_44_161 VDD VSS sg13g2_decap_8
XFILLER_60_665 VDD VSS sg13g2_decap_8
XFILLER_32_378 VDD VSS sg13g2_decap_8
XFILLER_20_518 VDD VSS sg13g2_decap_8
XFILLER_71_91 VDD VSS sg13g2_decap_8
XFILLER_13_581 VDD VSS sg13g2_decap_8
XFILLER_9_574 VDD VSS sg13g2_decap_8
XFILLER_87_518 VDD VSS sg13g2_decap_8
XFILLER_67_275 VDD VSS sg13g2_decap_8
XFILLER_95_595 VDD VSS sg13g2_decap_8
XFILLER_83_735 VDD VSS sg13g2_decap_8
XFILLER_55_448 VDD VSS sg13g2_decap_8
XFILLER_82_245 VDD VSS sg13g2_decap_8
XFILLER_70_418 VDD VSS sg13g2_decap_8
XFILLER_36_651 VDD VSS sg13g2_decap_8
XFILLER_23_301 VDD VSS sg13g2_decap_8
XFILLER_35_161 VDD VSS sg13g2_decap_8
XFILLER_51_665 VDD VSS sg13g2_decap_8
XFILLER_11_518 VDD VSS sg13g2_decap_8
XFILLER_23_378 VDD VSS sg13g2_decap_8
XFILLER_50_175 VDD VSS sg13g2_decap_8
XFILLER_51_28 VDD VSS sg13g2_decap_8
XFILLER_3_728 VDD VSS sg13g2_decap_8
XFILLER_4_7 VDD VSS sg13g2_decap_8
XFILLER_2_238 VDD VSS sg13g2_decap_8
XFILLER_78_518 VDD VSS sg13g2_decap_8
XFILLER_76_14 VDD VSS sg13g2_decap_8
XFILLER_59_721 VDD VSS sg13g2_decap_8
XFILLER_58_231 VDD VSS sg13g2_decap_8
XFILLER_86_595 VDD VSS sg13g2_decap_8
XFILLER_74_735 VDD VSS sg13g2_decap_8
XFILLER_46_448 VDD VSS sg13g2_decap_8
XFILLER_73_245 VDD VSS sg13g2_decap_8
XFILLER_92_35 VDD VSS sg13g2_decap_8
XFILLER_27_651 VDD VSS sg13g2_decap_8
XFILLER_14_301 VDD VSS sg13g2_decap_8
XFILLER_26_161 VDD VSS sg13g2_decap_8
XFILLER_42_665 VDD VSS sg13g2_decap_8
XFILLER_25_84 VDD VSS sg13g2_decap_8
XFILLER_14_378 VDD VSS sg13g2_decap_8
XFILLER_41_175 VDD VSS sg13g2_decap_8
XFILLER_6_511 VDD VSS sg13g2_decap_8
XFILLER_10_595 VDD VSS sg13g2_decap_8
XFILLER_6_588 VDD VSS sg13g2_decap_8
XFILLER_37_7 VDD VSS sg13g2_decap_8
XFILLER_49_231 VDD VSS sg13g2_decap_8
XFILLER_77_562 VDD VSS sg13g2_decap_8
XFILLER_65_724 VDD VSS sg13g2_decap_8
X_53_ _75_/A VDD _53_/Y VSS _76_/Q _55_/A2 sg13g2_o21ai_1
XFILLER_2_77 VDD VSS sg13g2_decap_8
XFILLER_92_532 VDD VSS sg13g2_decap_8
XFILLER_37_448 VDD VSS sg13g2_decap_8
XFILLER_64_245 VDD VSS sg13g2_decap_8
XFILLER_66_91 VDD VSS sg13g2_decap_8
XFILLER_18_651 VDD VSS sg13g2_decap_8
XFILLER_80_749 VDD VSS sg13g2_decap_8
XFILLER_17_161 VDD VSS sg13g2_decap_8
XFILLER_33_665 VDD VSS sg13g2_decap_8
XFILLER_20_315 VDD VSS sg13g2_decap_8
XFILLER_60_462 VDD VSS sg13g2_decap_8
XFILLER_32_175 VDD VSS sg13g2_decap_8
XFILLER_9_371 VDD VSS sg13g2_decap_8
XFILLER_63_0 VDD VSS sg13g2_decap_8
XFILLER_87_315 VDD VSS sg13g2_decap_8
XFILLER_68_573 VDD VSS sg13g2_decap_8
XFILLER_83_532 VDD VSS sg13g2_decap_8
XFILLER_95_392 VDD VSS sg13g2_decap_8
XFILLER_56_735 VDD VSS sg13g2_decap_8
XFILLER_46_28 VDD VSS sg13g2_decap_8
XFILLER_28_448 VDD VSS sg13g2_decap_8
XFILLER_71_716 VDD VSS sg13g2_decap_8
XFILLER_55_245 VDD VSS sg13g2_decap_8
XFILLER_62_49 VDD VSS sg13g2_decap_8
XFILLER_51_462 VDD VSS sg13g2_decap_8
XFILLER_24_665 VDD VSS sg13g2_decap_8
XFILLER_11_315 VDD VSS sg13g2_decap_8
XFILLER_23_175 VDD VSS sg13g2_decap_8
XFILLER_7_308 VDD VSS sg13g2_decap_8
XFILLER_11_42 VDD VSS sg13g2_decap_8
XFILLER_3_525 VDD VSS sg13g2_decap_8
XFILLER_78_315 VDD VSS sg13g2_decap_8
XFILLER_87_35 VDD VSS sg13g2_decap_8
XFILLER_93_329 VDD VSS sg13g2_decap_8
XFILLER_74_532 VDD VSS sg13g2_decap_8
XFILLER_86_392 VDD VSS sg13g2_decap_8
XFILLER_59_595 VDD VSS sg13g2_decap_8
XFILLER_47_735 VDD VSS sg13g2_decap_8
XFILLER_19_448 VDD VSS sg13g2_decap_8
XFILLER_46_245 VDD VSS sg13g2_decap_8
XFILLER_62_749 VDD VSS sg13g2_decap_8
XFILLER_61_259 VDD VSS sg13g2_decap_8
XFILLER_42_462 VDD VSS sg13g2_decap_8
XFILLER_15_665 VDD VSS sg13g2_decap_8
XFILLER_30_602 VDD VSS sg13g2_decap_8
XFILLER_14_175 VDD VSS sg13g2_decap_8
XFILLER_30_679 VDD VSS sg13g2_decap_8
XFILLER_10_392 VDD VSS sg13g2_decap_8
XFILLER_6_385 VDD VSS sg13g2_decap_8
XFILLER_69_359 VDD VSS sg13g2_decap_8
XFILLER_65_521 VDD VSS sg13g2_decap_8
XFILLER_84_329 VDD VSS sg13g2_decap_8
XFILLER_38_735 VDD VSS sg13g2_decap_8
XFILLER_37_245 VDD VSS sg13g2_decap_8
XFILLER_65_598 VDD VSS sg13g2_decap_8
XFILLER_53_749 VDD VSS sg13g2_decap_8
XFILLER_80_546 VDD VSS sg13g2_decap_8
XFILLER_52_259 VDD VSS sg13g2_decap_8
XFILLER_33_462 VDD VSS sg13g2_decap_8
XFILLER_21_602 VDD VSS sg13g2_decap_8
XFILLER_20_112 VDD VSS sg13g2_decap_8
XFILLER_21_679 VDD VSS sg13g2_decap_8
XFILLER_20_189 VDD VSS sg13g2_decap_8
XFILLER_88_602 VDD VSS sg13g2_decap_8
XFILLER_87_112 VDD VSS sg13g2_decap_8
XFILLER_0_539 VDD VSS sg13g2_decap_8
XFILLER_88_679 VDD VSS sg13g2_decap_8
XFILLER_57_49 VDD VSS sg13g2_decap_8
XFILLER_87_189 VDD VSS sg13g2_decap_8
XFILLER_68_370 VDD VSS sg13g2_decap_8
XFILLER_56_532 VDD VSS sg13g2_decap_8
XFILLER_29_735 VDD VSS sg13g2_decap_8
XFILLER_28_245 VDD VSS sg13g2_decap_8
XFILLER_71_513 VDD VSS sg13g2_decap_8
XFILLER_44_749 VDD VSS sg13g2_decap_8
XFILLER_43_259 VDD VSS sg13g2_decap_8
XFILLER_12_602 VDD VSS sg13g2_decap_8
XFILLER_24_462 VDD VSS sg13g2_decap_8
XFILLER_11_112 VDD VSS sg13g2_decap_8
XFILLER_12_679 VDD VSS sg13g2_decap_8
XFILLER_7_105 VDD VSS sg13g2_decap_8
XFILLER_11_189 VDD VSS sg13g2_decap_8
XFILLER_22_63 VDD VSS sg13g2_decap_8
XFILLER_3_322 VDD VSS sg13g2_decap_8
XFILLER_79_602 VDD VSS sg13g2_decap_8
XFILLER_78_112 VDD VSS sg13g2_decap_8
XFILLER_3_399 VDD VSS sg13g2_decap_8
XFILLER_94_616 VDD VSS sg13g2_decap_8
XFILLER_79_679 VDD VSS sg13g2_decap_8
XFILLER_93_126 VDD VSS sg13g2_decap_8
XFILLER_78_189 VDD VSS sg13g2_decap_8
XFILLER_66_329 VDD VSS sg13g2_decap_8
XFILLER_47_532 VDD VSS sg13g2_decap_8
XFILLER_59_392 VDD VSS sg13g2_decap_8
XFILLER_19_245 VDD VSS sg13g2_decap_8
XFILLER_62_546 VDD VSS sg13g2_decap_8
XFILLER_74_395 VDD VSS sg13g2_decap_8
XFILLER_35_749 VDD VSS sg13g2_decap_8
XFILLER_63_70 VDD VSS sg13g2_decap_8
XFILLER_15_462 VDD VSS sg13g2_decap_8
XFILLER_34_259 VDD VSS sg13g2_decap_8
XFILLER_8_21 VDD VSS sg13g2_decap_8
XFILLER_30_476 VDD VSS sg13g2_decap_8
XFILLER_8_98 VDD VSS sg13g2_decap_8
XFILLER_7_672 VDD VSS sg13g2_decap_8
XFILLER_6_182 VDD VSS sg13g2_decap_8
XFILLER_69_112 VDD VSS sg13g2_decap_8
XFILLER_85_616 VDD VSS sg13g2_decap_8
XFILLER_26_0 VDD VSS sg13g2_decap_8
XFILLER_84_126 VDD VSS sg13g2_decap_8
XFILLER_69_189 VDD VSS sg13g2_decap_8
XFILLER_57_329 VDD VSS sg13g2_decap_8
XFILLER_38_532 VDD VSS sg13g2_decap_8
XFILLER_93_693 VDD VSS sg13g2_decap_8
XFILLER_26_727 VDD VSS sg13g2_decap_8
XFILLER_80_343 VDD VSS sg13g2_decap_8
XFILLER_53_546 VDD VSS sg13g2_decap_8
XFILLER_25_259 VDD VSS sg13g2_decap_8
XFILLER_21_476 VDD VSS sg13g2_decap_8
XFILLER_5_609 VDD VSS sg13g2_decap_8
XFILLER_4_119 VDD VSS sg13g2_decap_8
XFILLER_0_336 VDD VSS sg13g2_decap_8
XFILLER_88_476 VDD VSS sg13g2_decap_8
XFILLER_48_329 VDD VSS sg13g2_decap_8
XFILLER_75_137 VDD VSS sg13g2_decap_8
XFILLER_84_14 VDD VSS sg13g2_decap_8
XFILLER_29_532 VDD VSS sg13g2_decap_8
XFILLER_84_693 VDD VSS sg13g2_decap_8
XFILLER_17_63 VDD VSS sg13g2_decap_8
XFILLER_17_749 VDD VSS sg13g2_decap_8
XFILLER_44_546 VDD VSS sg13g2_decap_8
XFILLER_16_259 VDD VSS sg13g2_decap_8
XFILLER_71_387 VDD VSS sg13g2_decap_8
XFILLER_12_476 VDD VSS sg13g2_decap_8
XFILLER_33_84 VDD VSS sg13g2_decap_8
XFILLER_8_469 VDD VSS sg13g2_decap_8
XFILLER_4_686 VDD VSS sg13g2_decap_8
XFILLER_3_196 VDD VSS sg13g2_decap_8
XFILLER_79_476 VDD VSS sg13g2_decap_8
XFILLER_94_413 VDD VSS sg13g2_decap_8
XFILLER_66_126 VDD VSS sg13g2_decap_8
XFILLER_58_70 VDD VSS sg13g2_decap_8
XFILLER_39_329 VDD VSS sg13g2_decap_8
XFILLER_90_630 VDD VSS sg13g2_decap_8
XFILLER_35_546 VDD VSS sg13g2_decap_8
XFILLER_62_343 VDD VSS sg13g2_decap_8
XFILLER_74_91 VDD VSS sg13g2_decap_8
XFILLER_30_273 VDD VSS sg13g2_decap_8
XFILLER_58_616 VDD VSS sg13g2_decap_8
XFILLER_85_413 VDD VSS sg13g2_decap_8
XFILLER_57_126 VDD VSS sg13g2_decap_8
XFILLER_66_660 VDD VSS sg13g2_decap_8
XFILLER_93_490 VDD VSS sg13g2_decap_8
XFILLER_81_630 VDD VSS sg13g2_decap_8
XFILLER_54_28 VDD VSS sg13g2_decap_8
XFILLER_26_524 VDD VSS sg13g2_decap_8
XFILLER_80_140 VDD VSS sg13g2_decap_8
XFILLER_53_343 VDD VSS sg13g2_decap_8
XFILLER_70_49 VDD VSS sg13g2_decap_8
XFILLER_21_273 VDD VSS sg13g2_decap_8
XFILLER_5_406 VDD VSS sg13g2_decap_8
XFILLER_79_14 VDD VSS sg13g2_decap_8
XFILLER_1_623 VDD VSS sg13g2_decap_8
XFILLER_49_616 VDD VSS sg13g2_decap_8
XFILLER_0_133 VDD VSS sg13g2_decap_8
XFILLER_88_273 VDD VSS sg13g2_decap_8
XFILLER_95_35 VDD VSS sg13g2_decap_8
XFILLER_48_126 VDD VSS sg13g2_decap_8
XFILLER_91_427 VDD VSS sg13g2_decap_8
XFILLER_28_84 VDD VSS sg13g2_decap_8
XFILLER_84_490 VDD VSS sg13g2_decap_8
XFILLER_57_693 VDD VSS sg13g2_decap_8
XFILLER_17_546 VDD VSS sg13g2_decap_8
XFILLER_72_663 VDD VSS sg13g2_decap_8
XFILLER_71_140 VDD VSS sg13g2_decap_8
XFILLER_44_343 VDD VSS sg13g2_decap_8
XFILLER_40_560 VDD VSS sg13g2_decap_8
XFILLER_9_756 VDD VSS sg13g2_fill_1
XFILLER_12_273 VDD VSS sg13g2_decap_8
XIO_BOND_outputs\[2\].output_pad output_PAD[2] bondpad_70x70_novias
XFILLER_67_7 VDD VSS sg13g2_decap_8
XFILLER_8_266 VDD VSS sg13g2_decap_8
XFILLER_4_483 VDD VSS sg13g2_decap_8
XFILLER_5_77 VDD VSS sg13g2_decap_8
XFILLER_95_700 VDD VSS sg13g2_decap_8
XFILLER_69_91 VDD VSS sg13g2_decap_8
XFILLER_94_210 VDD VSS sg13g2_decap_8
XFILLER_79_273 VDD VSS sg13g2_decap_8
XFILLER_67_457 VDD VSS sg13g2_decap_8
XFILLER_39_126 VDD VSS sg13g2_decap_8
XFILLER_94_287 VDD VSS sg13g2_decap_8
XFILLER_82_427 VDD VSS sg13g2_decap_8
XFILLER_63_641 VDD VSS sg13g2_decap_8
XFILLER_48_693 VDD VSS sg13g2_decap_8
XFILLER_62_140 VDD VSS sg13g2_decap_8
XFILLER_35_343 VDD VSS sg13g2_decap_8
XFILLER_93_0 VDD VSS sg13g2_decap_8
XFILLER_50_357 VDD VSS sg13g2_decap_8
XFILLER_31_560 VDD VSS sg13g2_decap_8
XFILLER_49_28 VDD VSS sg13g2_decap_8
XFILLER_86_700 VDD VSS sg13g2_decap_8
XFILLER_85_210 VDD VSS sg13g2_decap_8
XFILLER_58_413 VDD VSS sg13g2_decap_8
XFILLER_65_49 VDD VSS sg13g2_decap_8
XFILLER_85_287 VDD VSS sg13g2_decap_8
XFILLER_73_449 VDD VSS sg13g2_fill_2
XFILLER_54_630 VDD VSS sg13g2_decap_8
XFILLER_26_321 VDD VSS sg13g2_decap_8
XFILLER_39_693 VDD VSS sg13g2_decap_8
XFILLER_53_140 VDD VSS sg13g2_decap_8
XFILLER_26_398 VDD VSS sg13g2_decap_8
XFILLER_41_357 VDD VSS sg13g2_decap_8
XFILLER_10_700 VDD VSS sg13g2_decap_8
XFILLER_14_42 VDD VSS sg13g2_decap_8
XFILLER_22_560 VDD VSS sg13g2_decap_8
XFILLER_5_203 VDD VSS sg13g2_decap_8
XFILLER_30_63 VDD VSS sg13g2_decap_8
XFILLER_1_420 VDD VSS sg13g2_decap_8
XFILLER_89_560 VDD VSS sg13g2_decap_8
XFILLER_49_413 VDD VSS sg13g2_decap_8
XFILLER_77_755 VDD VSS sg13g2_fill_2
XFILLER_77_744 VDD VSS sg13g2_decap_8
XFILLER_76_243 VDD VSS sg13g2_decap_8
XFILLER_76_210 VDD VSS sg13g2_decap_8
XFILLER_1_497 VDD VSS sg13g2_decap_8
XFILLER_92_714 VDD VSS sg13g2_decap_8
XFILLER_91_224 VDD VSS sg13g2_decap_8
XFILLER_64_427 VDD VSS sg13g2_decap_8
XFILLER_57_490 VDD VSS sg13g2_decap_8
XFILLER_45_630 VDD VSS sg13g2_decap_8
XFILLER_17_343 VDD VSS sg13g2_decap_8
XFILLER_44_140 VDD VSS sg13g2_decap_8
XFILLER_72_460 VDD VSS sg13g2_decap_8
XFILLER_60_644 VDD VSS sg13g2_decap_8
XFILLER_32_357 VDD VSS sg13g2_decap_8
XFILLER_13_560 VDD VSS sg13g2_decap_8
XFILLER_71_70 VDD VSS sg13g2_decap_8
XFILLER_9_553 VDD VSS sg13g2_decap_8
XFILLER_4_280 VDD VSS sg13g2_decap_8
XFILLER_68_755 VDD VSS sg13g2_fill_2
XFILLER_95_574 VDD VSS sg13g2_decap_8
XFILLER_83_714 VDD VSS sg13g2_decap_8
XFILLER_67_254 VDD VSS sg13g2_decap_8
XFILLER_82_224 VDD VSS sg13g2_decap_8
XFILLER_48_490 VDD VSS sg13g2_decap_8
XFILLER_55_427 VDD VSS sg13g2_decap_8
XFILLER_36_630 VDD VSS sg13g2_decap_8
XFILLER_35_140 VDD VSS sg13g2_decap_8
XFILLER_51_644 VDD VSS sg13g2_decap_8
XFILLER_23_357 VDD VSS sg13g2_decap_8
XFILLER_50_154 VDD VSS sg13g2_decap_8
XFILLER_3_707 VDD VSS sg13g2_decap_8
XFILLER_2_217 VDD VSS sg13g2_decap_8
XFILLER_59_700 VDD VSS sg13g2_decap_8
XFILLER_58_210 VDD VSS sg13g2_decap_8
XFILLER_86_574 VDD VSS sg13g2_decap_8
XFILLER_74_714 VDD VSS sg13g2_decap_8
XFILLER_73_224 VDD VSS sg13g2_decap_8
XFILLER_46_427 VDD VSS sg13g2_decap_8
XFILLER_58_287 VDD VSS sg13g2_decap_8
XFILLER_27_630 VDD VSS sg13g2_decap_8
XFILLER_73_268 VDD VSS sg13g2_decap_4
XFILLER_92_14 VDD VSS sg13g2_decap_8
XFILLER_26_140 VDD VSS sg13g2_decap_8
XFILLER_39_490 VDD VSS sg13g2_decap_8
XFILLER_25_63 VDD VSS sg13g2_decap_8
XFILLER_42_644 VDD VSS sg13g2_decap_8
XFILLER_14_357 VDD VSS sg13g2_decap_8
XFILLER_41_154 VDD VSS sg13g2_decap_8
XFILLER_10_574 VDD VSS sg13g2_decap_8
XFILLER_41_84 VDD VSS sg13g2_decap_8
XFILLER_6_567 VDD VSS sg13g2_decap_8
XFILLER_77_541 VDD VSS sg13g2_decap_8
XFILLER_1_294 VDD VSS sg13g2_decap_8
XFILLER_49_210 VDD VSS sg13g2_decap_8
XFILLER_65_703 VDD VSS sg13g2_decap_8
X_52_ _52_/B _52_/C _52_/A _52_/Y VDD VSS _52_/D sg13g2_nand4_1
XFILLER_2_56 VDD VSS sg13g2_decap_8
XFILLER_92_511 VDD VSS sg13g2_decap_8
XFILLER_64_224 VDD VSS sg13g2_decap_8
XFILLER_66_70 VDD VSS sg13g2_decap_8
XFILLER_37_427 VDD VSS sg13g2_decap_8
XFILLER_49_287 VDD VSS sg13g2_decap_8
XFILLER_18_630 VDD VSS sg13g2_decap_8
XFILLER_92_588 VDD VSS sg13g2_decap_8
XFILLER_80_728 VDD VSS sg13g2_decap_8
XFILLER_17_140 VDD VSS sg13g2_decap_8
XFILLER_60_441 VDD VSS sg13g2_decap_8
XFILLER_33_644 VDD VSS sg13g2_decap_8
XFILLER_82_91 VDD VSS sg13g2_decap_8
XFILLER_32_154 VDD VSS sg13g2_decap_8
XFILLER_9_350 VDD VSS sg13g2_decap_8
XFILLER_56_0 VDD VSS sg13g2_decap_8
XFILLER_68_552 VDD VSS sg13g2_decap_8
XFILLER_56_714 VDD VSS sg13g2_decap_8
XFILLER_83_511 VDD VSS sg13g2_decap_8
XFILLER_95_371 VDD VSS sg13g2_decap_8
XFILLER_28_427 VDD VSS sg13g2_decap_8
XFILLER_55_224 VDD VSS sg13g2_decap_8
XFILLER_83_588 VDD VSS sg13g2_decap_8
XFILLER_70_249 VDD VSS sg13g2_decap_8
XFILLER_62_28 VDD VSS sg13g2_decap_8
XFILLER_24_644 VDD VSS sg13g2_decap_8
XFILLER_23_154 VDD VSS sg13g2_decap_8
XFILLER_51_441 VDD VSS sg13g2_decap_8
XFILLER_11_21 VDD VSS sg13g2_decap_8
XFILLER_3_504 VDD VSS sg13g2_decap_8
XFILLER_87_14 VDD VSS sg13g2_decap_8
XFILLER_11_98 VDD VSS sg13g2_decap_8
XFILLER_93_308 VDD VSS sg13g2_decap_8
XFILLER_59_574 VDD VSS sg13g2_decap_8
XFILLER_47_714 VDD VSS sg13g2_decap_8
XFILLER_74_511 VDD VSS sg13g2_decap_8
XFILLER_86_371 VDD VSS sg13g2_decap_8
XFILLER_19_427 VDD VSS sg13g2_decap_8
XFILLER_46_224 VDD VSS sg13g2_decap_8
XFILLER_74_588 VDD VSS sg13g2_decap_8
XFILLER_62_728 VDD VSS sg13g2_decap_8
XFILLER_36_84 VDD VSS sg13g2_decap_8
XFILLER_61_238 VDD VSS sg13g2_decap_8
XFILLER_15_644 VDD VSS sg13g2_decap_8
XFILLER_70_750 VDD VSS sg13g2_decap_8
Xinputs\[7\].input_pad IOVDD IOVSS _52_/D input_PAD[7] VDD VSS sg13g2_IOPadIn
XFILLER_14_154 VDD VSS sg13g2_decap_8
XFILLER_42_441 VDD VSS sg13g2_decap_8
XFILLER_30_658 VDD VSS sg13g2_decap_8
XFILLER_10_371 VDD VSS sg13g2_decap_8
XFILLER_6_364 VDD VSS sg13g2_decap_8
XFILLER_69_338 VDD VSS sg13g2_decap_8
XFILLER_2_581 VDD VSS sg13g2_decap_8
XFILLER_84_308 VDD VSS sg13g2_decap_8
XFILLER_77_91 VDD VSS sg13g2_decap_8
XFILLER_38_714 VDD VSS sg13g2_decap_8
XFILLER_65_500 VDD VSS sg13g2_decap_8
XFILLER_77_393 VDD VSS sg13g2_fill_1
XFILLER_37_224 VDD VSS sg13g2_decap_8
XFILLER_80_525 VDD VSS sg13g2_decap_8
XFILLER_65_577 VDD VSS sg13g2_decap_8
XFILLER_92_385 VDD VSS sg13g2_decap_8
XFILLER_53_728 VDD VSS sg13g2_decap_8
XFILLER_52_238 VDD VSS sg13g2_decap_8
XFILLER_33_441 VDD VSS sg13g2_decap_8
XFILLER_21_658 VDD VSS sg13g2_decap_8
XFILLER_20_168 VDD VSS sg13g2_decap_8
XFILLER_0_518 VDD VSS sg13g2_decap_8
XFILLER_88_658 VDD VSS sg13g2_decap_8
XFILLER_87_168 VDD VSS sg13g2_decap_8
XFILLER_57_28 VDD VSS sg13g2_decap_8
XFILLER_56_511 VDD VSS sg13g2_decap_8
XFILLER_29_714 VDD VSS sg13g2_decap_8
XFILLER_28_224 VDD VSS sg13g2_decap_8
XFILLER_83_385 VDD VSS sg13g2_decap_8
XFILLER_56_588 VDD VSS sg13g2_decap_8
XFILLER_44_728 VDD VSS sg13g2_decap_8
XFILLER_73_49 VDD VSS sg13g2_decap_8
XFILLER_43_238 VDD VSS sg13g2_decap_8
XFILLER_71_569 VDD VSS sg13g2_decap_8
XFILLER_24_441 VDD VSS sg13g2_decap_8
XFILLER_12_658 VDD VSS sg13g2_decap_8
XFILLER_11_168 VDD VSS sg13g2_decap_8
XFILLER_22_42 VDD VSS sg13g2_decap_8
XFILLER_3_301 VDD VSS sg13g2_decap_8
XIO_BOND_outputs\[7\].output_pad output_PAD[7] bondpad_70x70_novias
XFILLER_3_378 VDD VSS sg13g2_decap_8
XFILLER_79_658 VDD VSS sg13g2_decap_8
XFILLER_78_168 VDD VSS sg13g2_decap_8
XFILLER_66_308 VDD VSS sg13g2_decap_8
XFILLER_93_105 VDD VSS sg13g2_decap_8
XFILLER_47_511 VDD VSS sg13g2_decap_8
XFILLER_59_371 VDD VSS sg13g2_decap_8
XFILLER_74_330 VDD VSS sg13g2_decap_8
XFILLER_19_224 VDD VSS sg13g2_decap_8
XFILLER_62_525 VDD VSS sg13g2_decap_8
XFILLER_47_588 VDD VSS sg13g2_decap_8
XFILLER_35_728 VDD VSS sg13g2_decap_8
XFILLER_34_238 VDD VSS sg13g2_decap_8
XFILLER_15_441 VDD VSS sg13g2_decap_8
XFILLER_30_455 VDD VSS sg13g2_decap_8
XFILLER_7_651 VDD VSS sg13g2_decap_8
XFILLER_8_77 VDD VSS sg13g2_decap_8
XFILLER_6_161 VDD VSS sg13g2_decap_8
XFILLER_69_168 VDD VSS sg13g2_decap_8
XFILLER_57_308 VDD VSS sg13g2_decap_8
XFILLER_84_105 VDD VSS sg13g2_decap_8
XFILLER_38_511 VDD VSS sg13g2_decap_8
XFILLER_19_0 VDD VSS sg13g2_decap_8
XFILLER_93_672 VDD VSS sg13g2_decap_8
XFILLER_26_706 VDD VSS sg13g2_decap_8
XFILLER_38_588 VDD VSS sg13g2_decap_8
XFILLER_92_182 VDD VSS sg13g2_decap_8
XFILLER_80_322 VDD VSS sg13g2_decap_8
XFILLER_65_385 VDD VSS sg13g2_decap_8
XFILLER_53_525 VDD VSS sg13g2_decap_8
XFILLER_25_238 VDD VSS sg13g2_decap_8
XFILLER_80_399 VDD VSS sg13g2_decap_8
XFILLER_21_455 VDD VSS sg13g2_decap_8
XFILLER_68_49 VDD VSS sg13g2_decap_8
XFILLER_0_315 VDD VSS sg13g2_decap_8
XFILLER_88_455 VDD VSS sg13g2_decap_8
XFILLER_48_308 VDD VSS sg13g2_decap_8
XFILLER_75_116 VDD VSS sg13g2_decap_8
XFILLER_29_511 VDD VSS sg13g2_decap_8
XFILLER_91_609 VDD VSS sg13g2_decap_8
XFILLER_84_672 VDD VSS sg13g2_decap_8
XFILLER_90_119 VDD VSS sg13g2_decap_8
XFILLER_17_728 VDD VSS sg13g2_decap_8
XFILLER_29_588 VDD VSS sg13g2_decap_8
XFILLER_83_182 VDD VSS sg13g2_decap_8
XFILLER_17_42 VDD VSS sg13g2_decap_8
XFILLER_16_238 VDD VSS sg13g2_decap_8
XFILLER_56_385 VDD VSS sg13g2_decap_8
XFILLER_44_525 VDD VSS sg13g2_decap_8
XFILLER_12_455 VDD VSS sg13g2_decap_8
XFILLER_40_742 VDD VSS sg13g2_decap_8
XFILLER_33_63 VDD VSS sg13g2_decap_8
XFILLER_8_448 VDD VSS sg13g2_decap_8
XFILLER_4_665 VDD VSS sg13g2_decap_8
XFILLER_3_175 VDD VSS sg13g2_decap_8
XFILLER_79_455 VDD VSS sg13g2_decap_8
XFILLER_39_308 VDD VSS sg13g2_decap_8
XFILLER_67_639 VDD VSS sg13g2_decap_8
XFILLER_66_105 VDD VSS sg13g2_decap_8
XFILLER_82_609 VDD VSS sg13g2_decap_8
XFILLER_94_469 VDD VSS sg13g2_decap_8
XFILLER_12_7 VDD VSS sg13g2_decap_8
XFILLER_75_683 VDD VSS sg13g2_decap_8
XFILLER_81_119 VDD VSS sg13g2_decap_8
XFILLER_74_182 VDD VSS sg13g2_decap_8
XFILLER_62_322 VDD VSS sg13g2_decap_8
XFILLER_74_70 VDD VSS sg13g2_decap_8
XFILLER_47_385 VDD VSS sg13g2_decap_8
XFILLER_35_525 VDD VSS sg13g2_decap_8
XFILLER_90_686 VDD VSS sg13g2_decap_8
XFILLER_62_399 VDD VSS sg13g2_decap_8
XFILLER_50_539 VDD VSS sg13g2_decap_8
XFILLER_31_742 VDD VSS sg13g2_decap_8
XFILLER_90_91 VDD VSS sg13g2_decap_8
XFILLER_30_252 VDD VSS sg13g2_decap_8
XFILLER_57_105 VDD VSS sg13g2_decap_8
XFILLER_85_469 VDD VSS sg13g2_decap_8
XFILLER_72_119 VDD VSS sg13g2_decap_8
XFILLER_26_503 VDD VSS sg13g2_decap_8
XFILLER_65_182 VDD VSS sg13g2_decap_8
XFILLER_38_385 VDD VSS sg13g2_decap_8
XFILLER_53_322 VDD VSS sg13g2_decap_8
XFILLER_81_686 VDD VSS sg13g2_decap_8
XFILLER_53_399 VDD VSS sg13g2_decap_8
XFILLER_41_539 VDD VSS sg13g2_decap_8
XFILLER_80_196 VDD VSS sg13g2_decap_8
XFILLER_22_742 VDD VSS sg13g2_decap_8
XFILLER_70_28 VDD VSS sg13g2_decap_8
XFILLER_21_252 VDD VSS sg13g2_decap_8
XFILLER_1_602 VDD VSS sg13g2_decap_8
XFILLER_89_742 VDD VSS sg13g2_decap_8
XFILLER_0_112 VDD VSS sg13g2_decap_8
XFILLER_88_252 VDD VSS sg13g2_decap_8
XFILLER_95_14 VDD VSS sg13g2_decap_8
XFILLER_1_679 VDD VSS sg13g2_decap_8
XFILLER_48_105 VDD VSS sg13g2_decap_8
XFILLER_64_609 VDD VSS sg13g2_decap_8
XFILLER_76_447 VDD VSS sg13g2_decap_8
XFILLER_0_189 VDD VSS sg13g2_decap_8
XFILLER_91_406 VDD VSS sg13g2_decap_8
XFILLER_63_119 VDD VSS sg13g2_decap_8
XFILLER_57_672 VDD VSS sg13g2_decap_8
XFILLER_28_63 VDD VSS sg13g2_decap_8
XFILLER_29_385 VDD VSS sg13g2_decap_8
XFILLER_44_322 VDD VSS sg13g2_decap_8
XFILLER_56_182 VDD VSS sg13g2_decap_8
XFILLER_17_525 VDD VSS sg13g2_decap_8
XFILLER_72_642 VDD VSS sg13g2_decap_8
XFILLER_44_399 VDD VSS sg13g2_decap_8
XFILLER_32_539 VDD VSS sg13g2_decap_8
XFILLER_71_196 VDD VSS sg13g2_decap_8
XFILLER_13_742 VDD VSS sg13g2_decap_8
XFILLER_44_84 VDD VSS sg13g2_decap_8
XFILLER_9_735 VDD VSS sg13g2_decap_8
XFILLER_12_252 VDD VSS sg13g2_decap_8
XFILLER_8_245 VDD VSS sg13g2_decap_8
XFILLER_4_462 VDD VSS sg13g2_decap_8
XFILLER_5_56 VDD VSS sg13g2_decap_8
XFILLER_69_70 VDD VSS sg13g2_decap_8
XFILLER_79_252 VDD VSS sg13g2_decap_8
XFILLER_39_105 VDD VSS sg13g2_decap_8
XFILLER_95_756 VDD VSS sg13g2_fill_1
XFILLER_67_436 VDD VSS sg13g2_decap_8
XFILLER_94_266 VDD VSS sg13g2_decap_8
XFILLER_82_406 VDD VSS sg13g2_decap_8
XFILLER_55_609 VDD VSS sg13g2_decap_8
XFILLER_48_672 VDD VSS sg13g2_decap_8
XFILLER_63_620 VDD VSS sg13g2_decap_8
XFILLER_75_480 VDD VSS sg13g2_decap_8
XFILLER_85_91 VDD VSS sg13g2_decap_8
XFILLER_35_322 VDD VSS sg13g2_decap_8
XFILLER_47_182 VDD VSS sg13g2_decap_8
XFILLER_54_119 VDD VSS sg13g2_decap_8
XFILLER_90_483 VDD VSS sg13g2_decap_8
XFILLER_63_697 VDD VSS sg13g2_decap_8
XFILLER_35_399 VDD VSS sg13g2_decap_8
XFILLER_23_539 VDD VSS sg13g2_decap_8
XFILLER_62_196 VDD VSS sg13g2_decap_8
XFILLER_50_336 VDD VSS sg13g2_decap_8
XFILLER_86_0 VDD VSS sg13g2_decap_8
XFILLER_86_756 VDD VSS sg13g2_fill_1
XFILLER_85_266 VDD VSS sg13g2_decap_8
XFILLER_65_28 VDD VSS sg13g2_decap_8
XFILLER_46_609 VDD VSS sg13g2_decap_8
XFILLER_58_469 VDD VSS sg13g2_decap_8
XFILLER_39_672 VDD VSS sg13g2_decap_8
XFILLER_73_428 VDD VSS sg13g2_decap_8
XFILLER_26_300 VDD VSS sg13g2_decap_8
XFILLER_38_182 VDD VSS sg13g2_decap_8
XFILLER_45_119 VDD VSS sg13g2_decap_8
XFILLER_81_483 VDD VSS sg13g2_decap_8
XFILLER_54_686 VDD VSS sg13g2_decap_8
XFILLER_26_377 VDD VSS sg13g2_decap_8
XFILLER_14_539 VDD VSS sg13g2_decap_8
XFILLER_81_49 VDD VSS sg13g2_decap_8
XFILLER_41_336 VDD VSS sg13g2_decap_8
XFILLER_53_196 VDD VSS sg13g2_decap_8
XFILLER_14_21 VDD VSS sg13g2_decap_8
XFILLER_10_756 VDD VSS sg13g2_fill_1
XFILLER_14_98 VDD VSS sg13g2_decap_8
XFILLER_6_749 VDD VSS sg13g2_decap_8
XFILLER_5_259 VDD VSS sg13g2_decap_8
XFILLER_30_42 VDD VSS sg13g2_decap_8
XFILLER_77_723 VDD VSS sg13g2_decap_8
XFILLER_1_476 VDD VSS sg13g2_decap_8
XFILLER_39_84 VDD VSS sg13g2_decap_8
XFILLER_64_406 VDD VSS sg13g2_decap_8
XFILLER_49_469 VDD VSS sg13g2_decap_8
XFILLER_37_609 VDD VSS sg13g2_decap_8
XFILLER_91_203 VDD VSS sg13g2_decap_8
XFILLER_76_299 VDD VSS sg13g2_decap_8
XFILLER_17_322 VDD VSS sg13g2_decap_8
XFILLER_36_119 VDD VSS sg13g2_decap_8
XFILLER_29_182 VDD VSS sg13g2_decap_8
XFILLER_60_623 VDD VSS sg13g2_decap_8
XFILLER_45_686 VDD VSS sg13g2_decap_8
XFILLER_17_399 VDD VSS sg13g2_decap_8
XFILLER_32_336 VDD VSS sg13g2_decap_8
XFILLER_44_196 VDD VSS sg13g2_decap_8
XFILLER_9_532 VDD VSS sg13g2_decap_8
XFILLER_68_734 VDD VSS sg13g2_decap_8
XFILLER_67_233 VDD VSS sg13g2_decap_8
XFILLER_95_553 VDD VSS sg13g2_decap_8
XFILLER_55_406 VDD VSS sg13g2_decap_8
XFILLER_28_609 VDD VSS sg13g2_decap_8
XFILLER_82_203 VDD VSS sg13g2_decap_8
XFILLER_27_119 VDD VSS sg13g2_decap_8
XFILLER_51_623 VDD VSS sg13g2_decap_8
XFILLER_36_686 VDD VSS sg13g2_decap_8
XFILLER_63_494 VDD VSS sg13g2_decap_8
XFILLER_90_280 VDD VSS sg13g2_decap_8
XFILLER_23_336 VDD VSS sg13g2_decap_8
XFILLER_35_196 VDD VSS sg13g2_decap_8
XFILLER_50_133 VDD VSS sg13g2_decap_8
XFILLER_76_49 VDD VSS sg13g2_decap_8
XFILLER_59_756 VDD VSS sg13g2_fill_1
XFILLER_86_553 VDD VSS sg13g2_decap_8
XFILLER_46_406 VDD VSS sg13g2_decap_8
XFILLER_58_266 VDD VSS sg13g2_decap_8
XFILLER_19_609 VDD VSS sg13g2_decap_8
XFILLER_73_203 VDD VSS sg13g2_decap_8
XFILLER_18_119 VDD VSS sg13g2_decap_8
XFILLER_27_686 VDD VSS sg13g2_decap_8
XFILLER_81_280 VDD VSS sg13g2_decap_8
XFILLER_54_483 VDD VSS sg13g2_decap_8
Xinputs\[6\].input_pad IOVDD IOVSS _51_/D input_PAD[6] VDD VSS sg13g2_IOPadIn
XFILLER_25_42 VDD VSS sg13g2_decap_8
XFILLER_14_336 VDD VSS sg13g2_decap_8
XFILLER_26_196 VDD VSS sg13g2_decap_8
XFILLER_42_623 VDD VSS sg13g2_decap_8
XFILLER_41_133 VDD VSS sg13g2_decap_8
XFILLER_10_553 VDD VSS sg13g2_decap_8
XFILLER_41_63 VDD VSS sg13g2_decap_8
XFILLER_6_546 VDD VSS sg13g2_decap_8
XFILLER_77_520 VDD VSS sg13g2_decap_8
XFILLER_2_35 VDD VSS sg13g2_decap_8
XFILLER_1_273 VDD VSS sg13g2_decap_8
X_51_ _51_/B _51_/C _51_/A _57_/A VDD VSS _51_/D sg13g2_nand4_1
XFILLER_37_406 VDD VSS sg13g2_decap_8
XFILLER_49_266 VDD VSS sg13g2_decap_8
XFILLER_77_597 VDD VSS sg13g2_decap_8
XFILLER_64_203 VDD VSS sg13g2_decap_8
XFILLER_92_567 VDD VSS sg13g2_decap_8
XFILLER_80_707 VDD VSS sg13g2_decap_8
XFILLER_18_686 VDD VSS sg13g2_decap_8
XFILLER_17_196 VDD VSS sg13g2_decap_8
XFILLER_60_420 VDD VSS sg13g2_decap_8
XFILLER_33_623 VDD VSS sg13g2_decap_8
XFILLER_45_483 VDD VSS sg13g2_decap_8
XFILLER_82_70 VDD VSS sg13g2_decap_8
XFILLER_32_133 VDD VSS sg13g2_decap_8
XFILLER_60_497 VDD VSS sg13g2_decap_8
XFILLER_49_0 VDD VSS sg13g2_decap_8
XFILLER_68_531 VDD VSS sg13g2_decap_8
XFILLER_95_350 VDD VSS sg13g2_decap_8
XFILLER_28_406 VDD VSS sg13g2_decap_8
XFILLER_55_203 VDD VSS sg13g2_decap_8
XFILLER_83_567 VDD VSS sg13g2_decap_8
XFILLER_70_228 VDD VSS sg13g2_decap_8
XFILLER_63_280 VDD VSS sg13g2_decap_8
XFILLER_51_420 VDD VSS sg13g2_decap_8
XFILLER_24_623 VDD VSS sg13g2_decap_8
XFILLER_36_483 VDD VSS sg13g2_decap_8
XFILLER_23_133 VDD VSS sg13g2_decap_8
XFILLER_51_497 VDD VSS sg13g2_decap_8
XFILLER_11_77 VDD VSS sg13g2_decap_8
XFILLER_86_350 VDD VSS sg13g2_decap_8
XFILLER_59_553 VDD VSS sg13g2_decap_8
XFILLER_19_406 VDD VSS sg13g2_decap_8
XFILLER_46_203 VDD VSS sg13g2_decap_8
XFILLER_74_567 VDD VSS sg13g2_decap_8
XFILLER_62_707 VDD VSS sg13g2_decap_8
XFILLER_36_63 VDD VSS sg13g2_decap_8
XFILLER_61_217 VDD VSS sg13g2_decap_8
XFILLER_42_420 VDD VSS sg13g2_decap_8
XFILLER_54_280 VDD VSS sg13g2_decap_8
XFILLER_15_623 VDD VSS sg13g2_decap_8
XFILLER_27_483 VDD VSS sg13g2_decap_8
XFILLER_14_133 VDD VSS sg13g2_decap_8
XFILLER_30_637 VDD VSS sg13g2_decap_8
XFILLER_42_497 VDD VSS sg13g2_decap_8
XFILLER_52_84 VDD VSS sg13g2_decap_8
XFILLER_10_350 VDD VSS sg13g2_decap_8
XFILLER_6_343 VDD VSS sg13g2_decap_8
XFILLER_69_317 VDD VSS sg13g2_decap_8
XFILLER_2_560 VDD VSS sg13g2_decap_8
XFILLER_42_7 VDD VSS sg13g2_decap_8
XFILLER_77_70 VDD VSS sg13g2_decap_8
XFILLER_77_372 VDD VSS sg13g2_decap_8
XFILLER_37_203 VDD VSS sg13g2_decap_8
XFILLER_65_556 VDD VSS sg13g2_decap_8
XFILLER_53_707 VDD VSS sg13g2_decap_8
XFILLER_80_504 VDD VSS sg13g2_decap_8
XFILLER_92_364 VDD VSS sg13g2_decap_8
XFILLER_52_217 VDD VSS sg13g2_decap_8
XFILLER_93_91 VDD VSS sg13g2_decap_8
XFILLER_33_420 VDD VSS sg13g2_decap_8
XFILLER_45_280 VDD VSS sg13g2_decap_8
XFILLER_18_483 VDD VSS sg13g2_decap_8
XFILLER_21_637 VDD VSS sg13g2_decap_8
XFILLER_33_497 VDD VSS sg13g2_decap_8
XFILLER_20_147 VDD VSS sg13g2_decap_8
XFILLER_60_294 VDD VSS sg13g2_decap_8
XFILLER_88_637 VDD VSS sg13g2_decap_8
XIO_BOND_clk_pad clk_PAD bondpad_70x70_novias
XFILLER_87_147 VDD VSS sg13g2_decap_8
XFILLER_28_203 VDD VSS sg13g2_decap_8
XFILLER_83_364 VDD VSS sg13g2_decap_8
XFILLER_73_28 VDD VSS sg13g2_decap_8
XFILLER_56_567 VDD VSS sg13g2_decap_8
XFILLER_44_707 VDD VSS sg13g2_decap_8
XFILLER_71_548 VDD VSS sg13g2_decap_8
XFILLER_24_420 VDD VSS sg13g2_decap_8
XFILLER_36_280 VDD VSS sg13g2_decap_8
XFILLER_43_217 VDD VSS sg13g2_decap_8
XFILLER_12_637 VDD VSS sg13g2_decap_8
XFILLER_24_497 VDD VSS sg13g2_decap_8
XFILLER_11_147 VDD VSS sg13g2_decap_8
XFILLER_51_294 VDD VSS sg13g2_decap_8
XFILLER_22_21 VDD VSS sg13g2_decap_8
XFILLER_22_98 VDD VSS sg13g2_decap_8
XFILLER_3_357 VDD VSS sg13g2_decap_8
XFILLER_79_637 VDD VSS sg13g2_decap_8
XFILLER_78_147 VDD VSS sg13g2_decap_8
XFILLER_19_203 VDD VSS sg13g2_decap_8
XFILLER_59_350 VDD VSS sg13g2_decap_8
XFILLER_62_504 VDD VSS sg13g2_decap_8
XFILLER_47_567 VDD VSS sg13g2_decap_8
XFILLER_47_84 VDD VSS sg13g2_decap_8
XFILLER_35_707 VDD VSS sg13g2_decap_8
XFILLER_15_420 VDD VSS sg13g2_decap_8
XFILLER_27_280 VDD VSS sg13g2_decap_8
XFILLER_34_217 VDD VSS sg13g2_decap_8
XFILLER_30_434 VDD VSS sg13g2_decap_8
XFILLER_42_294 VDD VSS sg13g2_decap_8
XFILLER_15_497 VDD VSS sg13g2_decap_8
XFILLER_8_56 VDD VSS sg13g2_decap_8
XFILLER_7_630 VDD VSS sg13g2_decap_8
XFILLER_6_140 VDD VSS sg13g2_decap_8
XFILLER_88_91 VDD VSS sg13g2_decap_8
XFILLER_69_147 VDD VSS sg13g2_decap_8
XFILLER_93_651 VDD VSS sg13g2_decap_8
XFILLER_80_301 VDD VSS sg13g2_decap_8
XFILLER_65_364 VDD VSS sg13g2_decap_8
XFILLER_53_504 VDD VSS sg13g2_decap_8
XFILLER_38_567 VDD VSS sg13g2_decap_8
XFILLER_92_161 VDD VSS sg13g2_decap_8
XFILLER_25_217 VDD VSS sg13g2_decap_8
XFILLER_18_280 VDD VSS sg13g2_decap_8
XFILLER_80_378 VDD VSS sg13g2_decap_8
XFILLER_61_581 VDD VSS sg13g2_decap_8
XFILLER_21_434 VDD VSS sg13g2_decap_8
XFILLER_33_294 VDD VSS sg13g2_decap_8
XFILLER_88_434 VDD VSS sg13g2_decap_8
XFILLER_68_28 VDD VSS sg13g2_decap_8
XFILLER_76_629 VDD VSS sg13g2_decap_8
XFILLER_69_692 VDD VSS sg13g2_decap_8
XFILLER_84_651 VDD VSS sg13g2_decap_8
XFILLER_84_49 VDD VSS sg13g2_decap_8
XFILLER_17_21 VDD VSS sg13g2_decap_8
XFILLER_56_364 VDD VSS sg13g2_decap_8
XFILLER_17_707 VDD VSS sg13g2_decap_8
XFILLER_29_567 VDD VSS sg13g2_decap_8
XFILLER_44_504 VDD VSS sg13g2_decap_8
XFILLER_83_161 VDD VSS sg13g2_decap_8
XFILLER_16_217 VDD VSS sg13g2_decap_8
XFILLER_71_345 VDD VSS sg13g2_decap_8
XFILLER_17_98 VDD VSS sg13g2_decap_8
XFILLER_52_581 VDD VSS sg13g2_decap_8
XFILLER_40_721 VDD VSS sg13g2_decap_8
XFILLER_12_434 VDD VSS sg13g2_decap_8
XFILLER_33_42 VDD VSS sg13g2_decap_8
XFILLER_24_294 VDD VSS sg13g2_decap_8
XFILLER_8_427 VDD VSS sg13g2_decap_8
XFILLER_4_644 VDD VSS sg13g2_decap_8
XFILLER_3_154 VDD VSS sg13g2_decap_8
XFILLER_79_434 VDD VSS sg13g2_decap_8
XFILLER_67_618 VDD VSS sg13g2_decap_8
XFILLER_94_448 VDD VSS sg13g2_decap_8
XFILLER_75_662 VDD VSS sg13g2_decap_8
XFILLER_47_364 VDD VSS sg13g2_decap_8
XFILLER_35_504 VDD VSS sg13g2_decap_8
XFILLER_74_161 VDD VSS sg13g2_decap_8
XFILLER_62_301 VDD VSS sg13g2_decap_8
XFILLER_90_665 VDD VSS sg13g2_decap_8
XFILLER_62_378 VDD VSS sg13g2_decap_8
XFILLER_50_518 VDD VSS sg13g2_decap_8
XFILLER_31_721 VDD VSS sg13g2_decap_8
XFILLER_15_294 VDD VSS sg13g2_decap_8
XFILLER_30_231 VDD VSS sg13g2_decap_8
XFILLER_43_581 VDD VSS sg13g2_decap_8
XFILLER_90_70 VDD VSS sg13g2_decap_8
XFILLER_31_0 VDD VSS sg13g2_decap_8
XFILLER_85_448 VDD VSS sg13g2_decap_8
XFILLER_38_364 VDD VSS sg13g2_decap_8
XFILLER_66_695 VDD VSS sg13g2_decap_8
XFILLER_65_161 VDD VSS sg13g2_decap_8
XFILLER_53_301 VDD VSS sg13g2_decap_8
XFILLER_81_665 VDD VSS sg13g2_decap_8
XFILLER_26_559 VDD VSS sg13g2_decap_8
XFILLER_80_175 VDD VSS sg13g2_decap_8
XFILLER_53_378 VDD VSS sg13g2_decap_8
XFILLER_41_518 VDD VSS sg13g2_decap_8
XFILLER_22_721 VDD VSS sg13g2_decap_8
XFILLER_34_581 VDD VSS sg13g2_decap_8
XFILLER_21_231 VDD VSS sg13g2_decap_8
XFILLER_79_49 VDD VSS sg13g2_decap_8
XFILLER_89_721 VDD VSS sg13g2_decap_8
XFILLER_88_231 VDD VSS sg13g2_decap_8
XFILLER_1_658 VDD VSS sg13g2_decap_8
XFILLER_76_426 VDD VSS sg13g2_decap_8
XFILLER_0_168 VDD VSS sg13g2_decap_8
XFILLER_57_651 VDD VSS sg13g2_decap_8
XFILLER_28_42 VDD VSS sg13g2_decap_8
XFILLER_29_364 VDD VSS sg13g2_decap_8
XFILLER_17_504 VDD VSS sg13g2_decap_8
XFILLER_72_621 VDD VSS sg13g2_decap_8
XFILLER_44_301 VDD VSS sg13g2_decap_8
XFILLER_56_161 VDD VSS sg13g2_decap_8
XFILLER_72_698 VDD VSS sg13g2_decap_8
XFILLER_71_175 VDD VSS sg13g2_decap_8
XFILLER_44_378 VDD VSS sg13g2_decap_8
XFILLER_32_518 VDD VSS sg13g2_decap_8
XFILLER_13_721 VDD VSS sg13g2_decap_8
XFILLER_44_63 VDD VSS sg13g2_decap_8
XFILLER_25_581 VDD VSS sg13g2_decap_8
XFILLER_9_714 VDD VSS sg13g2_decap_8
XFILLER_12_231 VDD VSS sg13g2_decap_8
XFILLER_8_224 VDD VSS sg13g2_decap_8
XFILLER_40_595 VDD VSS sg13g2_decap_8
XFILLER_60_84 VDD VSS sg13g2_decap_8
XFILLER_4_441 VDD VSS sg13g2_decap_8
XFILLER_5_35 VDD VSS sg13g2_decap_8
XFILLER_79_231 VDD VSS sg13g2_decap_8
XFILLER_67_415 VDD VSS sg13g2_decap_8
XFILLER_95_735 VDD VSS sg13g2_decap_8
XFILLER_94_245 VDD VSS sg13g2_decap_8
XFILLER_85_70 VDD VSS sg13g2_decap_8
XFILLER_48_651 VDD VSS sg13g2_decap_8
XFILLER_35_301 VDD VSS sg13g2_decap_8
XFILLER_47_161 VDD VSS sg13g2_decap_8
XFILLER_63_676 VDD VSS sg13g2_decap_8
XFILLER_90_462 VDD VSS sg13g2_decap_8
XFILLER_62_175 VDD VSS sg13g2_decap_8
XFILLER_35_378 VDD VSS sg13g2_decap_8
XFILLER_50_315 VDD VSS sg13g2_decap_8
XFILLER_23_518 VDD VSS sg13g2_decap_8
XFILLER_16_581 VDD VSS sg13g2_decap_8
XFILLER_31_595 VDD VSS sg13g2_decap_8
XFILLER_79_0 VDD VSS sg13g2_decap_8
XFILLER_86_735 VDD VSS sg13g2_decap_8
XFILLER_58_448 VDD VSS sg13g2_decap_8
XFILLER_85_245 VDD VSS sg13g2_decap_8
XFILLER_39_651 VDD VSS sg13g2_decap_8
XFILLER_38_161 VDD VSS sg13g2_decap_8
XFILLER_66_492 VDD VSS sg13g2_decap_8
XFILLER_54_665 VDD VSS sg13g2_decap_8
Xinputs\[5\].input_pad IOVDD IOVSS _51_/C input_PAD[5] VDD VSS sg13g2_IOPadIn
XFILLER_26_356 VDD VSS sg13g2_decap_8
XFILLER_81_462 VDD VSS sg13g2_decap_8
XFILLER_41_315 VDD VSS sg13g2_decap_8
XFILLER_53_175 VDD VSS sg13g2_decap_8
XFILLER_14_518 VDD VSS sg13g2_decap_8
XFILLER_81_28 VDD VSS sg13g2_decap_8
XFILLER_10_735 VDD VSS sg13g2_decap_8
XFILLER_14_77 VDD VSS sg13g2_decap_8
XFILLER_22_595 VDD VSS sg13g2_decap_8
XFILLER_6_728 VDD VSS sg13g2_decap_8
XFILLER_30_21 VDD VSS sg13g2_decap_8
XFILLER_5_238 VDD VSS sg13g2_decap_8
XFILLER_30_98 VDD VSS sg13g2_decap_8
XFILLER_77_702 VDD VSS sg13g2_decap_8
Xclk_pad IOVDD IOVSS clk_pad/p2c clk_PAD VDD VSS sg13g2_IOPadIn
XFILLER_1_455 VDD VSS sg13g2_decap_8
XFILLER_89_595 VDD VSS sg13g2_decap_8
XFILLER_39_63 VDD VSS sg13g2_decap_8
XFILLER_49_448 VDD VSS sg13g2_decap_8
XFILLER_92_749 VDD VSS sg13g2_decap_8
XFILLER_76_278 VDD VSS sg13g2_decap_8
XFILLER_17_301 VDD VSS sg13g2_decap_8
XFILLER_29_161 VDD VSS sg13g2_decap_8
XFILLER_91_259 VDD VSS sg13g2_decap_8
XFILLER_60_602 VDD VSS sg13g2_decap_8
XFILLER_55_84 VDD VSS sg13g2_decap_8
XFILLER_17_378 VDD VSS sg13g2_decap_8
XFILLER_45_665 VDD VSS sg13g2_decap_8
XFILLER_72_495 VDD VSS sg13g2_decap_8
XFILLER_32_315 VDD VSS sg13g2_decap_8
XFILLER_44_175 VDD VSS sg13g2_decap_8
XFILLER_60_679 VDD VSS sg13g2_decap_8
XFILLER_13_595 VDD VSS sg13g2_decap_8
XFILLER_9_511 VDD VSS sg13g2_decap_8
XFILLER_72_7 VDD VSS sg13g2_decap_8
XFILLER_40_392 VDD VSS sg13g2_decap_8
XFILLER_9_588 VDD VSS sg13g2_decap_8
XFILLER_68_713 VDD VSS sg13g2_decap_8
XFILLER_95_532 VDD VSS sg13g2_decap_8
XFILLER_67_212 VDD VSS sg13g2_decap_8
XFILLER_83_749 VDD VSS sg13g2_decap_8
XFILLER_67_289 VDD VSS sg13g2_decap_8
XFILLER_82_259 VDD VSS sg13g2_decap_8
XFILLER_51_602 VDD VSS sg13g2_decap_8
XFILLER_36_665 VDD VSS sg13g2_decap_8
XFILLER_23_315 VDD VSS sg13g2_decap_8
XFILLER_35_175 VDD VSS sg13g2_decap_8
XFILLER_50_112 VDD VSS sg13g2_decap_8
XFILLER_51_679 VDD VSS sg13g2_decap_8
XFILLER_50_189 VDD VSS sg13g2_decap_8
XFILLER_31_392 VDD VSS sg13g2_decap_8
XFILLER_86_532 VDD VSS sg13g2_decap_8
XFILLER_76_28 VDD VSS sg13g2_decap_8
XFILLER_59_735 VDD VSS sg13g2_decap_8
XFILLER_58_245 VDD VSS sg13g2_decap_8
XFILLER_74_749 VDD VSS sg13g2_decap_8
XFILLER_92_49 VDD VSS sg13g2_decap_8
XFILLER_25_21 VDD VSS sg13g2_decap_8
XFILLER_54_462 VDD VSS sg13g2_decap_8
XFILLER_27_665 VDD VSS sg13g2_decap_8
XFILLER_42_602 VDD VSS sg13g2_decap_8
XFILLER_14_315 VDD VSS sg13g2_decap_8
XFILLER_26_175 VDD VSS sg13g2_decap_8
XFILLER_41_112 VDD VSS sg13g2_decap_8
XFILLER_42_679 VDD VSS sg13g2_decap_8
XFILLER_25_98 VDD VSS sg13g2_decap_8
XFILLER_41_189 VDD VSS sg13g2_decap_8
XFILLER_10_532 VDD VSS sg13g2_decap_8
XFILLER_22_392 VDD VSS sg13g2_decap_8
XFILLER_6_525 VDD VSS sg13g2_decap_8
XFILLER_41_42 VDD VSS sg13g2_decap_8
XFILLER_2_742 VDD VSS sg13g2_decap_8
XFILLER_9_0 VDD VSS sg13g2_decap_8
XFILLER_1_252 VDD VSS sg13g2_decap_8
XFILLER_89_392 VDD VSS sg13g2_decap_8
XFILLER_2_14 VDD VSS sg13g2_decap_8
X_50_ _60_/B _60_/C _50_/Y VDD VSS sg13g2_nor2_1
XFILLER_49_245 VDD VSS sg13g2_decap_8
XFILLER_77_576 VDD VSS sg13g2_decap_8
XFILLER_65_738 VDD VSS sg13g2_decap_8
XFILLER_92_546 VDD VSS sg13g2_decap_8
XFILLER_64_259 VDD VSS sg13g2_decap_8
XFILLER_45_462 VDD VSS sg13g2_decap_8
XFILLER_18_665 VDD VSS sg13g2_decap_8
XFILLER_33_602 VDD VSS sg13g2_decap_8
XFILLER_72_270 VDD VSS sg13g2_decap_8
XFILLER_17_175 VDD VSS sg13g2_decap_8
XFILLER_32_112 VDD VSS sg13g2_decap_8
XFILLER_33_679 VDD VSS sg13g2_decap_8
XFILLER_20_329 VDD VSS sg13g2_decap_8
XFILLER_32_189 VDD VSS sg13g2_decap_8
XFILLER_60_476 VDD VSS sg13g2_decap_8
XFILLER_13_392 VDD VSS sg13g2_decap_8
XFILLER_9_385 VDD VSS sg13g2_decap_8
XFILLER_68_510 VDD VSS sg13g2_decap_8
XFILLER_87_329 VDD VSS sg13g2_decap_8
XFILLER_68_587 VDD VSS sg13g2_decap_8
XFILLER_56_749 VDD VSS sg13g2_decap_8
XFILLER_83_546 VDD VSS sg13g2_decap_8
XFILLER_36_462 VDD VSS sg13g2_decap_8
XFILLER_55_259 VDD VSS sg13g2_decap_8
XFILLER_24_602 VDD VSS sg13g2_decap_8
XFILLER_23_112 VDD VSS sg13g2_decap_8
XFILLER_24_679 VDD VSS sg13g2_decap_8
XFILLER_11_329 VDD VSS sg13g2_decap_8
XFILLER_23_189 VDD VSS sg13g2_decap_8
XFILLER_51_476 VDD VSS sg13g2_decap_8
XFILLER_11_56 VDD VSS sg13g2_decap_8
XFILLER_3_539 VDD VSS sg13g2_decap_8
XFILLER_87_49 VDD VSS sg13g2_decap_8
XFILLER_2_7 VDD VSS sg13g2_decap_8
XFILLER_78_329 VDD VSS sg13g2_decap_8
XFILLER_59_532 VDD VSS sg13g2_decap_8
XFILLER_74_546 VDD VSS sg13g2_decap_8
XFILLER_47_749 VDD VSS sg13g2_decap_8
XFILLER_36_42 VDD VSS sg13g2_decap_8
XFILLER_27_462 VDD VSS sg13g2_decap_8
XFILLER_46_259 VDD VSS sg13g2_decap_8
XFILLER_15_602 VDD VSS sg13g2_decap_8
XFILLER_14_112 VDD VSS sg13g2_decap_8
XFILLER_15_679 VDD VSS sg13g2_decap_8
XFILLER_14_189 VDD VSS sg13g2_decap_8
XFILLER_42_476 VDD VSS sg13g2_decap_8
XFILLER_30_616 VDD VSS sg13g2_decap_8
XFILLER_52_63 VDD VSS sg13g2_decap_8
XFILLER_6_322 VDD VSS sg13g2_decap_8
XFILLER_6_399 VDD VSS sg13g2_decap_8
XFILLER_35_7 VDD VSS sg13g2_decap_8
XFILLER_77_351 VDD VSS sg13g2_decap_8
XFILLER_65_535 VDD VSS sg13g2_decap_8
XFILLER_92_343 VDD VSS sg13g2_decap_8
XFILLER_38_749 VDD VSS sg13g2_decap_8
XFILLER_18_462 VDD VSS sg13g2_decap_8
XFILLER_37_259 VDD VSS sg13g2_decap_8
XFILLER_73_590 VDD VSS sg13g2_decap_8
XFILLER_93_70 VDD VSS sg13g2_decap_8
XFILLER_33_476 VDD VSS sg13g2_decap_8
XFILLER_60_273 VDD VSS sg13g2_decap_8
XFILLER_21_616 VDD VSS sg13g2_decap_8
XFILLER_20_126 VDD VSS sg13g2_decap_8
XFILLER_9_182 VDD VSS sg13g2_decap_8
XFILLER_61_0 VDD VSS sg13g2_decap_8
XFILLER_88_616 VDD VSS sg13g2_decap_8
XFILLER_87_126 VDD VSS sg13g2_decap_8
XFILLER_68_384 VDD VSS sg13g2_decap_8
XFILLER_56_546 VDD VSS sg13g2_decap_8
XFILLER_29_749 VDD VSS sg13g2_decap_8
XFILLER_83_343 VDD VSS sg13g2_decap_8
XFILLER_28_259 VDD VSS sg13g2_decap_8
XFILLER_71_527 VDD VSS sg13g2_decap_8
XFILLER_12_616 VDD VSS sg13g2_decap_8
XFILLER_24_476 VDD VSS sg13g2_decap_8
XFILLER_51_273 VDD VSS sg13g2_decap_8
XFILLER_8_609 VDD VSS sg13g2_decap_8
XFILLER_11_126 VDD VSS sg13g2_decap_8
XFILLER_7_119 VDD VSS sg13g2_decap_8
XIO_BOND_vss_pads\[0\].vss_pad VSS bondpad_70x70_novias
XFILLER_20_693 VDD VSS sg13g2_decap_8
XFILLER_22_77 VDD VSS sg13g2_decap_8
XFILLER_3_336 VDD VSS sg13g2_decap_8
XFILLER_79_616 VDD VSS sg13g2_decap_8
XFILLER_78_126 VDD VSS sg13g2_decap_8
XFILLER_87_693 VDD VSS sg13g2_decap_8
XFILLER_47_546 VDD VSS sg13g2_decap_8
XFILLER_47_63 VDD VSS sg13g2_decap_8
XFILLER_19_259 VDD VSS sg13g2_decap_8
XFILLER_70_582 VDD VSS sg13g2_decap_8
XFILLER_63_84 VDD VSS sg13g2_decap_8
XFILLER_15_476 VDD VSS sg13g2_decap_8
XFILLER_30_413 VDD VSS sg13g2_decap_8
XFILLER_42_273 VDD VSS sg13g2_decap_8
XFILLER_8_35 VDD VSS sg13g2_decap_8
XFILLER_11_693 VDD VSS sg13g2_decap_8
XFILLER_7_686 VDD VSS sg13g2_decap_8
XFILLER_6_196 VDD VSS sg13g2_decap_8
XFILLER_69_126 VDD VSS sg13g2_decap_8
XFILLER_88_70 VDD VSS sg13g2_decap_8
XFILLER_93_630 VDD VSS sg13g2_decap_8
XFILLER_78_693 VDD VSS sg13g2_decap_8
XFILLER_38_546 VDD VSS sg13g2_decap_8
XFILLER_92_140 VDD VSS sg13g2_decap_8
XFILLER_65_343 VDD VSS sg13g2_decap_8
XFILLER_80_357 VDD VSS sg13g2_decap_8
XFILLER_61_560 VDD VSS sg13g2_decap_8
XFILLER_21_413 VDD VSS sg13g2_decap_8
XFILLER_33_273 VDD VSS sg13g2_decap_8
XFILLER_88_413 VDD VSS sg13g2_decap_8
XFILLER_76_608 VDD VSS sg13g2_decap_8
XFILLER_69_671 VDD VSS sg13g2_decap_8
XFILLER_84_630 VDD VSS sg13g2_decap_8
XFILLER_84_28 VDD VSS sg13g2_decap_8
XFILLER_29_546 VDD VSS sg13g2_decap_8
XFILLER_83_140 VDD VSS sg13g2_decap_8
XFILLER_56_343 VDD VSS sg13g2_decap_8
XFILLER_71_324 VDD VSS sg13g2_decap_8
XFILLER_17_77 VDD VSS sg13g2_decap_8
XFILLER_52_560 VDD VSS sg13g2_decap_8
XFILLER_40_700 VDD VSS sg13g2_decap_8
XFILLER_12_413 VDD VSS sg13g2_decap_8
XFILLER_33_21 VDD VSS sg13g2_decap_8
XFILLER_24_273 VDD VSS sg13g2_decap_8
XFILLER_8_406 VDD VSS sg13g2_decap_8
XFILLER_33_98 VDD VSS sg13g2_decap_8
XFILLER_20_490 VDD VSS sg13g2_decap_8
XFILLER_4_623 VDD VSS sg13g2_decap_8
XFILLER_3_133 VDD VSS sg13g2_decap_8
XFILLER_79_413 VDD VSS sg13g2_decap_8
XFILLER_94_427 VDD VSS sg13g2_decap_8
XFILLER_87_490 VDD VSS sg13g2_decap_8
XFILLER_58_84 VDD VSS sg13g2_decap_8
XFILLER_75_641 VDD VSS sg13g2_decap_8
XFILLER_74_140 VDD VSS sg13g2_decap_8
XFILLER_47_343 VDD VSS sg13g2_decap_8
XFILLER_90_644 VDD VSS sg13g2_decap_8
XFILLER_62_357 VDD VSS sg13g2_decap_8
XFILLER_31_700 VDD VSS sg13g2_decap_8
XFILLER_43_560 VDD VSS sg13g2_decap_8
XFILLER_70_390 VDD VSS sg13g2_decap_8
XFILLER_15_273 VDD VSS sg13g2_decap_8
XFILLER_30_210 VDD VSS sg13g2_decap_8
XFILLER_30_287 VDD VSS sg13g2_decap_8
XFILLER_11_490 VDD VSS sg13g2_decap_8
XFILLER_7_483 VDD VSS sg13g2_decap_8
XFILLER_24_0 VDD VSS sg13g2_decap_8
XFILLER_78_490 VDD VSS sg13g2_decap_8
XFILLER_85_427 VDD VSS sg13g2_decap_8
XFILLER_65_140 VDD VSS sg13g2_decap_8
XFILLER_38_343 VDD VSS sg13g2_decap_8
XFILLER_66_674 VDD VSS sg13g2_decap_8
Xinputs\[4\].input_pad IOVDD IOVSS _52_/C input_PAD[4] VDD VSS sg13g2_IOPadIn
XFILLER_26_538 VDD VSS sg13g2_decap_8
XFILLER_81_644 VDD VSS sg13g2_decap_8
XFILLER_53_357 VDD VSS sg13g2_decap_8
XFILLER_80_154 VDD VSS sg13g2_decap_8
XFILLER_0_91 VDD VSS sg13g2_decap_8
XFILLER_22_700 VDD VSS sg13g2_decap_8
XFILLER_34_560 VDD VSS sg13g2_decap_8
XFILLER_21_210 VDD VSS sg13g2_decap_8
XFILLER_21_287 VDD VSS sg13g2_decap_8
XFILLER_79_28 VDD VSS sg13g2_decap_8
XFILLER_89_700 VDD VSS sg13g2_decap_8
XFILLER_88_210 VDD VSS sg13g2_decap_8
XFILLER_1_637 VDD VSS sg13g2_decap_8
XFILLER_0_147 VDD VSS sg13g2_decap_8
XFILLER_88_287 VDD VSS sg13g2_decap_8
XFILLER_95_49 VDD VSS sg13g2_decap_8
XFILLER_57_630 VDD VSS sg13g2_decap_8
XFILLER_28_21 VDD VSS sg13g2_decap_8
XFILLER_29_343 VDD VSS sg13g2_decap_8
XFILLER_56_140 VDD VSS sg13g2_decap_8
XFILLER_72_600 VDD VSS sg13g2_decap_8
XFILLER_28_98 VDD VSS sg13g2_decap_8
XFILLER_44_357 VDD VSS sg13g2_decap_8
XFILLER_72_677 VDD VSS sg13g2_decap_8
XFILLER_71_154 VDD VSS sg13g2_decap_8
XFILLER_13_700 VDD VSS sg13g2_decap_8
XFILLER_44_42 VDD VSS sg13g2_decap_8
XFILLER_25_560 VDD VSS sg13g2_decap_8
XFILLER_12_210 VDD VSS sg13g2_decap_8
XFILLER_8_203 VDD VSS sg13g2_decap_8
XFILLER_12_287 VDD VSS sg13g2_decap_8
XFILLER_40_574 VDD VSS sg13g2_decap_8
XFILLER_60_63 VDD VSS sg13g2_decap_8
XFILLER_4_420 VDD VSS sg13g2_decap_8
XFILLER_5_14 VDD VSS sg13g2_decap_8
XFILLER_79_210 VDD VSS sg13g2_decap_8
XFILLER_4_497 VDD VSS sg13g2_decap_8
XFILLER_95_714 VDD VSS sg13g2_decap_8
XFILLER_94_224 VDD VSS sg13g2_decap_8
XFILLER_79_287 VDD VSS sg13g2_decap_8
XFILLER_48_630 VDD VSS sg13g2_decap_8
XFILLER_47_140 VDD VSS sg13g2_decap_8
XFILLER_63_655 VDD VSS sg13g2_decap_8
XFILLER_90_441 VDD VSS sg13g2_decap_8
XFILLER_62_154 VDD VSS sg13g2_decap_8
XFILLER_35_357 VDD VSS sg13g2_decap_8
XFILLER_16_560 VDD VSS sg13g2_decap_8
XFILLER_31_574 VDD VSS sg13g2_decap_8
XFILLER_7_280 VDD VSS sg13g2_decap_8
XFILLER_86_714 VDD VSS sg13g2_decap_8
XFILLER_85_224 VDD VSS sg13g2_decap_8
XFILLER_58_427 VDD VSS sg13g2_decap_8
XFILLER_39_630 VDD VSS sg13g2_decap_8
XFILLER_66_471 VDD VSS sg13g2_decap_8
XFILLER_38_140 VDD VSS sg13g2_decap_8
XFILLER_81_441 VDD VSS sg13g2_decap_8
XFILLER_54_644 VDD VSS sg13g2_decap_8
XFILLER_26_335 VDD VSS sg13g2_decap_8
XFILLER_53_154 VDD VSS sg13g2_decap_8
XFILLER_10_714 VDD VSS sg13g2_decap_8
XFILLER_14_56 VDD VSS sg13g2_decap_8
XFILLER_22_574 VDD VSS sg13g2_decap_8
XFILLER_6_707 VDD VSS sg13g2_decap_8
XFILLER_5_217 VDD VSS sg13g2_decap_8
XFILLER_30_77 VDD VSS sg13g2_decap_8
XFILLER_1_434 VDD VSS sg13g2_decap_8
XFILLER_89_574 VDD VSS sg13g2_decap_8
XFILLER_39_42 VDD VSS sg13g2_decap_8
XFILLER_76_224 VDD VSS sg13g2_decap_4
XFILLER_49_427 VDD VSS sg13g2_decap_8
XFILLER_76_257 VDD VSS sg13g2_decap_8
XFILLER_92_728 VDD VSS sg13g2_decap_8
XFILLER_29_140 VDD VSS sg13g2_decap_8
XFILLER_91_238 VDD VSS sg13g2_decap_8
XFILLER_72_430 VDD VSS sg13g2_decap_4
XFILLER_45_644 VDD VSS sg13g2_decap_8
XFILLER_72_474 VDD VSS sg13g2_decap_8
XFILLER_55_63 VDD VSS sg13g2_decap_8
XFILLER_17_357 VDD VSS sg13g2_decap_8
XFILLER_44_154 VDD VSS sg13g2_decap_8
XFILLER_60_658 VDD VSS sg13g2_decap_8
XFILLER_13_574 VDD VSS sg13g2_decap_8
XFILLER_40_371 VDD VSS sg13g2_decap_8
XFILLER_71_84 VDD VSS sg13g2_decap_8
XFILLER_9_567 VDD VSS sg13g2_decap_8
XFILLER_65_7 VDD VSS sg13g2_decap_8
XFILLER_4_294 VDD VSS sg13g2_decap_8
XFILLER_95_511 VDD VSS sg13g2_decap_8
XFILLER_67_202 VDD VSS sg13g2_decap_4
XFILLER_95_588 VDD VSS sg13g2_decap_8
XFILLER_83_728 VDD VSS sg13g2_decap_8
XFILLER_67_268 VDD VSS sg13g2_decap_8
XFILLER_82_238 VDD VSS sg13g2_decap_8
XFILLER_36_644 VDD VSS sg13g2_decap_8
XFILLER_63_441 VDD VSS sg13g2_decap_8
XFILLER_63_452 VDD VSS sg13g2_fill_1
XFILLER_35_154 VDD VSS sg13g2_decap_8
XFILLER_91_0 VDD VSS sg13g2_decap_8
XFILLER_51_658 VDD VSS sg13g2_decap_8
XFILLER_31_371 VDD VSS sg13g2_decap_8
XFILLER_50_168 VDD VSS sg13g2_decap_8
XFILLER_59_714 VDD VSS sg13g2_decap_8
XFILLER_86_511 VDD VSS sg13g2_decap_8
XFILLER_58_224 VDD VSS sg13g2_decap_8
XFILLER_86_588 VDD VSS sg13g2_decap_8
XFILLER_74_728 VDD VSS sg13g2_decap_8
XFILLER_73_238 VDD VSS sg13g2_decap_8
XFILLER_27_644 VDD VSS sg13g2_decap_8
XFILLER_92_28 VDD VSS sg13g2_decap_8
XFILLER_26_154 VDD VSS sg13g2_decap_8
XFILLER_54_441 VDD VSS sg13g2_decap_8
XFILLER_25_77 VDD VSS sg13g2_decap_8
XFILLER_42_658 VDD VSS sg13g2_decap_8
XFILLER_10_511 VDD VSS sg13g2_decap_8
XFILLER_22_371 VDD VSS sg13g2_decap_8
XFILLER_41_168 VDD VSS sg13g2_decap_8
XFILLER_41_21 VDD VSS sg13g2_decap_8
XFILLER_6_504 VDD VSS sg13g2_decap_8
XFILLER_10_588 VDD VSS sg13g2_decap_8
XFILLER_41_98 VDD VSS sg13g2_decap_8
XFILLER_2_721 VDD VSS sg13g2_decap_8
XFILLER_1_231 VDD VSS sg13g2_decap_8
XFILLER_89_371 VDD VSS sg13g2_decap_8
XFILLER_49_224 VDD VSS sg13g2_decap_8
XFILLER_77_555 VDD VSS sg13g2_decap_8
XFILLER_92_525 VDD VSS sg13g2_decap_8
XFILLER_65_717 VDD VSS sg13g2_decap_8
XFILLER_64_238 VDD VSS sg13g2_decap_8
XFILLER_66_84 VDD VSS sg13g2_decap_8
XFILLER_18_644 VDD VSS sg13g2_decap_8
XFILLER_17_154 VDD VSS sg13g2_decap_8
XFILLER_45_441 VDD VSS sg13g2_decap_8
XFILLER_60_455 VDD VSS sg13g2_decap_8
XFILLER_33_658 VDD VSS sg13g2_decap_8
XFILLER_20_308 VDD VSS sg13g2_decap_8
XFILLER_32_168 VDD VSS sg13g2_decap_8
XFILLER_13_371 VDD VSS sg13g2_decap_8
XFILLER_9_364 VDD VSS sg13g2_decap_8
XFILLER_5_581 VDD VSS sg13g2_decap_8
XFILLER_87_308 VDD VSS sg13g2_decap_8
XFILLER_68_566 VDD VSS sg13g2_decap_8
XFILLER_83_525 VDD VSS sg13g2_decap_8
XFILLER_95_385 VDD VSS sg13g2_decap_8
XFILLER_56_728 VDD VSS sg13g2_decap_8
XFILLER_55_238 VDD VSS sg13g2_decap_8
XFILLER_71_709 VDD VSS sg13g2_decap_8
XFILLER_36_441 VDD VSS sg13g2_decap_8
XFILLER_51_455 VDD VSS sg13g2_decap_8
XFILLER_24_658 VDD VSS sg13g2_decap_8
XFILLER_11_308 VDD VSS sg13g2_decap_8
XFILLER_23_168 VDD VSS sg13g2_decap_8
XFILLER_3_518 VDD VSS sg13g2_decap_8
XFILLER_11_35 VDD VSS sg13g2_decap_8
XFILLER_78_308 VDD VSS sg13g2_decap_8
XFILLER_87_28 VDD VSS sg13g2_decap_8
XFILLER_59_511 VDD VSS sg13g2_decap_8
XFILLER_59_588 VDD VSS sg13g2_decap_8
XFILLER_47_728 VDD VSS sg13g2_decap_8
XFILLER_74_525 VDD VSS sg13g2_decap_8
XFILLER_86_385 VDD VSS sg13g2_decap_8
XFILLER_36_21 VDD VSS sg13g2_decap_8
XFILLER_46_238 VDD VSS sg13g2_decap_8
XFILLER_27_441 VDD VSS sg13g2_decap_8
XFILLER_36_98 VDD VSS sg13g2_decap_8
XFILLER_42_455 VDD VSS sg13g2_decap_8
XFILLER_15_658 VDD VSS sg13g2_decap_8
XFILLER_52_42 VDD VSS sg13g2_decap_8
XFILLER_14_168 VDD VSS sg13g2_decap_8
XFILLER_6_301 VDD VSS sg13g2_decap_8
XFILLER_10_385 VDD VSS sg13g2_decap_8
XFILLER_6_378 VDD VSS sg13g2_decap_8
XFILLER_77_330 VDD VSS sg13g2_decap_8
XFILLER_2_595 VDD VSS sg13g2_decap_8
XFILLER_28_7 VDD VSS sg13g2_decap_8
XFILLER_65_514 VDD VSS sg13g2_decap_8
XFILLER_38_728 VDD VSS sg13g2_decap_8
XFILLER_92_322 VDD VSS sg13g2_decap_8
XFILLER_37_238 VDD VSS sg13g2_decap_8
XFILLER_18_441 VDD VSS sg13g2_decap_8
XFILLER_80_539 VDD VSS sg13g2_decap_8
XFILLER_92_399 VDD VSS sg13g2_decap_8
XFILLER_61_742 VDD VSS sg13g2_decap_8
XFILLER_33_455 VDD VSS sg13g2_decap_8
XFILLER_20_105 VDD VSS sg13g2_decap_8
XFILLER_60_252 VDD VSS sg13g2_decap_8
XFILLER_9_161 VDD VSS sg13g2_decap_8
Xoutputs\[0\].output_pad _76_/Q IOVDD IOVSS output_PAD[0] VDD VSS sg13g2_IOPadOut30mA
XFILLER_54_0 VDD VSS sg13g2_decap_8
XFILLER_87_105 VDD VSS sg13g2_decap_8
XFILLER_68_363 VDD VSS sg13g2_decap_8
XFILLER_3_91 VDD VSS sg13g2_decap_8
XFILLER_29_728 VDD VSS sg13g2_decap_8
XFILLER_95_182 VDD VSS sg13g2_decap_8
XFILLER_83_322 VDD VSS sg13g2_decap_8
XFILLER_56_525 VDD VSS sg13g2_decap_8
XFILLER_28_238 VDD VSS sg13g2_decap_8
XFILLER_71_506 VDD VSS sg13g2_decap_8
XFILLER_83_399 VDD VSS sg13g2_decap_8
XFILLER_52_742 VDD VSS sg13g2_decap_8
XFILLER_11_105 VDD VSS sg13g2_decap_8
XFILLER_24_455 VDD VSS sg13g2_decap_8
XFILLER_51_252 VDD VSS sg13g2_decap_8
XFILLER_22_56 VDD VSS sg13g2_decap_8
XFILLER_20_672 VDD VSS sg13g2_decap_8
XFILLER_3_315 VDD VSS sg13g2_decap_8
XFILLER_78_105 VDD VSS sg13g2_decap_8
XFILLER_94_609 VDD VSS sg13g2_decap_8
XFILLER_87_672 VDD VSS sg13g2_decap_8
XFILLER_93_119 VDD VSS sg13g2_decap_8
XFILLER_86_182 VDD VSS sg13g2_decap_8
XFILLER_47_525 VDD VSS sg13g2_decap_8
XFILLER_47_42 VDD VSS sg13g2_decap_8
XFILLER_19_238 VDD VSS sg13g2_decap_8
XFILLER_59_385 VDD VSS sg13g2_decap_8
XFILLER_74_344 VDD VSS sg13g2_decap_8
XFILLER_62_539 VDD VSS sg13g2_decap_8
XFILLER_43_742 VDD VSS sg13g2_decap_8
XFILLER_70_561 VDD VSS sg13g2_decap_8
XFILLER_63_63 VDD VSS sg13g2_decap_8
XFILLER_15_455 VDD VSS sg13g2_decap_8
XFILLER_42_252 VDD VSS sg13g2_decap_8
XFILLER_8_14 VDD VSS sg13g2_decap_8
XFILLER_30_469 VDD VSS sg13g2_decap_8
XFILLER_11_672 VDD VSS sg13g2_decap_8
XFILLER_7_665 VDD VSS sg13g2_decap_8
XFILLER_10_182 VDD VSS sg13g2_decap_8
XFILLER_6_175 VDD VSS sg13g2_decap_8
XFILLER_69_105 VDD VSS sg13g2_decap_8
XFILLER_85_609 VDD VSS sg13g2_decap_8
XFILLER_2_392 VDD VSS sg13g2_decap_8
XFILLER_78_672 VDD VSS sg13g2_decap_8
XFILLER_84_119 VDD VSS sg13g2_decap_8
XFILLER_77_182 VDD VSS sg13g2_decap_8
XFILLER_65_322 VDD VSS sg13g2_decap_8
XFILLER_38_525 VDD VSS sg13g2_decap_8
Xinputs\[3\].input_pad IOVDD IOVSS _51_/B input_PAD[3] VDD VSS sg13g2_IOPadIn
XFILLER_93_686 VDD VSS sg13g2_decap_8
XFILLER_65_399 VDD VSS sg13g2_decap_8
XFILLER_53_539 VDD VSS sg13g2_decap_8
XFILLER_92_196 VDD VSS sg13g2_decap_8
XFILLER_80_336 VDD VSS sg13g2_decap_8
XFILLER_34_742 VDD VSS sg13g2_decap_8
XFILLER_33_252 VDD VSS sg13g2_decap_8
XFILLER_21_469 VDD VSS sg13g2_decap_8
XFILLER_0_329 VDD VSS sg13g2_decap_8
XFILLER_69_650 VDD VSS sg13g2_decap_8
XFILLER_88_469 VDD VSS sg13g2_decap_8
XFILLER_68_182 VDD VSS sg13g2_decap_8
XFILLER_56_322 VDD VSS sg13g2_decap_8
XFILLER_29_525 VDD VSS sg13g2_decap_8
XFILLER_84_686 VDD VSS sg13g2_decap_8
XFILLER_17_56 VDD VSS sg13g2_decap_8
XFILLER_56_399 VDD VSS sg13g2_decap_8
XFILLER_44_539 VDD VSS sg13g2_decap_8
XFILLER_83_196 VDD VSS sg13g2_decap_8
XFILLER_25_742 VDD VSS sg13g2_decap_8
XFILLER_24_252 VDD VSS sg13g2_decap_8
XFILLER_12_469 VDD VSS sg13g2_decap_8
XFILLER_33_77 VDD VSS sg13g2_decap_8
XFILLER_40_756 VDD VSS sg13g2_fill_1
XFILLER_4_602 VDD VSS sg13g2_decap_8
XFILLER_3_112 VDD VSS sg13g2_decap_8
XFILLER_4_679 VDD VSS sg13g2_decap_8
XFILLER_3_189 VDD VSS sg13g2_decap_8
XFILLER_94_406 VDD VSS sg13g2_decap_8
XFILLER_79_469 VDD VSS sg13g2_decap_8
XFILLER_58_63 VDD VSS sg13g2_decap_8
XFILLER_75_620 VDD VSS sg13g2_decap_8
XFILLER_66_119 VDD VSS sg13g2_decap_8
XFILLER_47_322 VDD VSS sg13g2_decap_8
XFILLER_59_182 VDD VSS sg13g2_decap_8
XFILLER_90_623 VDD VSS sg13g2_decap_8
XFILLER_75_697 VDD VSS sg13g2_decap_8
XFILLER_35_539 VDD VSS sg13g2_decap_8
XFILLER_74_196 VDD VSS sg13g2_decap_8
XFILLER_62_336 VDD VSS sg13g2_decap_8
XFILLER_74_84 VDD VSS sg13g2_decap_8
XFILLER_47_399 VDD VSS sg13g2_decap_8
XFILLER_16_742 VDD VSS sg13g2_decap_8
XFILLER_15_252 VDD VSS sg13g2_decap_8
XFILLER_95_7 VDD VSS sg13g2_decap_8
XFILLER_31_756 VDD VSS sg13g2_fill_1
XFILLER_30_266 VDD VSS sg13g2_decap_8
XFILLER_7_462 VDD VSS sg13g2_decap_8
XFILLER_85_406 VDD VSS sg13g2_decap_8
XFILLER_58_609 VDD VSS sg13g2_decap_8
XFILLER_38_322 VDD VSS sg13g2_decap_8
XFILLER_57_119 VDD VSS sg13g2_decap_8
XFILLER_66_653 VDD VSS sg13g2_decap_8
XFILLER_17_0 VDD VSS sg13g2_decap_8
XFILLER_93_483 VDD VSS sg13g2_decap_8
XFILLER_81_623 VDD VSS sg13g2_decap_8
XFILLER_26_517 VDD VSS sg13g2_decap_8
XFILLER_80_133 VDD VSS sg13g2_decap_8
XFILLER_65_196 VDD VSS sg13g2_decap_8
XFILLER_0_70 VDD VSS sg13g2_decap_8
XFILLER_38_399 VDD VSS sg13g2_decap_8
XFILLER_53_336 VDD VSS sg13g2_decap_8
XFILLER_22_756 VDD VSS sg13g2_fill_1
XFILLER_21_266 VDD VSS sg13g2_decap_8
XFILLER_1_616 VDD VSS sg13g2_decap_8
XFILLER_89_756 VDD VSS sg13g2_fill_1
XFILLER_0_126 VDD VSS sg13g2_decap_8
XFILLER_88_266 VDD VSS sg13g2_decap_8
XFILLER_95_28 VDD VSS sg13g2_decap_8
XFILLER_49_609 VDD VSS sg13g2_decap_8
XFILLER_48_119 VDD VSS sg13g2_decap_8
XFILLER_29_322 VDD VSS sg13g2_decap_8
XFILLER_84_483 VDD VSS sg13g2_decap_8
XFILLER_57_686 VDD VSS sg13g2_decap_8
XFILLER_28_77 VDD VSS sg13g2_decap_8
XFILLER_72_656 VDD VSS sg13g2_decap_8
XFILLER_71_133 VDD VSS sg13g2_decap_8
XFILLER_29_399 VDD VSS sg13g2_decap_8
XFILLER_44_336 VDD VSS sg13g2_decap_8
XFILLER_56_196 VDD VSS sg13g2_decap_8
XFILLER_17_539 VDD VSS sg13g2_decap_8
XFILLER_44_21 VDD VSS sg13g2_decap_8
XFILLER_13_756 VDD VSS sg13g2_fill_1
XFILLER_44_98 VDD VSS sg13g2_decap_8
XFILLER_40_553 VDD VSS sg13g2_decap_8
XFILLER_9_749 VDD VSS sg13g2_decap_8
XFILLER_12_266 VDD VSS sg13g2_decap_8
XFILLER_8_259 VDD VSS sg13g2_decap_8
XFILLER_60_42 VDD VSS sg13g2_decap_8
XFILLER_4_476 VDD VSS sg13g2_decap_8
XFILLER_69_84 VDD VSS sg13g2_decap_8
XFILLER_79_266 VDD VSS sg13g2_decap_8
XFILLER_94_203 VDD VSS sg13g2_decap_8
XFILLER_39_119 VDD VSS sg13g2_decap_8
XFILLER_0_693 VDD VSS sg13g2_decap_8
XFILLER_10_7 VDD VSS sg13g2_decap_8
XFILLER_48_686 VDD VSS sg13g2_decap_8
XFILLER_75_494 VDD VSS sg13g2_decap_8
XFILLER_63_634 VDD VSS sg13g2_decap_8
XFILLER_90_420 VDD VSS sg13g2_decap_8
XFILLER_62_133 VDD VSS sg13g2_decap_8
XFILLER_35_336 VDD VSS sg13g2_decap_8
XFILLER_47_196 VDD VSS sg13g2_decap_8
XFILLER_90_497 VDD VSS sg13g2_decap_8
XFILLER_31_553 VDD VSS sg13g2_decap_8
XFILLER_58_406 VDD VSS sg13g2_decap_8
XFILLER_85_203 VDD VSS sg13g2_decap_8
XFILLER_39_686 VDD VSS sg13g2_decap_8
XFILLER_93_280 VDD VSS sg13g2_decap_8
XFILLER_81_420 VDD VSS sg13g2_decap_8
XFILLER_54_623 VDD VSS sg13g2_decap_8
XFILLER_26_314 VDD VSS sg13g2_decap_8
XFILLER_38_196 VDD VSS sg13g2_decap_8
XFILLER_53_133 VDD VSS sg13g2_decap_8
XFILLER_81_497 VDD VSS sg13g2_decap_8
XFILLER_14_35 VDD VSS sg13g2_decap_8
XFILLER_22_553 VDD VSS sg13g2_decap_8
XFILLER_30_56 VDD VSS sg13g2_decap_8
XFILLER_1_413 VDD VSS sg13g2_decap_8
XFILLER_89_553 VDD VSS sg13g2_decap_8
XFILLER_39_21 VDD VSS sg13g2_decap_8
XFILLER_49_406 VDD VSS sg13g2_decap_8
XFILLER_77_737 VDD VSS sg13g2_decap_8
XFILLER_76_203 VDD VSS sg13g2_decap_8
XFILLER_92_707 VDD VSS sg13g2_decap_8
XFILLER_39_98 VDD VSS sg13g2_decap_8
XFILLER_91_217 VDD VSS sg13g2_decap_8
XFILLER_84_280 VDD VSS sg13g2_decap_8
XFILLER_57_483 VDD VSS sg13g2_decap_8
XFILLER_55_42 VDD VSS sg13g2_decap_8
XFILLER_17_336 VDD VSS sg13g2_decap_8
XFILLER_29_196 VDD VSS sg13g2_decap_8
XFILLER_45_623 VDD VSS sg13g2_decap_8
XFILLER_72_453 VDD VSS sg13g2_decap_8
XFILLER_44_133 VDD VSS sg13g2_decap_8
XFILLER_60_637 VDD VSS sg13g2_decap_8
XFILLER_13_553 VDD VSS sg13g2_decap_8
XFILLER_71_63 VDD VSS sg13g2_decap_8
XFILLER_40_350 VDD VSS sg13g2_decap_8
XFILLER_9_546 VDD VSS sg13g2_decap_8
Xoutputs\[5\].output_pad _81_/Q IOVDD IOVSS output_PAD[5] VDD VSS sg13g2_IOPadOut30mA
XFILLER_58_7 VDD VSS sg13g2_decap_8
XFILLER_4_273 VDD VSS sg13g2_decap_8
XFILLER_68_748 VDD VSS sg13g2_decap_8
XFILLER_95_567 VDD VSS sg13g2_decap_8
XFILLER_83_707 VDD VSS sg13g2_decap_8
XFILLER_67_247 VDD VSS sg13g2_decap_8
XFILLER_0_490 VDD VSS sg13g2_decap_8
XFILLER_82_217 VDD VSS sg13g2_decap_8
XFILLER_63_420 VDD VSS sg13g2_decap_8
XFILLER_48_483 VDD VSS sg13g2_decap_8
XFILLER_36_623 VDD VSS sg13g2_decap_8
XFILLER_35_133 VDD VSS sg13g2_decap_8
XFILLER_51_637 VDD VSS sg13g2_decap_8
XFILLER_90_294 VDD VSS sg13g2_decap_8
XFILLER_50_147 VDD VSS sg13g2_decap_8
XFILLER_31_350 VDD VSS sg13g2_decap_8
XFILLER_84_0 VDD VSS sg13g2_decap_8
XFILLER_6_91 VDD VSS sg13g2_decap_8
XFILLER_58_203 VDD VSS sg13g2_decap_8
XFILLER_86_567 VDD VSS sg13g2_decap_8
XFILLER_74_707 VDD VSS sg13g2_decap_8
XFILLER_73_217 VDD VSS sg13g2_decap_8
XFILLER_66_280 VDD VSS sg13g2_decap_8
XFILLER_54_420 VDD VSS sg13g2_decap_8
XFILLER_27_623 VDD VSS sg13g2_decap_8
XFILLER_39_483 VDD VSS sg13g2_decap_8
XFILLER_26_133 VDD VSS sg13g2_decap_8
XFILLER_54_497 VDD VSS sg13g2_decap_8
XFILLER_42_637 VDD VSS sg13g2_decap_8
XFILLER_81_294 VDD VSS sg13g2_decap_8
XFILLER_25_56 VDD VSS sg13g2_decap_8
XFILLER_41_147 VDD VSS sg13g2_decap_8
XFILLER_22_350 VDD VSS sg13g2_decap_8
XFILLER_10_567 VDD VSS sg13g2_decap_8
XFILLER_41_77 VDD VSS sg13g2_decap_8
XFILLER_2_700 VDD VSS sg13g2_decap_8
XFILLER_1_210 VDD VSS sg13g2_decap_8
XFILLER_89_350 VDD VSS sg13g2_decap_8
XFILLER_49_203 VDD VSS sg13g2_decap_8
XFILLER_77_534 VDD VSS sg13g2_decap_8
XFILLER_2_49 VDD VSS sg13g2_decap_8
XFILLER_1_287 VDD VSS sg13g2_decap_8
XFILLER_92_504 VDD VSS sg13g2_decap_8
XFILLER_66_63 VDD VSS sg13g2_decap_8
XFILLER_64_217 VDD VSS sg13g2_decap_8
XFILLER_45_420 VDD VSS sg13g2_decap_8
XFILLER_57_280 VDD VSS sg13g2_decap_8
XFILLER_18_623 VDD VSS sg13g2_decap_8
XFILLER_73_751 VDD VSS sg13g2_decap_4
XFILLER_17_133 VDD VSS sg13g2_decap_8
XFILLER_33_637 VDD VSS sg13g2_decap_8
XFILLER_45_497 VDD VSS sg13g2_decap_8
XFILLER_72_294 VDD VSS sg13g2_decap_8
XFILLER_82_84 VDD VSS sg13g2_decap_8
XFILLER_32_147 VDD VSS sg13g2_decap_8
XFILLER_60_434 VDD VSS sg13g2_decap_8
XFILLER_13_350 VDD VSS sg13g2_decap_8
XFILLER_9_343 VDD VSS sg13g2_decap_8
XFILLER_5_560 VDD VSS sg13g2_decap_8
XFILLER_68_545 VDD VSS sg13g2_decap_8
XFILLER_83_504 VDD VSS sg13g2_decap_8
XFILLER_95_364 VDD VSS sg13g2_decap_8
XFILLER_56_707 VDD VSS sg13g2_decap_8
XFILLER_36_420 VDD VSS sg13g2_decap_8
XFILLER_48_280 VDD VSS sg13g2_decap_8
XFILLER_55_217 VDD VSS sg13g2_decap_8
XFILLER_70_209 VDD VSS sg13g2_fill_2
XFILLER_91_581 VDD VSS sg13g2_decap_8
XFILLER_24_637 VDD VSS sg13g2_decap_8
XFILLER_36_497 VDD VSS sg13g2_decap_8
XFILLER_63_294 VDD VSS sg13g2_decap_8
XFILLER_23_147 VDD VSS sg13g2_decap_8
XFILLER_51_434 VDD VSS sg13g2_decap_8
XFILLER_11_14 VDD VSS sg13g2_decap_8
XFILLER_74_504 VDD VSS sg13g2_decap_8
XFILLER_86_364 VDD VSS sg13g2_decap_8
XFILLER_59_567 VDD VSS sg13g2_decap_8
XFILLER_47_707 VDD VSS sg13g2_decap_8
XFILLER_27_420 VDD VSS sg13g2_decap_8
XFILLER_39_280 VDD VSS sg13g2_decap_8
XFILLER_46_217 VDD VSS sg13g2_decap_8
XFILLER_82_581 VDD VSS sg13g2_decap_8
XFILLER_36_77 VDD VSS sg13g2_decap_8
XFILLER_70_743 VDD VSS sg13g2_decap_8
XFILLER_42_434 VDD VSS sg13g2_decap_8
XFILLER_54_294 VDD VSS sg13g2_decap_8
XFILLER_15_637 VDD VSS sg13g2_decap_8
XFILLER_27_497 VDD VSS sg13g2_decap_8
XFILLER_52_21 VDD VSS sg13g2_decap_8
XFILLER_14_147 VDD VSS sg13g2_decap_8
XFILLER_52_98 VDD VSS sg13g2_decap_8
XFILLER_10_364 VDD VSS sg13g2_decap_8
XFILLER_6_357 VDD VSS sg13g2_decap_8
XFILLER_2_574 VDD VSS sg13g2_decap_8
XFILLER_77_84 VDD VSS sg13g2_decap_8
Xinputs\[2\].input_pad IOVDD IOVSS _49_/D input_PAD[2] VDD VSS sg13g2_IOPadIn
XFILLER_38_707 VDD VSS sg13g2_decap_8
XFILLER_92_301 VDD VSS sg13g2_decap_8
XFILLER_77_386 VDD VSS sg13g2_decap_8
XFILLER_37_217 VDD VSS sg13g2_decap_8
XFILLER_18_420 VDD VSS sg13g2_decap_8
XFILLER_80_518 VDD VSS sg13g2_decap_8
XFILLER_92_378 VDD VSS sg13g2_decap_8
XFILLER_61_721 VDD VSS sg13g2_decap_8
XFILLER_33_434 VDD VSS sg13g2_decap_8
XFILLER_45_294 VDD VSS sg13g2_decap_8
XFILLER_60_231 VDD VSS sg13g2_decap_8
XFILLER_18_497 VDD VSS sg13g2_decap_8
XFILLER_9_140 VDD VSS sg13g2_decap_8
XFILLER_47_0 VDD VSS sg13g2_decap_8
XFILLER_68_342 VDD VSS sg13g2_decap_8
XFILLER_56_504 VDD VSS sg13g2_decap_8
XFILLER_3_70 VDD VSS sg13g2_decap_8
XFILLER_29_707 VDD VSS sg13g2_decap_8
XFILLER_95_161 VDD VSS sg13g2_decap_8
XFILLER_83_301 VDD VSS sg13g2_decap_8
XFILLER_28_217 VDD VSS sg13g2_decap_8
XFILLER_83_378 VDD VSS sg13g2_decap_8
XFILLER_52_721 VDD VSS sg13g2_decap_8
XFILLER_64_581 VDD VSS sg13g2_decap_8
XFILLER_24_434 VDD VSS sg13g2_decap_8
XFILLER_36_294 VDD VSS sg13g2_decap_8
XFILLER_51_231 VDD VSS sg13g2_decap_8
XFILLER_20_651 VDD VSS sg13g2_decap_8
XFILLER_22_35 VDD VSS sg13g2_decap_8
XFILLER_87_651 VDD VSS sg13g2_decap_8
XFILLER_47_504 VDD VSS sg13g2_decap_8
XFILLER_47_21 VDD VSS sg13g2_decap_8
XFILLER_59_364 VDD VSS sg13g2_decap_8
XFILLER_86_161 VDD VSS sg13g2_decap_8
XFILLER_74_323 VDD VSS sg13g2_decap_8
XFILLER_19_217 VDD VSS sg13g2_decap_8
XFILLER_47_98 VDD VSS sg13g2_decap_8
XFILLER_62_518 VDD VSS sg13g2_decap_8
XFILLER_74_378 VDD VSS sg13g2_fill_2
XFILLER_63_42 VDD VSS sg13g2_decap_8
XFILLER_55_581 VDD VSS sg13g2_decap_8
XFILLER_15_434 VDD VSS sg13g2_decap_8
XFILLER_27_294 VDD VSS sg13g2_decap_8
XFILLER_43_721 VDD VSS sg13g2_decap_8
XFILLER_70_540 VDD VSS sg13g2_decap_8
XFILLER_42_231 VDD VSS sg13g2_decap_8
XFILLER_11_651 VDD VSS sg13g2_decap_8
XFILLER_30_448 VDD VSS sg13g2_decap_8
XFILLER_10_161 VDD VSS sg13g2_decap_8
XFILLER_7_644 VDD VSS sg13g2_decap_8
XFILLER_6_154 VDD VSS sg13g2_decap_8
XFILLER_40_7 VDD VSS sg13g2_decap_8
XFILLER_2_371 VDD VSS sg13g2_decap_8
XFILLER_78_651 VDD VSS sg13g2_decap_8
XFILLER_38_504 VDD VSS sg13g2_decap_8
XFILLER_77_161 VDD VSS sg13g2_decap_8
XFILLER_65_301 VDD VSS sg13g2_decap_8
XFILLER_93_665 VDD VSS sg13g2_decap_8
XFILLER_92_175 VDD VSS sg13g2_decap_8
XFILLER_80_315 VDD VSS sg13g2_decap_8
XFILLER_65_378 VDD VSS sg13g2_decap_8
XFILLER_53_518 VDD VSS sg13g2_decap_8
XFILLER_46_581 VDD VSS sg13g2_decap_8
XFILLER_18_294 VDD VSS sg13g2_decap_8
XFILLER_34_721 VDD VSS sg13g2_decap_8
XFILLER_33_231 VDD VSS sg13g2_decap_8
XFILLER_61_595 VDD VSS sg13g2_decap_8
XFILLER_21_448 VDD VSS sg13g2_decap_8
XFILLER_0_308 VDD VSS sg13g2_decap_8
XFILLER_88_448 VDD VSS sg13g2_decap_8
XFILLER_75_109 VDD VSS sg13g2_decap_8
XFILLER_29_504 VDD VSS sg13g2_decap_8
XFILLER_68_161 VDD VSS sg13g2_decap_8
XFILLER_56_301 VDD VSS sg13g2_decap_8
XFILLER_84_665 VDD VSS sg13g2_decap_8
XFILLER_83_175 VDD VSS sg13g2_decap_8
XFILLER_17_35 VDD VSS sg13g2_decap_8
XFILLER_56_378 VDD VSS sg13g2_decap_8
XFILLER_44_518 VDD VSS sg13g2_decap_8
XFILLER_25_721 VDD VSS sg13g2_decap_8
XFILLER_37_581 VDD VSS sg13g2_decap_8
XFILLER_71_359 VDD VSS sg13g2_fill_2
XFILLER_24_231 VDD VSS sg13g2_decap_8
XFILLER_52_595 VDD VSS sg13g2_decap_8
XFILLER_40_735 VDD VSS sg13g2_decap_8
XFILLER_12_448 VDD VSS sg13g2_decap_8
XFILLER_33_56 VDD VSS sg13g2_decap_8
XFILLER_4_658 VDD VSS sg13g2_decap_8
XFILLER_3_168 VDD VSS sg13g2_decap_8
XFILLER_79_448 VDD VSS sg13g2_decap_8
XFILLER_58_42 VDD VSS sg13g2_decap_8
XFILLER_47_301 VDD VSS sg13g2_decap_8
XFILLER_59_161 VDD VSS sg13g2_decap_8
XFILLER_90_602 VDD VSS sg13g2_decap_8
XFILLER_75_676 VDD VSS sg13g2_decap_8
XFILLER_74_175 VDD VSS sg13g2_decap_8
XFILLER_62_315 VDD VSS sg13g2_decap_8
XFILLER_47_378 VDD VSS sg13g2_decap_8
XFILLER_35_518 VDD VSS sg13g2_decap_8
XFILLER_74_63 VDD VSS sg13g2_decap_8
XFILLER_16_721 VDD VSS sg13g2_decap_8
XFILLER_28_581 VDD VSS sg13g2_decap_8
XFILLER_90_679 VDD VSS sg13g2_decap_8
XFILLER_15_231 VDD VSS sg13g2_decap_8
XFILLER_31_735 VDD VSS sg13g2_decap_8
XFILLER_43_595 VDD VSS sg13g2_decap_8
XFILLER_88_7 VDD VSS sg13g2_decap_8
XFILLER_30_245 VDD VSS sg13g2_decap_8
XFILLER_90_84 VDD VSS sg13g2_decap_8
XFILLER_7_441 VDD VSS sg13g2_decap_8
XFILLER_38_301 VDD VSS sg13g2_decap_8
XFILLER_66_632 VDD VSS sg13g2_decap_8
XFILLER_81_602 VDD VSS sg13g2_decap_8
XFILLER_93_462 VDD VSS sg13g2_decap_8
XFILLER_38_378 VDD VSS sg13g2_decap_8
XFILLER_53_315 VDD VSS sg13g2_decap_8
XFILLER_80_112 VDD VSS sg13g2_decap_8
XFILLER_65_175 VDD VSS sg13g2_decap_8
XFILLER_19_581 VDD VSS sg13g2_decap_8
XFILLER_81_679 VDD VSS sg13g2_decap_8
XFILLER_80_189 VDD VSS sg13g2_decap_8
XFILLER_22_735 VDD VSS sg13g2_decap_8
XFILLER_34_595 VDD VSS sg13g2_decap_8
XFILLER_21_245 VDD VSS sg13g2_decap_8
XFILLER_61_392 VDD VSS sg13g2_decap_8
XFILLER_9_91 VDD VSS sg13g2_decap_8
XFILLER_89_735 VDD VSS sg13g2_decap_8
XFILLER_0_105 VDD VSS sg13g2_decap_8
XFILLER_88_245 VDD VSS sg13g2_decap_8
XFILLER_29_301 VDD VSS sg13g2_decap_8
XFILLER_28_56 VDD VSS sg13g2_decap_8
XFILLER_84_462 VDD VSS sg13g2_decap_8
XFILLER_57_665 VDD VSS sg13g2_decap_8
XFILLER_29_378 VDD VSS sg13g2_decap_8
XFILLER_17_518 VDD VSS sg13g2_decap_8
XFILLER_72_635 VDD VSS sg13g2_decap_8
XFILLER_71_112 VDD VSS sg13g2_decap_8
XFILLER_44_315 VDD VSS sg13g2_decap_8
XFILLER_56_175 VDD VSS sg13g2_decap_8
XFILLER_71_189 VDD VSS sg13g2_decap_8
XFILLER_13_735 VDD VSS sg13g2_decap_8
XFILLER_44_77 VDD VSS sg13g2_decap_8
XFILLER_25_595 VDD VSS sg13g2_decap_8
XFILLER_12_245 VDD VSS sg13g2_decap_8
XFILLER_52_392 VDD VSS sg13g2_decap_8
XFILLER_40_532 VDD VSS sg13g2_decap_8
XFILLER_9_728 VDD VSS sg13g2_decap_8
XFILLER_60_21 VDD VSS sg13g2_decap_8
XFILLER_8_238 VDD VSS sg13g2_decap_8
XFILLER_60_98 VDD VSS sg13g2_decap_8
XFILLER_4_455 VDD VSS sg13g2_decap_8
XFILLER_5_49 VDD VSS sg13g2_decap_8
XFILLER_69_63 VDD VSS sg13g2_decap_8
XFILLER_79_245 VDD VSS sg13g2_decap_8
XFILLER_95_749 VDD VSS sg13g2_decap_8
XFILLER_67_429 VDD VSS sg13g2_decap_8
XFILLER_0_672 VDD VSS sg13g2_decap_8
XFILLER_94_259 VDD VSS sg13g2_decap_8
XFILLER_63_613 VDD VSS sg13g2_decap_8
XFILLER_75_473 VDD VSS sg13g2_decap_8
XFILLER_75_451 VDD VSS sg13g2_decap_4
XFILLER_85_84 VDD VSS sg13g2_decap_8
XFILLER_48_665 VDD VSS sg13g2_decap_8
XFILLER_62_112 VDD VSS sg13g2_decap_8
XFILLER_35_315 VDD VSS sg13g2_decap_8
XFILLER_47_175 VDD VSS sg13g2_decap_8
XFILLER_90_476 VDD VSS sg13g2_decap_8
XFILLER_62_189 VDD VSS sg13g2_decap_8
XFILLER_50_329 VDD VSS sg13g2_decap_8
XFILLER_43_392 VDD VSS sg13g2_decap_8
XFILLER_16_595 VDD VSS sg13g2_decap_8
XFILLER_31_532 VDD VSS sg13g2_decap_8
XFILLER_86_749 VDD VSS sg13g2_decap_8
XFILLER_85_259 VDD VSS sg13g2_decap_8
XFILLER_54_602 VDD VSS sg13g2_decap_8
XFILLER_39_665 VDD VSS sg13g2_decap_8
XFILLER_38_175 VDD VSS sg13g2_decap_8
XFILLER_53_112 VDD VSS sg13g2_decap_8
XFILLER_54_679 VDD VSS sg13g2_decap_8
XFILLER_81_476 VDD VSS sg13g2_decap_8
XFILLER_41_329 VDD VSS sg13g2_decap_8
XFILLER_53_189 VDD VSS sg13g2_decap_8
XFILLER_14_14 VDD VSS sg13g2_decap_8
XFILLER_34_392 VDD VSS sg13g2_decap_8
XFILLER_22_532 VDD VSS sg13g2_decap_8
XFILLER_10_749 VDD VSS sg13g2_decap_8
XFILLER_30_35 VDD VSS sg13g2_decap_8
XFILLER_89_532 VDD VSS sg13g2_decap_8
XFILLER_77_716 VDD VSS sg13g2_decap_8
XFILLER_1_469 VDD VSS sg13g2_decap_8
XFILLER_39_77 VDD VSS sg13g2_decap_8
XFILLER_57_462 VDD VSS sg13g2_decap_8
XFILLER_45_602 VDD VSS sg13g2_decap_8
XFILLER_55_21 VDD VSS sg13g2_decap_8
XFILLER_17_315 VDD VSS sg13g2_decap_8
XFILLER_29_175 VDD VSS sg13g2_decap_8
XFILLER_44_112 VDD VSS sg13g2_decap_8
XFILLER_45_679 VDD VSS sg13g2_decap_8
XFILLER_60_616 VDD VSS sg13g2_decap_8
XFILLER_55_98 VDD VSS sg13g2_decap_8
XFILLER_32_329 VDD VSS sg13g2_decap_8
XFILLER_44_189 VDD VSS sg13g2_decap_8
XFILLER_13_532 VDD VSS sg13g2_decap_8
XFILLER_25_392 VDD VSS sg13g2_decap_8
XFILLER_71_42 VDD VSS sg13g2_decap_8
XFILLER_9_525 VDD VSS sg13g2_decap_8
XFILLER_5_742 VDD VSS sg13g2_decap_8
XFILLER_4_252 VDD VSS sg13g2_decap_8
XFILLER_68_727 VDD VSS sg13g2_decap_8
XFILLER_95_546 VDD VSS sg13g2_decap_8
Xclkbuf_1_0__f_clk_PAD2CORE _79_/CLK clkbuf_0_clk_PAD2CORE/X VDD VSS sg13g2_buf_16
XFILLER_67_226 VDD VSS sg13g2_decap_8
XFILLER_48_462 VDD VSS sg13g2_decap_8
XFILLER_36_602 VDD VSS sg13g2_decap_8
XFILLER_35_112 VDD VSS sg13g2_decap_8
XFILLER_36_679 VDD VSS sg13g2_decap_8
XFILLER_63_487 VDD VSS sg13g2_decap_8
XFILLER_90_273 VDD VSS sg13g2_decap_8
XFILLER_51_616 VDD VSS sg13g2_decap_8
XFILLER_23_329 VDD VSS sg13g2_decap_8
XFILLER_35_189 VDD VSS sg13g2_decap_8
XFILLER_16_392 VDD VSS sg13g2_decap_8
XFILLER_50_126 VDD VSS sg13g2_decap_8
XFILLER_77_0 VDD VSS sg13g2_decap_8
XFILLER_6_70 VDD VSS sg13g2_decap_8
XFILLER_86_546 VDD VSS sg13g2_decap_8
XFILLER_59_749 VDD VSS sg13g2_decap_8
XFILLER_39_462 VDD VSS sg13g2_decap_8
XFILLER_58_259 VDD VSS sg13g2_decap_8
XFILLER_27_602 VDD VSS sg13g2_decap_8
XFILLER_26_112 VDD VSS sg13g2_decap_8
XFILLER_27_679 VDD VSS sg13g2_decap_8
XFILLER_81_273 VDD VSS sg13g2_decap_8
XFILLER_25_35 VDD VSS sg13g2_decap_8
XFILLER_14_329 VDD VSS sg13g2_decap_8
XFILLER_26_189 VDD VSS sg13g2_decap_8
XFILLER_54_476 VDD VSS sg13g2_decap_8
XFILLER_42_616 VDD VSS sg13g2_decap_8
XFILLER_41_126 VDD VSS sg13g2_decap_8
XFILLER_50_693 VDD VSS sg13g2_decap_8
XFILLER_10_546 VDD VSS sg13g2_decap_8
XFILLER_41_56 VDD VSS sg13g2_decap_8
XFILLER_6_539 VDD VSS sg13g2_decap_8
XFILLER_2_756 VDD VSS sg13g2_fill_1
XFILLER_77_513 VDD VSS sg13g2_decap_8
XFILLER_1_266 VDD VSS sg13g2_decap_8
Xinputs\[1\].input_pad IOVDD IOVSS hold14/A input_PAD[1] VDD VSS sg13g2_IOPadIn
XFILLER_2_28 VDD VSS sg13g2_decap_8
XFILLER_66_42 VDD VSS sg13g2_decap_8
XFILLER_49_259 VDD VSS sg13g2_decap_8
XFILLER_18_602 VDD VSS sg13g2_decap_8
XFILLER_73_730 VDD VSS sg13g2_decap_8
XFILLER_17_112 VDD VSS sg13g2_decap_8
XFILLER_45_476 VDD VSS sg13g2_decap_8
XFILLER_60_413 VDD VSS sg13g2_decap_8
XFILLER_18_679 VDD VSS sg13g2_decap_8
XFILLER_33_616 VDD VSS sg13g2_decap_8
XFILLER_82_63 VDD VSS sg13g2_decap_8
XFILLER_17_189 VDD VSS sg13g2_decap_8
XFILLER_32_126 VDD VSS sg13g2_decap_8
XFILLER_9_322 VDD VSS sg13g2_decap_8
XFILLER_41_693 VDD VSS sg13g2_decap_8
XFILLER_70_7 VDD VSS sg13g2_decap_8
XFILLER_9_399 VDD VSS sg13g2_decap_8
XFILLER_68_524 VDD VSS sg13g2_decap_8
XFILLER_95_343 VDD VSS sg13g2_decap_8
XFILLER_91_560 VDD VSS sg13g2_decap_8
XFILLER_63_273 VDD VSS sg13g2_decap_8
XFILLER_36_476 VDD VSS sg13g2_decap_8
XFILLER_51_413 VDD VSS sg13g2_decap_8
XFILLER_24_616 VDD VSS sg13g2_decap_8
XFILLER_23_126 VDD VSS sg13g2_decap_8
XFILLER_32_693 VDD VSS sg13g2_decap_8
XFILLER_59_546 VDD VSS sg13g2_decap_8
XFILLER_86_343 VDD VSS sg13g2_decap_8
XFILLER_67_590 VDD VSS sg13g2_decap_8
XFILLER_82_560 VDD VSS sg13g2_decap_8
XFILLER_70_722 VDD VSS sg13g2_decap_8
XFILLER_36_56 VDD VSS sg13g2_decap_8
XFILLER_27_476 VDD VSS sg13g2_decap_8
XFILLER_42_413 VDD VSS sg13g2_decap_8
XFILLER_15_616 VDD VSS sg13g2_decap_8
XFILLER_14_126 VDD VSS sg13g2_decap_8
XFILLER_54_273 VDD VSS sg13g2_decap_8
XFILLER_23_693 VDD VSS sg13g2_decap_8
XFILLER_50_490 VDD VSS sg13g2_decap_8
XFILLER_10_343 VDD VSS sg13g2_decap_8
XFILLER_52_77 VDD VSS sg13g2_decap_8
XFILLER_6_336 VDD VSS sg13g2_decap_8
XFILLER_7_0 VDD VSS sg13g2_decap_8
XFILLER_2_553 VDD VSS sg13g2_decap_8
XFILLER_77_63 VDD VSS sg13g2_decap_8
XFILLER_77_365 VDD VSS sg13g2_decap_8
XFILLER_65_549 VDD VSS sg13g2_decap_8
XFILLER_92_357 VDD VSS sg13g2_decap_8
XFILLER_93_84 VDD VSS sg13g2_decap_8
XFILLER_61_700 VDD VSS sg13g2_decap_8
XFILLER_18_476 VDD VSS sg13g2_decap_8
XFILLER_33_413 VDD VSS sg13g2_decap_8
XFILLER_45_273 VDD VSS sg13g2_decap_8
XFILLER_60_210 VDD VSS sg13g2_decap_8
XFILLER_60_287 VDD VSS sg13g2_decap_8
XFILLER_14_693 VDD VSS sg13g2_decap_8
XFILLER_41_490 VDD VSS sg13g2_decap_8
XFILLER_9_196 VDD VSS sg13g2_decap_8
XFILLER_68_321 VDD VSS sg13g2_decap_8
XFILLER_95_140 VDD VSS sg13g2_decap_8
XFILLER_68_398 VDD VSS sg13g2_decap_8
XFILLER_83_357 VDD VSS sg13g2_decap_8
XFILLER_64_560 VDD VSS sg13g2_decap_8
XFILLER_52_700 VDD VSS sg13g2_decap_8
XFILLER_24_413 VDD VSS sg13g2_decap_8
XFILLER_36_273 VDD VSS sg13g2_decap_8
XFILLER_51_210 VDD VSS sg13g2_decap_8
XFILLER_51_287 VDD VSS sg13g2_decap_8
XFILLER_22_14 VDD VSS sg13g2_decap_8
XFILLER_20_630 VDD VSS sg13g2_decap_8
XFILLER_32_490 VDD VSS sg13g2_decap_8
XFILLER_0_7 VDD VSS sg13g2_decap_8
XFILLER_87_630 VDD VSS sg13g2_decap_8
XFILLER_86_140 VDD VSS sg13g2_decap_8
XFILLER_59_343 VDD VSS sg13g2_decap_8
XFILLER_74_302 VDD VSS sg13g2_decap_8
XFILLER_47_77 VDD VSS sg13g2_decap_8
XFILLER_55_560 VDD VSS sg13g2_decap_8
XFILLER_43_700 VDD VSS sg13g2_decap_8
XFILLER_63_21 VDD VSS sg13g2_decap_8
XFILLER_15_413 VDD VSS sg13g2_decap_8
XFILLER_27_273 VDD VSS sg13g2_decap_8
XFILLER_42_210 VDD VSS sg13g2_decap_8
XFILLER_70_596 VDD VSS sg13g2_decap_8
XFILLER_63_98 VDD VSS sg13g2_decap_8
XFILLER_30_427 VDD VSS sg13g2_decap_8
XFILLER_42_287 VDD VSS sg13g2_decap_8
XFILLER_11_630 VDD VSS sg13g2_decap_8
XFILLER_8_49 VDD VSS sg13g2_decap_8
XFILLER_23_490 VDD VSS sg13g2_decap_8
XFILLER_7_623 VDD VSS sg13g2_decap_8
XFILLER_10_140 VDD VSS sg13g2_decap_8
XFILLER_6_133 VDD VSS sg13g2_decap_8
XFILLER_12_91 VDD VSS sg13g2_decap_8
XFILLER_2_350 VDD VSS sg13g2_decap_8
XFILLER_78_630 VDD VSS sg13g2_decap_8
XFILLER_88_84 VDD VSS sg13g2_decap_8
XFILLER_33_7 VDD VSS sg13g2_decap_8
XFILLER_77_140 VDD VSS sg13g2_decap_8
XFILLER_93_644 VDD VSS sg13g2_decap_8
XFILLER_65_357 VDD VSS sg13g2_decap_8
XFILLER_92_154 VDD VSS sg13g2_decap_8
XFILLER_46_560 VDD VSS sg13g2_decap_8
XFILLER_34_700 VDD VSS sg13g2_decap_8
XFILLER_18_273 VDD VSS sg13g2_decap_8
XFILLER_33_210 VDD VSS sg13g2_decap_8
XFILLER_61_574 VDD VSS sg13g2_decap_8
XFILLER_21_427 VDD VSS sg13g2_decap_8
XFILLER_33_287 VDD VSS sg13g2_decap_8
XFILLER_14_490 VDD VSS sg13g2_decap_8
XFILLER_88_427 VDD VSS sg13g2_decap_8
XFILLER_68_140 VDD VSS sg13g2_decap_8
XFILLER_69_685 VDD VSS sg13g2_decap_8
XFILLER_84_644 VDD VSS sg13g2_decap_8
XFILLER_17_14 VDD VSS sg13g2_decap_8
XFILLER_83_154 VDD VSS sg13g2_decap_8
XFILLER_56_357 VDD VSS sg13g2_decap_8
XFILLER_25_700 VDD VSS sg13g2_decap_8
XFILLER_37_560 VDD VSS sg13g2_decap_8
XFILLER_71_338 VDD VSS sg13g2_decap_8
XFILLER_24_210 VDD VSS sg13g2_decap_8
XFILLER_52_574 VDD VSS sg13g2_decap_8
XFILLER_12_427 VDD VSS sg13g2_decap_8
XFILLER_24_287 VDD VSS sg13g2_decap_8
XFILLER_40_714 VDD VSS sg13g2_decap_8
XFILLER_33_35 VDD VSS sg13g2_decap_8
XFILLER_4_637 VDD VSS sg13g2_decap_8
XFILLER_3_147 VDD VSS sg13g2_decap_8
XFILLER_79_427 VDD VSS sg13g2_decap_8
XFILLER_58_21 VDD VSS sg13g2_decap_8
XFILLER_58_98 VDD VSS sg13g2_decap_8
XFILLER_59_140 VDD VSS sg13g2_decap_8
XFILLER_75_655 VDD VSS sg13g2_decap_8
XFILLER_74_154 VDD VSS sg13g2_decap_8
XFILLER_74_42 VDD VSS sg13g2_decap_8
XFILLER_47_357 VDD VSS sg13g2_decap_8
XFILLER_16_700 VDD VSS sg13g2_decap_8
XFILLER_28_560 VDD VSS sg13g2_decap_8
XFILLER_90_658 VDD VSS sg13g2_decap_8
XFILLER_15_210 VDD VSS sg13g2_decap_8
XFILLER_15_287 VDD VSS sg13g2_decap_8
XFILLER_31_714 VDD VSS sg13g2_decap_8
XFILLER_43_574 VDD VSS sg13g2_decap_8
XFILLER_90_63 VDD VSS sg13g2_decap_8
XFILLER_30_224 VDD VSS sg13g2_decap_8
XFILLER_7_420 VDD VSS sg13g2_decap_8
XFILLER_7_497 VDD VSS sg13g2_decap_8
XFILLER_66_611 VDD VSS sg13g2_decap_8
XFILLER_93_441 VDD VSS sg13g2_decap_8
XFILLER_66_688 VDD VSS sg13g2_decap_8
XFILLER_65_154 VDD VSS sg13g2_decap_8
XFILLER_38_357 VDD VSS sg13g2_decap_8
XFILLER_19_560 VDD VSS sg13g2_decap_8
XFILLER_81_658 VDD VSS sg13g2_decap_8
XFILLER_80_168 VDD VSS sg13g2_decap_8
XFILLER_61_371 VDD VSS sg13g2_decap_8
XFILLER_22_714 VDD VSS sg13g2_decap_8
XFILLER_34_574 VDD VSS sg13g2_decap_8
XFILLER_21_224 VDD VSS sg13g2_decap_8
XFILLER_9_70 VDD VSS sg13g2_decap_8
XFILLER_89_714 VDD VSS sg13g2_decap_8
XFILLER_88_224 VDD VSS sg13g2_decap_8
XFILLER_76_419 VDD VSS sg13g2_decap_8
XFILLER_57_644 VDD VSS sg13g2_decap_8
XFILLER_28_35 VDD VSS sg13g2_decap_8
XFILLER_72_614 VDD VSS sg13g2_decap_8
XFILLER_84_441 VDD VSS sg13g2_decap_8
XFILLER_29_357 VDD VSS sg13g2_decap_8
XFILLER_56_154 VDD VSS sg13g2_decap_8
XFILLER_71_168 VDD VSS sg13g2_decap_8
XFILLER_13_714 VDD VSS sg13g2_decap_8
XFILLER_44_56 VDD VSS sg13g2_decap_8
XFILLER_52_371 VDD VSS sg13g2_decap_8
XFILLER_25_574 VDD VSS sg13g2_decap_8
XFILLER_40_511 VDD VSS sg13g2_decap_8
XFILLER_9_707 VDD VSS sg13g2_decap_8
XFILLER_12_224 VDD VSS sg13g2_decap_8
XFILLER_8_217 VDD VSS sg13g2_decap_8
XFILLER_40_588 VDD VSS sg13g2_decap_8
XFILLER_60_77 VDD VSS sg13g2_decap_8
XFILLER_4_434 VDD VSS sg13g2_decap_8
XFILLER_5_28 VDD VSS sg13g2_decap_8
XFILLER_79_224 VDD VSS sg13g2_decap_8
XFILLER_69_42 VDD VSS sg13g2_decap_8
XFILLER_95_728 VDD VSS sg13g2_decap_8
XFILLER_67_408 VDD VSS sg13g2_decap_8
XFILLER_0_651 VDD VSS sg13g2_decap_8
XFILLER_94_238 VDD VSS sg13g2_decap_8
XFILLER_75_430 VDD VSS sg13g2_decap_8
XFILLER_48_644 VDD VSS sg13g2_decap_8
XFILLER_85_63 VDD VSS sg13g2_decap_8
XFILLER_47_154 VDD VSS sg13g2_decap_8
XFILLER_63_669 VDD VSS sg13g2_decap_8
XFILLER_90_455 VDD VSS sg13g2_decap_8
XFILLER_62_168 VDD VSS sg13g2_decap_8
XFILLER_43_371 VDD VSS sg13g2_decap_8
XFILLER_50_308 VDD VSS sg13g2_decap_8
XFILLER_16_574 VDD VSS sg13g2_decap_8
XFILLER_31_511 VDD VSS sg13g2_decap_8
XFILLER_31_588 VDD VSS sg13g2_decap_8
XFILLER_7_294 VDD VSS sg13g2_decap_8
XFILLER_86_728 VDD VSS sg13g2_decap_8
XFILLER_22_0 VDD VSS sg13g2_decap_8
XFILLER_85_238 VDD VSS sg13g2_decap_8
XFILLER_39_644 VDD VSS sg13g2_decap_8
XFILLER_66_441 VDD VSS sg13g2_decap_8
XFILLER_38_154 VDD VSS sg13g2_decap_8
XFILLER_66_485 VDD VSS sg13g2_decap_8
XFILLER_81_455 VDD VSS sg13g2_decap_8
XFILLER_54_658 VDD VSS sg13g2_decap_8
XFILLER_26_349 VDD VSS sg13g2_decap_8
XFILLER_41_308 VDD VSS sg13g2_decap_8
XFILLER_53_168 VDD VSS sg13g2_decap_8
XFILLER_34_371 VDD VSS sg13g2_decap_8
XFILLER_22_511 VDD VSS sg13g2_decap_8
XFILLER_10_728 VDD VSS sg13g2_decap_8
XFILLER_22_588 VDD VSS sg13g2_decap_8
XFILLER_30_14 VDD VSS sg13g2_decap_8
XFILLER_89_511 VDD VSS sg13g2_decap_8
XFILLER_1_448 VDD VSS sg13g2_decap_8
XFILLER_89_588 VDD VSS sg13g2_decap_8
Xinputs\[0\].input_pad IOVDD IOVSS _51_/A input_PAD[0] VDD VSS sg13g2_IOPadIn
XFILLER_39_56 VDD VSS sg13g2_decap_8
XFILLER_29_154 VDD VSS sg13g2_decap_8
XFILLER_57_441 VDD VSS sg13g2_decap_8
XFILLER_55_77 VDD VSS sg13g2_decap_8
XFILLER_45_658 VDD VSS sg13g2_decap_8
XFILLER_72_488 VDD VSS sg13g2_decap_8
XFILLER_32_308 VDD VSS sg13g2_decap_8
XFILLER_44_168 VDD VSS sg13g2_decap_8
XFILLER_71_21 VDD VSS sg13g2_decap_8
XFILLER_13_511 VDD VSS sg13g2_decap_8
XFILLER_25_371 VDD VSS sg13g2_decap_8
XFILLER_9_504 VDD VSS sg13g2_decap_8
XFILLER_71_98 VDD VSS sg13g2_decap_8
XFILLER_13_588 VDD VSS sg13g2_decap_8
XFILLER_40_385 VDD VSS sg13g2_decap_8
XFILLER_5_721 VDD VSS sg13g2_decap_8
XFILLER_4_231 VDD VSS sg13g2_decap_8
XFILLER_68_706 VDD VSS sg13g2_decap_8
XFILLER_20_91 VDD VSS sg13g2_decap_8
XFILLER_95_525 VDD VSS sg13g2_decap_8
XFILLER_48_441 VDD VSS sg13g2_decap_8
XFILLER_75_271 VDD VSS sg13g2_decap_8
XFILLER_75_282 VDD VSS sg13g2_fill_2
XFILLER_91_742 VDD VSS sg13g2_decap_8
XFILLER_36_658 VDD VSS sg13g2_decap_8
XFILLER_90_252 VDD VSS sg13g2_decap_8
XFILLER_50_105 VDD VSS sg13g2_decap_8
XFILLER_23_308 VDD VSS sg13g2_decap_8
XFILLER_35_168 VDD VSS sg13g2_decap_8
XFILLER_16_371 VDD VSS sg13g2_decap_8
XFILLER_31_385 VDD VSS sg13g2_decap_8
XFILLER_8_581 VDD VSS sg13g2_decap_8
XFILLER_59_728 VDD VSS sg13g2_decap_8
XFILLER_86_525 VDD VSS sg13g2_decap_8
XFILLER_58_238 VDD VSS sg13g2_decap_8
XFILLER_39_441 VDD VSS sg13g2_decap_8
XFILLER_82_742 VDD VSS sg13g2_decap_8
XFILLER_54_455 VDD VSS sg13g2_decap_8
XFILLER_27_658 VDD VSS sg13g2_decap_8
XFILLER_81_252 VDD VSS sg13g2_decap_8
XFILLER_25_14 VDD VSS sg13g2_decap_8
XFILLER_41_105 VDD VSS sg13g2_decap_8
XFILLER_14_308 VDD VSS sg13g2_decap_8
XFILLER_26_168 VDD VSS sg13g2_decap_8
XFILLER_50_672 VDD VSS sg13g2_decap_8
XFILLER_10_525 VDD VSS sg13g2_decap_8
XFILLER_22_385 VDD VSS sg13g2_decap_8
XFILLER_6_518 VDD VSS sg13g2_decap_8
XFILLER_41_35 VDD VSS sg13g2_decap_8
XFILLER_2_735 VDD VSS sg13g2_decap_8
XFILLER_1_245 VDD VSS sg13g2_decap_8
XFILLER_89_385 VDD VSS sg13g2_decap_8
XFILLER_49_238 VDD VSS sg13g2_decap_8
XFILLER_77_569 VDD VSS sg13g2_decap_8
XFILLER_66_21 VDD VSS sg13g2_decap_8
XFILLER_92_539 VDD VSS sg13g2_decap_8
XFILLER_66_98 VDD VSS sg13g2_decap_8
XFILLER_45_455 VDD VSS sg13g2_decap_8
XFILLER_18_658 VDD VSS sg13g2_decap_8
XFILLER_72_263 VDD VSS sg13g2_decap_8
XFILLER_32_105 VDD VSS sg13g2_decap_8
XFILLER_17_168 VDD VSS sg13g2_decap_8
XFILLER_82_42 VDD VSS sg13g2_decap_8
XFILLER_9_301 VDD VSS sg13g2_decap_8
XFILLER_60_469 VDD VSS sg13g2_decap_8
XFILLER_13_385 VDD VSS sg13g2_decap_8
XFILLER_15_91 VDD VSS sg13g2_decap_8
XFILLER_41_672 VDD VSS sg13g2_decap_8
XFILLER_40_182 VDD VSS sg13g2_decap_8
XFILLER_9_378 VDD VSS sg13g2_decap_8
XFILLER_63_7 VDD VSS sg13g2_decap_8
XFILLER_5_595 VDD VSS sg13g2_decap_8
XFILLER_68_503 VDD VSS sg13g2_decap_8
XFILLER_95_322 VDD VSS sg13g2_decap_8
XFILLER_83_539 VDD VSS sg13g2_decap_8
XFILLER_76_580 VDD VSS sg13g2_decap_8
XFILLER_95_399 VDD VSS sg13g2_decap_8
XFILLER_64_742 VDD VSS sg13g2_decap_8
XFILLER_63_252 VDD VSS sg13g2_decap_8
XFILLER_36_455 VDD VSS sg13g2_decap_8
XFILLER_23_105 VDD VSS sg13g2_decap_8
XFILLER_51_469 VDD VSS sg13g2_decap_8
XFILLER_32_672 VDD VSS sg13g2_decap_8
XFILLER_31_182 VDD VSS sg13g2_decap_8
XFILLER_11_49 VDD VSS sg13g2_decap_8
XFILLER_86_322 VDD VSS sg13g2_decap_8
XFILLER_59_525 VDD VSS sg13g2_decap_8
XFILLER_74_539 VDD VSS sg13g2_decap_8
XFILLER_86_399 VDD VSS sg13g2_decap_8
XFILLER_55_742 VDD VSS sg13g2_decap_8
XFILLER_36_35 VDD VSS sg13g2_decap_8
XFILLER_70_701 VDD VSS sg13g2_decap_8
XFILLER_27_455 VDD VSS sg13g2_decap_8
XFILLER_54_252 VDD VSS sg13g2_decap_8
XFILLER_14_105 VDD VSS sg13g2_decap_8
XFILLER_42_469 VDD VSS sg13g2_decap_8
XFILLER_30_609 VDD VSS sg13g2_decap_8
XFILLER_52_56 VDD VSS sg13g2_decap_8
XFILLER_23_672 VDD VSS sg13g2_decap_8
XFILLER_10_322 VDD VSS sg13g2_decap_8
XFILLER_22_182 VDD VSS sg13g2_decap_8
XFILLER_6_315 VDD VSS sg13g2_decap_8
XFILLER_10_399 VDD VSS sg13g2_decap_8
XFILLER_2_532 VDD VSS sg13g2_decap_8
XFILLER_89_182 VDD VSS sg13g2_decap_8
XFILLER_77_42 VDD VSS sg13g2_decap_8
XFILLER_77_344 VDD VSS sg13g2_decap_8
XFILLER_65_528 VDD VSS sg13g2_decap_8
XFILLER_92_336 VDD VSS sg13g2_decap_8
XFILLER_46_742 VDD VSS sg13g2_decap_8
XFILLER_93_63 VDD VSS sg13g2_decap_8
XFILLER_18_455 VDD VSS sg13g2_decap_8
XFILLER_45_252 VDD VSS sg13g2_decap_8
XFILLER_73_583 VDD VSS sg13g2_decap_8
XFILLER_61_756 VDD VSS sg13g2_fill_1
XFILLER_33_469 VDD VSS sg13g2_decap_8
XFILLER_21_609 VDD VSS sg13g2_decap_8
XFILLER_20_119 VDD VSS sg13g2_decap_8
XFILLER_60_266 VDD VSS sg13g2_decap_8
XFILLER_14_672 VDD VSS sg13g2_decap_8
XFILLER_13_182 VDD VSS sg13g2_decap_8
XFILLER_9_175 VDD VSS sg13g2_decap_8
XFILLER_5_392 VDD VSS sg13g2_decap_8
XFILLER_88_609 VDD VSS sg13g2_decap_8
XFILLER_87_119 VDD VSS sg13g2_decap_8
XFILLER_68_300 VDD VSS sg13g2_decap_8
XFILLER_68_377 VDD VSS sg13g2_decap_8
XFILLER_56_539 VDD VSS sg13g2_decap_8
XFILLER_95_196 VDD VSS sg13g2_decap_8
XFILLER_83_336 VDD VSS sg13g2_decap_8
XFILLER_37_742 VDD VSS sg13g2_decap_8
XFILLER_36_252 VDD VSS sg13g2_decap_8
XFILLER_52_756 VDD VSS sg13g2_fill_1
XFILLER_12_609 VDD VSS sg13g2_decap_8
XFILLER_24_469 VDD VSS sg13g2_decap_8
XFILLER_11_119 VDD VSS sg13g2_decap_8
XFILLER_51_266 VDD VSS sg13g2_decap_8
XFILLER_20_686 VDD VSS sg13g2_decap_8
XFILLER_3_329 VDD VSS sg13g2_decap_8
XFILLER_79_609 VDD VSS sg13g2_decap_8
XFILLER_78_119 VDD VSS sg13g2_decap_8
XFILLER_59_322 VDD VSS sg13g2_decap_8
XFILLER_87_686 VDD VSS sg13g2_decap_8
XFILLER_86_196 VDD VSS sg13g2_decap_8
XFILLER_47_539 VDD VSS sg13g2_decap_8
XFILLER_47_56 VDD VSS sg13g2_decap_8
XFILLER_59_399 VDD VSS sg13g2_decap_8
XFILLER_28_742 VDD VSS sg13g2_decap_8
XFILLER_27_252 VDD VSS sg13g2_decap_8
XFILLER_15_469 VDD VSS sg13g2_decap_8
XFILLER_43_756 VDD VSS sg13g2_fill_1
XFILLER_70_575 VDD VSS sg13g2_decap_8
XFILLER_63_77 VDD VSS sg13g2_decap_8
XFILLER_30_406 VDD VSS sg13g2_decap_8
XFILLER_42_266 VDD VSS sg13g2_decap_8
XFILLER_8_28 VDD VSS sg13g2_decap_8
XFILLER_7_602 VDD VSS sg13g2_decap_8
XFILLER_11_686 VDD VSS sg13g2_decap_8
XFILLER_6_112 VDD VSS sg13g2_decap_8
XFILLER_7_679 VDD VSS sg13g2_decap_8
XFILLER_10_196 VDD VSS sg13g2_decap_8
XFILLER_12_70 VDD VSS sg13g2_decap_8
XFILLER_6_189 VDD VSS sg13g2_decap_8
XFILLER_88_63 VDD VSS sg13g2_decap_8
XFILLER_69_119 VDD VSS sg13g2_decap_8
XFILLER_26_7 VDD VSS sg13g2_decap_8
XFILLER_93_623 VDD VSS sg13g2_decap_8
XFILLER_78_686 VDD VSS sg13g2_decap_8
XFILLER_92_133 VDD VSS sg13g2_decap_8
XFILLER_77_196 VDD VSS sg13g2_decap_8
XFILLER_65_336 VDD VSS sg13g2_decap_8
XFILLER_19_742 VDD VSS sg13g2_decap_8
XFILLER_38_539 VDD VSS sg13g2_decap_8
XFILLER_18_252 VDD VSS sg13g2_decap_8
XFILLER_61_553 VDD VSS sg13g2_decap_8
XFILLER_34_756 VDD VSS sg13g2_fill_1
XFILLER_21_406 VDD VSS sg13g2_decap_8
XFILLER_33_266 VDD VSS sg13g2_decap_8
XFILLER_52_0 VDD VSS sg13g2_decap_8
XFILLER_88_406 VDD VSS sg13g2_decap_8
XFILLER_84_623 VDD VSS sg13g2_decap_8
XFILLER_69_664 VDD VSS sg13g2_decap_8
XFILLER_83_133 VDD VSS sg13g2_decap_8
XFILLER_56_336 VDD VSS sg13g2_decap_8
XFILLER_29_539 VDD VSS sg13g2_decap_8
XFILLER_71_317 VDD VSS sg13g2_decap_8
XFILLER_52_553 VDD VSS sg13g2_decap_8
XFILLER_25_756 VDD VSS sg13g2_fill_1
XFILLER_12_406 VDD VSS sg13g2_decap_8
XFILLER_33_14 VDD VSS sg13g2_decap_8
XFILLER_24_266 VDD VSS sg13g2_decap_8
XFILLER_20_483 VDD VSS sg13g2_decap_8
XFILLER_4_616 VDD VSS sg13g2_decap_8
XFILLER_3_126 VDD VSS sg13g2_decap_8
XFILLER_79_406 VDD VSS sg13g2_decap_8
XFILLER_58_77 VDD VSS sg13g2_decap_8
XFILLER_87_483 VDD VSS sg13g2_decap_8
XFILLER_75_634 VDD VSS sg13g2_decap_8
XFILLER_47_336 VDD VSS sg13g2_decap_8
XFILLER_59_196 VDD VSS sg13g2_decap_8
XFILLER_74_133 VDD VSS sg13g2_decap_8
XFILLER_74_21 VDD VSS sg13g2_decap_8
XFILLER_90_637 VDD VSS sg13g2_decap_8
XFILLER_74_98 VDD VSS sg13g2_decap_8
XFILLER_43_553 VDD VSS sg13g2_decap_8
XFILLER_15_266 VDD VSS sg13g2_decap_8
XFILLER_30_203 VDD VSS sg13g2_decap_8
XFILLER_70_383 VDD VSS sg13g2_decap_8
XFILLER_90_42 VDD VSS sg13g2_decap_8
XFILLER_11_483 VDD VSS sg13g2_decap_8
XFILLER_23_91 VDD VSS sg13g2_decap_8
XFILLER_7_476 VDD VSS sg13g2_decap_8
XFILLER_3_693 VDD VSS sg13g2_decap_8
XFILLER_78_483 VDD VSS sg13g2_decap_8
XFILLER_93_420 VDD VSS sg13g2_decap_8
XFILLER_38_336 VDD VSS sg13g2_decap_8
XFILLER_66_667 VDD VSS sg13g2_decap_8
XFILLER_65_133 VDD VSS sg13g2_decap_8
Xoutputs\[8\].output_pad_1 VDD VSS outputs\[8\].output_pad/c2p sg13g2_tielo
XFILLER_93_497 VDD VSS sg13g2_decap_8
XFILLER_81_637 VDD VSS sg13g2_decap_8
XFILLER_80_147 VDD VSS sg13g2_decap_8
XFILLER_0_84 VDD VSS sg13g2_decap_8
XFILLER_34_553 VDD VSS sg13g2_decap_8
XFILLER_21_203 VDD VSS sg13g2_decap_8
XFILLER_61_350 VDD VSS sg13g2_decap_8
XFILLER_88_203 VDD VSS sg13g2_decap_8
XFILLER_28_14 VDD VSS sg13g2_decap_8
XFILLER_84_420 VDD VSS sg13g2_decap_8
XFILLER_57_623 VDD VSS sg13g2_decap_8
XFILLER_29_336 VDD VSS sg13g2_decap_8
XFILLER_56_133 VDD VSS sg13g2_decap_8
XFILLER_84_497 VDD VSS sg13g2_decap_8
XFILLER_71_147 VDD VSS sg13g2_decap_8
XFILLER_44_35 VDD VSS sg13g2_decap_8
XFILLER_12_203 VDD VSS sg13g2_decap_8
XFILLER_52_350 VDD VSS sg13g2_decap_8
XFILLER_25_553 VDD VSS sg13g2_decap_8
XFILLER_40_567 VDD VSS sg13g2_decap_8
XFILLER_60_56 VDD VSS sg13g2_decap_8
XFILLER_20_280 VDD VSS sg13g2_decap_8
XFILLER_4_413 VDD VSS sg13g2_decap_8
XFILLER_69_21 VDD VSS sg13g2_decap_8
XFILLER_79_203 VDD VSS sg13g2_decap_8
XFILLER_95_707 VDD VSS sg13g2_decap_8
XFILLER_69_98 VDD VSS sg13g2_decap_8
XFILLER_0_630 VDD VSS sg13g2_decap_8
XFILLER_94_217 VDD VSS sg13g2_decap_8
XFILLER_87_280 VDD VSS sg13g2_decap_8
XFILLER_85_42 VDD VSS sg13g2_decap_8
XFILLER_48_623 VDD VSS sg13g2_decap_8
XFILLER_47_133 VDD VSS sg13g2_decap_8
XFILLER_63_648 VDD VSS sg13g2_decap_8
XFILLER_90_434 VDD VSS sg13g2_decap_8
XFILLER_62_147 VDD VSS sg13g2_decap_8
XFILLER_18_91 VDD VSS sg13g2_decap_8
XFILLER_43_350 VDD VSS sg13g2_decap_8
XFILLER_16_553 VDD VSS sg13g2_decap_8
XFILLER_71_681 VDD VSS sg13g2_decap_8
XFILLER_93_7 VDD VSS sg13g2_decap_8
XFILLER_31_567 VDD VSS sg13g2_decap_8
XFILLER_11_280 VDD VSS sg13g2_decap_8
XFILLER_7_273 VDD VSS sg13g2_decap_8
XFILLER_86_707 VDD VSS sg13g2_decap_8
XFILLER_3_490 VDD VSS sg13g2_decap_8
XFILLER_85_217 VDD VSS sg13g2_decap_8
XFILLER_78_280 VDD VSS sg13g2_decap_8
XFILLER_66_420 VDD VSS sg13g2_decap_8
XFILLER_39_623 VDD VSS sg13g2_decap_8
XFILLER_66_464 VDD VSS sg13g2_decap_8
XFILLER_15_0 VDD VSS sg13g2_decap_8
XFILLER_38_133 VDD VSS sg13g2_decap_8
XFILLER_54_637 VDD VSS sg13g2_decap_8
XFILLER_26_328 VDD VSS sg13g2_decap_8
XFILLER_93_294 VDD VSS sg13g2_decap_8
XFILLER_81_434 VDD VSS sg13g2_decap_8
XFILLER_53_147 VDD VSS sg13g2_decap_8
XFILLER_34_350 VDD VSS sg13g2_decap_8
XFILLER_10_707 VDD VSS sg13g2_decap_8
XFILLER_14_49 VDD VSS sg13g2_decap_8
XFILLER_22_567 VDD VSS sg13g2_decap_8
XFILLER_1_427 VDD VSS sg13g2_decap_8
XFILLER_89_567 VDD VSS sg13g2_decap_8
XFILLER_39_35 VDD VSS sg13g2_decap_8
XFILLER_76_217 VDD VSS sg13g2_decap_8
XFILLER_76_228 VDD VSS sg13g2_fill_2
XFILLER_57_420 VDD VSS sg13g2_decap_8
XFILLER_29_133 VDD VSS sg13g2_decap_8
XFILLER_57_497 VDD VSS sg13g2_decap_8
XFILLER_45_637 VDD VSS sg13g2_decap_8
XFILLER_84_294 VDD VSS sg13g2_decap_8
XFILLER_72_434 VDD VSS sg13g2_fill_1
XFILLER_72_423 VDD VSS sg13g2_decap_8
XFILLER_55_56 VDD VSS sg13g2_decap_8
XFILLER_44_147 VDD VSS sg13g2_decap_8
XFILLER_72_467 VDD VSS sg13g2_decap_8
XFILLER_25_350 VDD VSS sg13g2_decap_8
XFILLER_13_567 VDD VSS sg13g2_decap_8
XFILLER_71_77 VDD VSS sg13g2_decap_8
XFILLER_40_364 VDD VSS sg13g2_decap_8
XFILLER_5_700 VDD VSS sg13g2_decap_8
XFILLER_4_210 VDD VSS sg13g2_decap_8
XFILLER_20_70 VDD VSS sg13g2_decap_8
XFILLER_4_287 VDD VSS sg13g2_decap_8
XFILLER_95_504 VDD VSS sg13g2_decap_8
XFILLER_48_420 VDD VSS sg13g2_decap_8
XFILLER_91_721 VDD VSS sg13g2_decap_8
XFILLER_75_250 VDD VSS sg13g2_decap_8
XFILLER_36_637 VDD VSS sg13g2_decap_8
XFILLER_90_231 VDD VSS sg13g2_decap_8
XFILLER_63_434 VDD VSS sg13g2_decap_8
XFILLER_48_497 VDD VSS sg13g2_decap_8
XFILLER_35_147 VDD VSS sg13g2_decap_8
XFILLER_16_350 VDD VSS sg13g2_decap_8
XFILLER_31_364 VDD VSS sg13g2_decap_8
XFILLER_8_560 VDD VSS sg13g2_decap_8
XFILLER_86_504 VDD VSS sg13g2_decap_8
XFILLER_59_707 VDD VSS sg13g2_decap_8
XFILLER_39_420 VDD VSS sg13g2_decap_8
XFILLER_58_217 VDD VSS sg13g2_decap_8
XFILLER_67_751 VDD VSS sg13g2_decap_4
XFILLER_94_581 VDD VSS sg13g2_decap_8
XFILLER_82_721 VDD VSS sg13g2_decap_8
XFILLER_81_231 VDD VSS sg13g2_decap_8
XFILLER_66_294 VDD VSS sg13g2_decap_8
XFILLER_54_434 VDD VSS sg13g2_decap_8
XFILLER_27_637 VDD VSS sg13g2_decap_8
XFILLER_39_497 VDD VSS sg13g2_decap_8
XFILLER_26_147 VDD VSS sg13g2_decap_8
XFILLER_50_651 VDD VSS sg13g2_decap_8
XFILLER_10_504 VDD VSS sg13g2_decap_8
XFILLER_41_14 VDD VSS sg13g2_decap_8
XFILLER_22_364 VDD VSS sg13g2_decap_8
XFILLER_2_714 VDD VSS sg13g2_decap_8
XFILLER_1_224 VDD VSS sg13g2_decap_8
XFILLER_89_364 VDD VSS sg13g2_decap_8
XFILLER_77_548 VDD VSS sg13g2_decap_8
XFILLER_49_217 VDD VSS sg13g2_decap_8
XIO_BOND_outputs\[3\].output_pad output_PAD[3] bondpad_70x70_novias
XFILLER_92_518 VDD VSS sg13g2_decap_8
XFILLER_85_581 VDD VSS sg13g2_decap_8
XFILLER_66_77 VDD VSS sg13g2_decap_8
XFILLER_45_434 VDD VSS sg13g2_decap_8
XFILLER_57_294 VDD VSS sg13g2_decap_8
XFILLER_18_637 VDD VSS sg13g2_decap_8
XFILLER_72_242 VDD VSS sg13g2_decap_8
XFILLER_82_21 VDD VSS sg13g2_decap_8
XFILLER_17_147 VDD VSS sg13g2_decap_8
XFILLER_26_692 VDD VSS sg13g2_decap_8
XFILLER_82_98 VDD VSS sg13g2_decap_8
XFILLER_60_448 VDD VSS sg13g2_decap_8
XFILLER_41_651 VDD VSS sg13g2_decap_8
XFILLER_13_364 VDD VSS sg13g2_decap_8
XFILLER_15_70 VDD VSS sg13g2_decap_8
XFILLER_40_161 VDD VSS sg13g2_decap_8
XFILLER_9_357 VDD VSS sg13g2_decap_8
XFILLER_5_574 VDD VSS sg13g2_decap_8
XFILLER_31_91 VDD VSS sg13g2_decap_8
XFILLER_56_7 VDD VSS sg13g2_decap_8
XFILLER_95_301 VDD VSS sg13g2_decap_8
XFILLER_68_559 VDD VSS sg13g2_decap_8
XFILLER_83_518 VDD VSS sg13g2_decap_8
XFILLER_95_378 VDD VSS sg13g2_decap_8
XFILLER_64_721 VDD VSS sg13g2_decap_8
XFILLER_36_434 VDD VSS sg13g2_decap_8
XFILLER_48_294 VDD VSS sg13g2_decap_8
XFILLER_63_231 VDD VSS sg13g2_decap_8
XFILLER_91_595 VDD VSS sg13g2_decap_8
XFILLER_51_448 VDD VSS sg13g2_decap_8
XFILLER_32_651 VDD VSS sg13g2_decap_8
XFILLER_31_161 VDD VSS sg13g2_decap_8
XFILLER_82_0 VDD VSS sg13g2_decap_8
XFILLER_11_28 VDD VSS sg13g2_decap_8
XFILLER_59_504 VDD VSS sg13g2_decap_8
XFILLER_86_301 VDD VSS sg13g2_decap_8
XFILLER_74_518 VDD VSS sg13g2_decap_8
XFILLER_86_378 VDD VSS sg13g2_decap_8
XFILLER_55_721 VDD VSS sg13g2_decap_8
XFILLER_36_14 VDD VSS sg13g2_decap_8
XFILLER_27_434 VDD VSS sg13g2_decap_8
XFILLER_39_294 VDD VSS sg13g2_decap_8
XFILLER_54_231 VDD VSS sg13g2_decap_8
XFILLER_82_595 VDD VSS sg13g2_decap_8
XFILLER_42_448 VDD VSS sg13g2_decap_8
XFILLER_23_651 VDD VSS sg13g2_decap_8
XFILLER_10_301 VDD VSS sg13g2_decap_8
XFILLER_52_35 VDD VSS sg13g2_decap_8
XFILLER_22_161 VDD VSS sg13g2_decap_8
XFILLER_10_378 VDD VSS sg13g2_decap_8
XFILLER_2_511 VDD VSS sg13g2_decap_8
XFILLER_77_21 VDD VSS sg13g2_decap_8
XFILLER_89_161 VDD VSS sg13g2_decap_8
XFILLER_77_323 VDD VSS sg13g2_decap_8
XFILLER_2_588 VDD VSS sg13g2_decap_8
XFILLER_65_507 VDD VSS sg13g2_decap_8
XFILLER_92_315 VDD VSS sg13g2_decap_8
XFILLER_77_98 VDD VSS sg13g2_decap_8
XFILLER_93_42 VDD VSS sg13g2_decap_8
XFILLER_58_581 VDD VSS sg13g2_decap_8
XFILLER_46_721 VDD VSS sg13g2_decap_8
XFILLER_18_434 VDD VSS sg13g2_decap_8
XFILLER_73_562 VDD VSS sg13g2_decap_8
XFILLER_45_231 VDD VSS sg13g2_decap_8
XFILLER_61_735 VDD VSS sg13g2_decap_8
XFILLER_26_91 VDD VSS sg13g2_decap_8
XFILLER_33_448 VDD VSS sg13g2_decap_8
XFILLER_60_245 VDD VSS sg13g2_decap_8
XFILLER_14_651 VDD VSS sg13g2_decap_8
XFILLER_13_161 VDD VSS sg13g2_decap_8
XFILLER_9_154 VDD VSS sg13g2_decap_8
XFILLER_5_371 VDD VSS sg13g2_decap_8
XFILLER_68_356 VDD VSS sg13g2_decap_8
XFILLER_95_175 VDD VSS sg13g2_decap_8
XFILLER_83_315 VDD VSS sg13g2_decap_8
XFILLER_56_518 VDD VSS sg13g2_decap_8
XFILLER_3_84 VDD VSS sg13g2_decap_8
XFILLER_49_581 VDD VSS sg13g2_decap_8
XFILLER_37_721 VDD VSS sg13g2_decap_8
XFILLER_36_231 VDD VSS sg13g2_decap_8
XFILLER_64_595 VDD VSS sg13g2_decap_8
XFILLER_52_735 VDD VSS sg13g2_decap_8
XFILLER_91_392 VDD VSS sg13g2_decap_8
XFILLER_24_448 VDD VSS sg13g2_decap_8
XFILLER_51_245 VDD VSS sg13g2_decap_8
XFILLER_22_49 VDD VSS sg13g2_decap_8
XFILLER_20_665 VDD VSS sg13g2_decap_8
XFILLER_3_308 VDD VSS sg13g2_decap_8
XFILLER_59_301 VDD VSS sg13g2_decap_8
XFILLER_87_665 VDD VSS sg13g2_decap_8
XFILLER_47_518 VDD VSS sg13g2_decap_8
XFILLER_47_35 VDD VSS sg13g2_decap_8
XFILLER_59_378 VDD VSS sg13g2_decap_8
XFILLER_86_175 VDD VSS sg13g2_decap_8
XFILLER_74_337 VDD VSS sg13g2_decap_8
XFILLER_28_721 VDD VSS sg13g2_decap_8
XFILLER_27_231 VDD VSS sg13g2_decap_8
XFILLER_55_595 VDD VSS sg13g2_decap_8
XFILLER_43_735 VDD VSS sg13g2_decap_8
XFILLER_70_554 VDD VSS sg13g2_decap_8
XFILLER_82_392 VDD VSS sg13g2_decap_8
XFILLER_63_56 VDD VSS sg13g2_decap_8
XFILLER_15_448 VDD VSS sg13g2_decap_8
XFILLER_42_245 VDD VSS sg13g2_decap_8
XFILLER_11_665 VDD VSS sg13g2_decap_8
XFILLER_7_658 VDD VSS sg13g2_decap_8
XFILLER_10_175 VDD VSS sg13g2_decap_8
XFILLER_6_168 VDD VSS sg13g2_decap_8
XFILLER_88_42 VDD VSS sg13g2_decap_8
XFILLER_2_385 VDD VSS sg13g2_decap_8
XFILLER_93_602 VDD VSS sg13g2_decap_8
XFILLER_78_665 VDD VSS sg13g2_decap_8
XFILLER_38_518 VDD VSS sg13g2_decap_8
XFILLER_92_112 VDD VSS sg13g2_decap_8
XFILLER_77_175 VDD VSS sg13g2_decap_8
XFILLER_65_315 VDD VSS sg13g2_decap_8
XFILLER_19_7 VDD VSS sg13g2_decap_8
XFILLER_19_721 VDD VSS sg13g2_decap_8
XFILLER_93_679 VDD VSS sg13g2_decap_8
XFILLER_18_231 VDD VSS sg13g2_decap_8
XFILLER_92_189 VDD VSS sg13g2_decap_8
XFILLER_80_329 VDD VSS sg13g2_decap_8
XFILLER_46_595 VDD VSS sg13g2_decap_8
XFILLER_34_735 VDD VSS sg13g2_decap_8
XFILLER_61_532 VDD VSS sg13g2_decap_8
XFILLER_33_245 VDD VSS sg13g2_decap_8
XFILLER_45_0 VDD VSS sg13g2_decap_8
XFILLER_69_643 VDD VSS sg13g2_decap_8
XFILLER_84_602 VDD VSS sg13g2_decap_8
XFILLER_29_518 VDD VSS sg13g2_decap_8
XFILLER_83_112 VDD VSS sg13g2_decap_8
XFILLER_68_175 VDD VSS sg13g2_decap_8
XFILLER_56_315 VDD VSS sg13g2_decap_8
XFILLER_84_679 VDD VSS sg13g2_decap_8
XFILLER_83_189 VDD VSS sg13g2_decap_8
XFILLER_17_49 VDD VSS sg13g2_decap_8
XFILLER_25_735 VDD VSS sg13g2_decap_8
XFILLER_64_392 VDD VSS sg13g2_decap_8
XFILLER_52_532 VDD VSS sg13g2_decap_8
XFILLER_24_245 VDD VSS sg13g2_decap_8
XFILLER_37_595 VDD VSS sg13g2_decap_8
XFILLER_40_749 VDD VSS sg13g2_decap_8
XFILLER_20_462 VDD VSS sg13g2_decap_8
XFILLER_3_105 VDD VSS sg13g2_decap_8
XFILLER_58_56 VDD VSS sg13g2_decap_8
XFILLER_75_613 VDD VSS sg13g2_decap_8
XFILLER_87_462 VDD VSS sg13g2_decap_8
XFILLER_74_112 VDD VSS sg13g2_decap_8
XFILLER_47_315 VDD VSS sg13g2_decap_8
XFILLER_59_175 VDD VSS sg13g2_decap_8
XFILLER_90_616 VDD VSS sg13g2_decap_8
XFILLER_74_189 VDD VSS sg13g2_decap_8
XFILLER_62_329 VDD VSS sg13g2_decap_8
XFILLER_74_77 VDD VSS sg13g2_decap_8
XFILLER_55_392 VDD VSS sg13g2_decap_8
XFILLER_16_735 VDD VSS sg13g2_decap_8
XFILLER_28_595 VDD VSS sg13g2_decap_8
XFILLER_43_532 VDD VSS sg13g2_decap_8
XFILLER_70_362 VDD VSS sg13g2_decap_8
XFILLER_90_21 VDD VSS sg13g2_decap_8
XFILLER_15_245 VDD VSS sg13g2_decap_8
XFILLER_31_749 VDD VSS sg13g2_decap_8
XFILLER_30_259 VDD VSS sg13g2_decap_8
XFILLER_90_98 VDD VSS sg13g2_decap_8
XFILLER_11_462 VDD VSS sg13g2_decap_8
XFILLER_23_70 VDD VSS sg13g2_decap_8
XFILLER_7_455 VDD VSS sg13g2_decap_8
XFILLER_3_672 VDD VSS sg13g2_decap_8
XFILLER_2_182 VDD VSS sg13g2_decap_8
XFILLER_78_462 VDD VSS sg13g2_decap_8
XFILLER_66_646 VDD VSS sg13g2_decap_8
XFILLER_65_112 VDD VSS sg13g2_decap_8
XFILLER_38_315 VDD VSS sg13g2_decap_8
XFILLER_81_616 VDD VSS sg13g2_decap_8
XFILLER_93_476 VDD VSS sg13g2_decap_8
XFILLER_65_189 VDD VSS sg13g2_decap_8
XFILLER_53_329 VDD VSS sg13g2_decap_8
XFILLER_80_126 VDD VSS sg13g2_decap_8
XFILLER_0_63 VDD VSS sg13g2_decap_8
XFILLER_46_392 VDD VSS sg13g2_decap_8
XFILLER_19_595 VDD VSS sg13g2_decap_8
XFILLER_34_532 VDD VSS sg13g2_decap_8
XFILLER_22_749 VDD VSS sg13g2_decap_8
XFILLER_21_259 VDD VSS sg13g2_decap_8
XFILLER_1_609 VDD VSS sg13g2_decap_8
XFILLER_89_749 VDD VSS sg13g2_decap_8
XFILLER_0_119 VDD VSS sg13g2_decap_8
XFILLER_88_259 VDD VSS sg13g2_decap_8
XFILLER_69_462 VDD VSS sg13g2_decap_8
XFILLER_57_602 VDD VSS sg13g2_decap_8
XFILLER_29_315 VDD VSS sg13g2_decap_8
XFILLER_56_112 VDD VSS sg13g2_decap_8
XFILLER_57_679 VDD VSS sg13g2_decap_8
XFILLER_84_476 VDD VSS sg13g2_decap_8
XIO_BOND_outputs\[8\].output_pad output_PAD[8] bondpad_70x70_novias
XFILLER_44_329 VDD VSS sg13g2_decap_8
XFILLER_56_189 VDD VSS sg13g2_decap_8
XFILLER_72_649 VDD VSS sg13g2_decap_8
XFILLER_71_126 VDD VSS sg13g2_decap_8
XFILLER_44_14 VDD VSS sg13g2_decap_8
XFILLER_37_392 VDD VSS sg13g2_decap_8
XFILLER_25_532 VDD VSS sg13g2_decap_8
XFILLER_80_693 VDD VSS sg13g2_decap_8
XFILLER_13_749 VDD VSS sg13g2_decap_8
XFILLER_12_259 VDD VSS sg13g2_decap_8
XFILLER_40_546 VDD VSS sg13g2_decap_8
XFILLER_60_35 VDD VSS sg13g2_decap_8
XFILLER_4_469 VDD VSS sg13g2_decap_8
XFILLER_69_77 VDD VSS sg13g2_decap_8
XFILLER_79_259 VDD VSS sg13g2_decap_8
XFILLER_48_602 VDD VSS sg13g2_decap_8
XFILLER_85_21 VDD VSS sg13g2_decap_8
XFILLER_0_686 VDD VSS sg13g2_decap_8
XFILLER_47_112 VDD VSS sg13g2_decap_8
XFILLER_48_679 VDD VSS sg13g2_decap_8
XFILLER_75_487 VDD VSS sg13g2_decap_8
XFILLER_63_627 VDD VSS sg13g2_decap_8
XFILLER_90_413 VDD VSS sg13g2_decap_8
XFILLER_85_98 VDD VSS sg13g2_decap_8
XFILLER_18_70 VDD VSS sg13g2_decap_8
XFILLER_35_329 VDD VSS sg13g2_decap_8
XFILLER_47_189 VDD VSS sg13g2_decap_8
XFILLER_62_126 VDD VSS sg13g2_decap_8
XFILLER_28_392 VDD VSS sg13g2_decap_8
XFILLER_16_532 VDD VSS sg13g2_decap_8
XFILLER_71_660 VDD VSS sg13g2_decap_8
XFILLER_34_91 VDD VSS sg13g2_decap_8
XFILLER_31_546 VDD VSS sg13g2_decap_8
XFILLER_86_7 VDD VSS sg13g2_decap_8
XFILLER_8_742 VDD VSS sg13g2_decap_8
XFILLER_7_252 VDD VSS sg13g2_decap_8
XFILLER_39_602 VDD VSS sg13g2_decap_8
XFILLER_38_112 VDD VSS sg13g2_decap_8
XFILLER_93_273 VDD VSS sg13g2_decap_8
XFILLER_81_413 VDD VSS sg13g2_decap_8
XFILLER_54_616 VDD VSS sg13g2_decap_8
XFILLER_26_307 VDD VSS sg13g2_decap_8
XFILLER_39_679 VDD VSS sg13g2_decap_8
XFILLER_19_392 VDD VSS sg13g2_decap_8
XFILLER_38_189 VDD VSS sg13g2_decap_8
XFILLER_53_126 VDD VSS sg13g2_decap_8
XFILLER_62_693 VDD VSS sg13g2_decap_8
XFILLER_14_28 VDD VSS sg13g2_decap_8
XFILLER_22_546 VDD VSS sg13g2_decap_8
XFILLER_30_49 VDD VSS sg13g2_decap_8
XFILLER_1_406 VDD VSS sg13g2_decap_8
XFILLER_89_546 VDD VSS sg13g2_decap_8
XFILLER_39_14 VDD VSS sg13g2_decap_8
XFILLER_29_112 VDD VSS sg13g2_decap_8
XFILLER_84_273 VDD VSS sg13g2_decap_8
XFILLER_72_402 VDD VSS sg13g2_decap_8
XFILLER_55_35 VDD VSS sg13g2_decap_8
XFILLER_57_476 VDD VSS sg13g2_decap_8
XFILLER_45_616 VDD VSS sg13g2_decap_8
XFILLER_72_446 VDD VSS sg13g2_decap_8
XFILLER_17_329 VDD VSS sg13g2_decap_8
XFILLER_29_189 VDD VSS sg13g2_decap_8
XFILLER_44_126 VDD VSS sg13g2_decap_8
XFILLER_53_693 VDD VSS sg13g2_decap_8
XFILLER_80_490 VDD VSS sg13g2_decap_8
XFILLER_71_56 VDD VSS sg13g2_decap_8
XFILLER_13_546 VDD VSS sg13g2_decap_8
XFILLER_40_343 VDD VSS sg13g2_decap_8
XFILLER_9_539 VDD VSS sg13g2_decap_8
XFILLER_5_756 VDD VSS sg13g2_fill_1
XFILLER_4_266 VDD VSS sg13g2_decap_8
XFILLER_76_741 VDD VSS sg13g2_decap_8
XFILLER_0_483 VDD VSS sg13g2_decap_8
XFILLER_91_700 VDD VSS sg13g2_decap_8
XFILLER_63_413 VDD VSS sg13g2_decap_8
XFILLER_29_91 VDD VSS sg13g2_decap_8
XFILLER_48_476 VDD VSS sg13g2_decap_8
XFILLER_36_616 VDD VSS sg13g2_decap_8
XFILLER_90_210 VDD VSS sg13g2_decap_8
XFILLER_35_126 VDD VSS sg13g2_decap_8
XFILLER_90_287 VDD VSS sg13g2_decap_8
XFILLER_44_693 VDD VSS sg13g2_decap_8
XFILLER_31_343 VDD VSS sg13g2_decap_8
XFILLER_6_84 VDD VSS sg13g2_decap_8
XFILLER_67_730 VDD VSS sg13g2_decap_8
XFILLER_94_560 VDD VSS sg13g2_decap_8
XFILLER_82_700 VDD VSS sg13g2_decap_8
XFILLER_39_476 VDD VSS sg13g2_decap_8
XFILLER_27_616 VDD VSS sg13g2_decap_8
XFILLER_81_210 VDD VSS sg13g2_decap_8
XFILLER_66_273 VDD VSS sg13g2_decap_8
XFILLER_26_126 VDD VSS sg13g2_decap_8
XFILLER_54_413 VDD VSS sg13g2_decap_8
XFILLER_81_287 VDD VSS sg13g2_decap_8
XFILLER_25_49 VDD VSS sg13g2_decap_8
XFILLER_35_693 VDD VSS sg13g2_decap_8
XFILLER_62_490 VDD VSS sg13g2_decap_8
XFILLER_50_630 VDD VSS sg13g2_decap_8
XFILLER_22_343 VDD VSS sg13g2_decap_8
XFILLER_1_203 VDD VSS sg13g2_decap_8
XFILLER_89_343 VDD VSS sg13g2_decap_8
XFILLER_77_527 VDD VSS sg13g2_decap_8
XFILLER_85_560 VDD VSS sg13g2_decap_8
XFILLER_66_56 VDD VSS sg13g2_decap_8
XFILLER_18_616 VDD VSS sg13g2_decap_8
XFILLER_73_744 VDD VSS sg13g2_decap_8
XFILLER_72_210 VDD VSS sg13g2_decap_8
XFILLER_17_126 VDD VSS sg13g2_decap_8
XFILLER_45_413 VDD VSS sg13g2_decap_8
XFILLER_57_273 VDD VSS sg13g2_decap_8
XFILLER_73_755 VDD VSS sg13g2_fill_2
XFILLER_72_287 VDD VSS sg13g2_decap_8
XFILLER_60_427 VDD VSS sg13g2_decap_8
XFILLER_26_671 VDD VSS sg13g2_decap_8
XFILLER_82_77 VDD VSS sg13g2_decap_8
XFILLER_53_490 VDD VSS sg13g2_decap_8
XFILLER_13_343 VDD VSS sg13g2_decap_8
XFILLER_41_630 VDD VSS sg13g2_decap_8
XFILLER_40_140 VDD VSS sg13g2_decap_8
XFILLER_9_336 VDD VSS sg13g2_decap_8
XFILLER_31_70 VDD VSS sg13g2_decap_8
XFILLER_5_553 VDD VSS sg13g2_decap_8
XFILLER_49_7 VDD VSS sg13g2_decap_8
XFILLER_68_538 VDD VSS sg13g2_decap_8
XFILLER_95_357 VDD VSS sg13g2_decap_8
XFILLER_0_280 VDD VSS sg13g2_decap_8
XFILLER_64_700 VDD VSS sg13g2_decap_8
XFILLER_63_210 VDD VSS sg13g2_decap_8
XFILLER_36_413 VDD VSS sg13g2_decap_8
XFILLER_48_273 VDD VSS sg13g2_decap_8
XFILLER_91_574 VDD VSS sg13g2_decap_8
XFILLER_63_287 VDD VSS sg13g2_decap_8
XFILLER_51_427 VDD VSS sg13g2_decap_8
XFILLER_17_693 VDD VSS sg13g2_decap_8
XFILLER_32_630 VDD VSS sg13g2_decap_8
XFILLER_44_490 VDD VSS sg13g2_decap_8
XFILLER_31_140 VDD VSS sg13g2_decap_8
XFILLER_75_0 VDD VSS sg13g2_decap_8
XFILLER_86_357 VDD VSS sg13g2_decap_8
XFILLER_55_700 VDD VSS sg13g2_decap_8
XFILLER_27_413 VDD VSS sg13g2_decap_8
XFILLER_39_273 VDD VSS sg13g2_decap_8
XFILLER_54_210 VDD VSS sg13g2_decap_8
XFILLER_82_574 VDD VSS sg13g2_decap_8
XFILLER_70_736 VDD VSS sg13g2_decap_8
XFILLER_42_427 VDD VSS sg13g2_decap_8
XFILLER_54_287 VDD VSS sg13g2_decap_8
XFILLER_52_14 VDD VSS sg13g2_decap_8
XFILLER_23_630 VDD VSS sg13g2_decap_8
XFILLER_35_490 VDD VSS sg13g2_decap_8
XFILLER_22_140 VDD VSS sg13g2_decap_8
XFILLER_10_357 VDD VSS sg13g2_decap_8
XFILLER_89_140 VDD VSS sg13g2_decap_8
XFILLER_77_302 VDD VSS sg13g2_decap_8
XFILLER_2_567 VDD VSS sg13g2_decap_8
XFILLER_77_77 VDD VSS sg13g2_decap_8
XFILLER_77_379 VDD VSS sg13g2_decap_8
XFILLER_58_560 VDD VSS sg13g2_decap_8
XFILLER_46_700 VDD VSS sg13g2_decap_8
XFILLER_93_21 VDD VSS sg13g2_decap_8
XFILLER_18_413 VDD VSS sg13g2_decap_8
XFILLER_45_210 VDD VSS sg13g2_decap_8
XFILLER_73_541 VDD VSS sg13g2_decap_8
XFILLER_93_98 VDD VSS sg13g2_decap_8
XFILLER_61_714 VDD VSS sg13g2_decap_8
XFILLER_33_427 VDD VSS sg13g2_decap_8
XFILLER_45_287 VDD VSS sg13g2_decap_8
XFILLER_26_70 VDD VSS sg13g2_decap_8
XFILLER_60_224 VDD VSS sg13g2_decap_8
XFILLER_14_630 VDD VSS sg13g2_decap_8
XFILLER_13_140 VDD VSS sg13g2_decap_8
XFILLER_9_133 VDD VSS sg13g2_decap_8
XFILLER_42_91 VDD VSS sg13g2_decap_8
XIO_BOND_iovss_pads\[0\].iovss_pad IOVSS bondpad_70x70_novias
XFILLER_5_350 VDD VSS sg13g2_decap_8
XFILLER_68_335 VDD VSS sg13g2_decap_8
XFILLER_3_63 VDD VSS sg13g2_decap_8
XFILLER_95_154 VDD VSS sg13g2_decap_8
XFILLER_49_560 VDD VSS sg13g2_decap_8
XFILLER_37_700 VDD VSS sg13g2_decap_8
XFILLER_36_210 VDD VSS sg13g2_decap_8
XFILLER_76_390 VDD VSS sg13g2_decap_8
XFILLER_64_574 VDD VSS sg13g2_decap_8
XFILLER_91_371 VDD VSS sg13g2_decap_8
XFILLER_52_714 VDD VSS sg13g2_decap_8
XFILLER_24_427 VDD VSS sg13g2_decap_8
XFILLER_36_287 VDD VSS sg13g2_decap_8
XFILLER_51_224 VDD VSS sg13g2_decap_8
XFILLER_17_490 VDD VSS sg13g2_decap_8
XFILLER_22_28 VDD VSS sg13g2_decap_8
XFILLER_20_644 VDD VSS sg13g2_decap_8
XFILLER_87_644 VDD VSS sg13g2_decap_8
XFILLER_86_154 VDD VSS sg13g2_decap_8
XFILLER_47_14 VDD VSS sg13g2_decap_8
XFILLER_59_357 VDD VSS sg13g2_decap_8
XFILLER_28_700 VDD VSS sg13g2_decap_8
XFILLER_74_316 VDD VSS sg13g2_decap_8
XFILLER_27_210 VDD VSS sg13g2_decap_8
XFILLER_82_371 VDD VSS sg13g2_decap_8
XFILLER_55_574 VDD VSS sg13g2_decap_8
XFILLER_15_427 VDD VSS sg13g2_decap_8
XFILLER_43_714 VDD VSS sg13g2_decap_8
XFILLER_70_533 VDD VSS sg13g2_decap_8
XFILLER_63_35 VDD VSS sg13g2_decap_8
XFILLER_27_287 VDD VSS sg13g2_decap_8
XFILLER_42_224 VDD VSS sg13g2_decap_8
XFILLER_11_644 VDD VSS sg13g2_decap_8
XFILLER_7_637 VDD VSS sg13g2_decap_8
XFILLER_10_154 VDD VSS sg13g2_decap_8
XFILLER_6_147 VDD VSS sg13g2_decap_8
XFILLER_88_21 VDD VSS sg13g2_decap_8
XFILLER_5_0 VDD VSS sg13g2_decap_8
XFILLER_88_98 VDD VSS sg13g2_decap_8
XFILLER_2_364 VDD VSS sg13g2_decap_8
XFILLER_78_644 VDD VSS sg13g2_decap_8
XFILLER_77_154 VDD VSS sg13g2_decap_8
XFILLER_19_700 VDD VSS sg13g2_decap_8
XFILLER_18_210 VDD VSS sg13g2_decap_8
XFILLER_93_658 VDD VSS sg13g2_decap_8
XFILLER_92_168 VDD VSS sg13g2_decap_8
XFILLER_80_308 VDD VSS sg13g2_decap_8
XFILLER_61_511 VDD VSS sg13g2_decap_8
XFILLER_46_574 VDD VSS sg13g2_decap_8
XFILLER_37_91 VDD VSS sg13g2_decap_8
XFILLER_34_714 VDD VSS sg13g2_decap_8
XFILLER_18_287 VDD VSS sg13g2_decap_8
XFILLER_33_224 VDD VSS sg13g2_decap_8
XFILLER_61_588 VDD VSS sg13g2_decap_8
XFILLER_69_622 VDD VSS sg13g2_decap_8
XFILLER_38_0 VDD VSS sg13g2_decap_8
XFILLER_68_154 VDD VSS sg13g2_decap_8
XFILLER_69_699 VDD VSS sg13g2_decap_8
XFILLER_84_658 VDD VSS sg13g2_decap_8
XFILLER_17_28 VDD VSS sg13g2_decap_8
XFILLER_83_168 VDD VSS sg13g2_decap_8
XFILLER_64_371 VDD VSS sg13g2_decap_8
XFILLER_52_511 VDD VSS sg13g2_decap_8
XFILLER_25_714 VDD VSS sg13g2_decap_8
XFILLER_37_574 VDD VSS sg13g2_decap_8
XFILLER_24_224 VDD VSS sg13g2_decap_8
XFILLER_40_728 VDD VSS sg13g2_decap_8
XFILLER_52_588 VDD VSS sg13g2_decap_8
XFILLER_33_49 VDD VSS sg13g2_decap_8
XFILLER_20_441 VDD VSS sg13g2_decap_8
XFILLER_58_35 VDD VSS sg13g2_decap_8
XFILLER_87_441 VDD VSS sg13g2_decap_8
XFILLER_59_154 VDD VSS sg13g2_decap_8
XFILLER_75_669 VDD VSS sg13g2_decap_8
XFILLER_74_168 VDD VSS sg13g2_decap_8
XFILLER_62_308 VDD VSS sg13g2_decap_8
XFILLER_74_56 VDD VSS sg13g2_decap_8
XFILLER_16_714 VDD VSS sg13g2_decap_8
XFILLER_28_574 VDD VSS sg13g2_decap_8
XFILLER_43_511 VDD VSS sg13g2_decap_8
XFILLER_15_224 VDD VSS sg13g2_decap_8
XFILLER_55_371 VDD VSS sg13g2_decap_8
XFILLER_70_341 VDD VSS sg13g2_decap_8
XFILLER_31_728 VDD VSS sg13g2_decap_8
XFILLER_43_588 VDD VSS sg13g2_decap_8
XFILLER_90_77 VDD VSS sg13g2_decap_8
XFILLER_11_441 VDD VSS sg13g2_decap_8
XFILLER_30_238 VDD VSS sg13g2_decap_8
XFILLER_7_434 VDD VSS sg13g2_decap_8
XFILLER_3_651 VDD VSS sg13g2_decap_8
XFILLER_2_161 VDD VSS sg13g2_decap_8
XFILLER_31_7 VDD VSS sg13g2_decap_8
XFILLER_78_441 VDD VSS sg13g2_decap_8
XFILLER_66_625 VDD VSS sg13g2_decap_8
XFILLER_93_455 VDD VSS sg13g2_decap_8
XFILLER_65_168 VDD VSS sg13g2_decap_8
XFILLER_80_105 VDD VSS sg13g2_decap_8
XFILLER_0_42 VDD VSS sg13g2_decap_8
XFILLER_53_308 VDD VSS sg13g2_decap_8
XFILLER_19_574 VDD VSS sg13g2_decap_8
XFILLER_46_371 VDD VSS sg13g2_decap_8
XFILLER_34_511 VDD VSS sg13g2_decap_8
XFILLER_61_385 VDD VSS sg13g2_decap_8
XFILLER_22_728 VDD VSS sg13g2_decap_8
XFILLER_34_588 VDD VSS sg13g2_decap_8
XFILLER_21_238 VDD VSS sg13g2_decap_8
XFILLER_9_84 VDD VSS sg13g2_decap_8
XFILLER_89_728 VDD VSS sg13g2_decap_8
XFILLER_88_238 VDD VSS sg13g2_decap_8
XFILLER_69_496 VDD VSS sg13g2_decap_8
XFILLER_84_455 VDD VSS sg13g2_decap_8
XFILLER_57_658 VDD VSS sg13g2_decap_8
XFILLER_28_49 VDD VSS sg13g2_decap_8
XFILLER_72_628 VDD VSS sg13g2_decap_8
XFILLER_71_105 VDD VSS sg13g2_decap_8
XFILLER_44_308 VDD VSS sg13g2_decap_8
XFILLER_56_168 VDD VSS sg13g2_decap_8
XFILLER_37_371 VDD VSS sg13g2_decap_8
XFILLER_25_511 VDD VSS sg13g2_decap_8
XFILLER_80_672 VDD VSS sg13g2_decap_8
XFILLER_13_728 VDD VSS sg13g2_decap_8
XFILLER_52_385 VDD VSS sg13g2_decap_8
XFILLER_25_588 VDD VSS sg13g2_decap_8
XFILLER_40_525 VDD VSS sg13g2_decap_8
XFILLER_12_238 VDD VSS sg13g2_decap_8
XFILLER_60_14 VDD VSS sg13g2_decap_8
XFILLER_4_448 VDD VSS sg13g2_decap_8
XFILLER_69_56 VDD VSS sg13g2_decap_8
XFILLER_79_238 VDD VSS sg13g2_decap_8
XFILLER_0_665 VDD VSS sg13g2_decap_8
XFILLER_75_444 VDD VSS sg13g2_decap_8
XFILLER_85_77 VDD VSS sg13g2_decap_8
XFILLER_48_658 VDD VSS sg13g2_decap_8
XFILLER_63_606 VDD VSS sg13g2_decap_8
XFILLER_62_105 VDD VSS sg13g2_decap_8
XFILLER_35_308 VDD VSS sg13g2_decap_8
XFILLER_47_168 VDD VSS sg13g2_decap_8
XFILLER_28_371 VDD VSS sg13g2_decap_8
XFILLER_16_511 VDD VSS sg13g2_decap_8
XFILLER_90_469 VDD VSS sg13g2_decap_8
XFILLER_43_385 VDD VSS sg13g2_decap_8
XFILLER_16_588 VDD VSS sg13g2_decap_8
XFILLER_31_525 VDD VSS sg13g2_decap_8
XFILLER_70_182 VDD VSS sg13g2_decap_8
XFILLER_34_70 VDD VSS sg13g2_decap_8
XFILLER_8_721 VDD VSS sg13g2_decap_8
XFILLER_79_7 VDD VSS sg13g2_decap_8
XFILLER_7_231 VDD VSS sg13g2_decap_8
XFILLER_50_91 VDD VSS sg13g2_decap_8
XFILLER_94_742 VDD VSS sg13g2_decap_8
XFILLER_39_658 VDD VSS sg13g2_decap_8
XFILLER_93_252 VDD VSS sg13g2_decap_8
XFILLER_53_105 VDD VSS sg13g2_decap_8
XFILLER_38_168 VDD VSS sg13g2_decap_8
XFILLER_66_499 VDD VSS sg13g2_decap_8
XFILLER_19_371 VDD VSS sg13g2_decap_8
XFILLER_81_469 VDD VSS sg13g2_decap_8
XFILLER_62_672 VDD VSS sg13g2_decap_8
XFILLER_34_385 VDD VSS sg13g2_decap_8
XFILLER_22_525 VDD VSS sg13g2_decap_8
XFILLER_61_182 VDD VSS sg13g2_decap_8
XFILLER_30_28 VDD VSS sg13g2_decap_8
XFILLER_89_525 VDD VSS sg13g2_decap_8
XFILLER_77_709 VDD VSS sg13g2_decap_8
XFILLER_85_742 VDD VSS sg13g2_decap_8
XFILLER_69_282 VDD VSS sg13g2_decap_8
XFILLER_84_252 VDD VSS sg13g2_decap_8
XFILLER_55_14 VDD VSS sg13g2_decap_8
XFILLER_17_308 VDD VSS sg13g2_decap_8
XFILLER_29_168 VDD VSS sg13g2_decap_8
XFILLER_57_455 VDD VSS sg13g2_decap_8
XFILLER_44_105 VDD VSS sg13g2_decap_8
XFILLER_60_609 VDD VSS sg13g2_decap_8
XFILLER_53_672 VDD VSS sg13g2_decap_8
XFILLER_13_525 VDD VSS sg13g2_decap_8
XFILLER_25_385 VDD VSS sg13g2_decap_8
XFILLER_71_35 VDD VSS sg13g2_decap_8
XFILLER_40_322 VDD VSS sg13g2_decap_8
XFILLER_52_182 VDD VSS sg13g2_decap_8
XFILLER_9_518 VDD VSS sg13g2_decap_8
XFILLER_40_399 VDD VSS sg13g2_decap_8
XFILLER_5_735 VDD VSS sg13g2_decap_8
XFILLER_4_245 VDD VSS sg13g2_decap_8
XFILLER_95_539 VDD VSS sg13g2_decap_8
XFILLER_76_720 VDD VSS sg13g2_decap_8
XFILLER_67_219 VDD VSS sg13g2_decap_8
XFILLER_0_462 VDD VSS sg13g2_decap_8
XFILLER_29_70 VDD VSS sg13g2_decap_8
XFILLER_48_455 VDD VSS sg13g2_decap_8
XFILLER_91_756 VDD VSS sg13g2_fill_1
XFILLER_35_105 VDD VSS sg13g2_decap_8
XFILLER_51_609 VDD VSS sg13g2_decap_8
XFILLER_90_266 VDD VSS sg13g2_decap_8
XFILLER_45_91 VDD VSS sg13g2_decap_8
XFILLER_16_385 VDD VSS sg13g2_decap_8
XFILLER_50_119 VDD VSS sg13g2_decap_8
XFILLER_44_672 VDD VSS sg13g2_decap_8
XFILLER_31_322 VDD VSS sg13g2_decap_8
XFILLER_43_182 VDD VSS sg13g2_decap_8
XFILLER_31_399 VDD VSS sg13g2_decap_8
XFILLER_8_595 VDD VSS sg13g2_decap_8
XFILLER_6_63 VDD VSS sg13g2_decap_8
XFILLER_86_539 VDD VSS sg13g2_decap_8
XFILLER_20_0 VDD VSS sg13g2_decap_8
XFILLER_66_252 VDD VSS sg13g2_decap_8
XFILLER_39_455 VDD VSS sg13g2_decap_8
XFILLER_26_105 VDD VSS sg13g2_decap_8
XFILLER_82_756 VDD VSS sg13g2_fill_1
XFILLER_54_469 VDD VSS sg13g2_decap_8
XFILLER_42_609 VDD VSS sg13g2_decap_8
XFILLER_81_266 VDD VSS sg13g2_decap_8
XFILLER_25_28 VDD VSS sg13g2_decap_8
XFILLER_41_119 VDD VSS sg13g2_decap_8
XFILLER_35_672 VDD VSS sg13g2_decap_8
XFILLER_22_322 VDD VSS sg13g2_decap_8
XFILLER_34_182 VDD VSS sg13g2_decap_8
XFILLER_50_686 VDD VSS sg13g2_decap_8
XFILLER_10_539 VDD VSS sg13g2_decap_8
XFILLER_22_399 VDD VSS sg13g2_decap_8
XFILLER_41_49 VDD VSS sg13g2_decap_8
XIO_BOND_iovdd_pads\[0\].iovdd_pad IOVDD bondpad_70x70_novias
XFILLER_89_322 VDD VSS sg13g2_decap_8
XFILLER_2_749 VDD VSS sg13g2_decap_8
XFILLER_9_7 VDD VSS sg13g2_decap_8
XFILLER_1_259 VDD VSS sg13g2_decap_8
XFILLER_77_506 VDD VSS sg13g2_decap_8
XFILLER_89_399 VDD VSS sg13g2_decap_8
XFILLER_66_35 VDD VSS sg13g2_decap_8
XFILLER_58_742 VDD VSS sg13g2_decap_8
XFILLER_57_252 VDD VSS sg13g2_decap_8
XFILLER_73_723 VDD VSS sg13g2_decap_8
XFILLER_17_105 VDD VSS sg13g2_decap_8
XFILLER_45_469 VDD VSS sg13g2_decap_8
XFILLER_26_650 VDD VSS sg13g2_decap_8
XFILLER_33_609 VDD VSS sg13g2_decap_8
XFILLER_72_277 VDD VSS sg13g2_fill_2
XFILLER_82_56 VDD VSS sg13g2_decap_8
XFILLER_32_119 VDD VSS sg13g2_decap_8
XFILLER_60_406 VDD VSS sg13g2_decap_8
XFILLER_13_322 VDD VSS sg13g2_decap_8
XFILLER_25_182 VDD VSS sg13g2_decap_8
XFILLER_9_315 VDD VSS sg13g2_decap_8
XFILLER_41_686 VDD VSS sg13g2_decap_8
XFILLER_13_399 VDD VSS sg13g2_decap_8
XFILLER_40_196 VDD VSS sg13g2_decap_8
XFILLER_5_532 VDD VSS sg13g2_decap_8
X_80__4 VDD VSS _80__4/L_HI sg13g2_tiehi
XFILLER_68_517 VDD VSS sg13g2_decap_8
XFILLER_95_336 VDD VSS sg13g2_decap_8
XFILLER_49_742 VDD VSS sg13g2_decap_8
XFILLER_48_252 VDD VSS sg13g2_decap_8
XFILLER_76_594 VDD VSS sg13g2_decap_8
XFILLER_91_553 VDD VSS sg13g2_decap_8
XFILLER_64_756 VDD VSS sg13g2_fill_1
XFILLER_36_469 VDD VSS sg13g2_decap_8
XFILLER_24_609 VDD VSS sg13g2_decap_8
XFILLER_63_266 VDD VSS sg13g2_decap_8
XFILLER_23_119 VDD VSS sg13g2_decap_8
XFILLER_51_406 VDD VSS sg13g2_decap_8
XFILLER_17_672 VDD VSS sg13g2_decap_8
XFILLER_16_182 VDD VSS sg13g2_decap_8
XFILLER_32_686 VDD VSS sg13g2_decap_8
XFILLER_31_196 VDD VSS sg13g2_decap_8
XFILLER_68_0 VDD VSS sg13g2_decap_8
XFILLER_8_392 VDD VSS sg13g2_decap_8
XFILLER_86_336 VDD VSS sg13g2_decap_8
XFILLER_59_539 VDD VSS sg13g2_decap_8
XFILLER_39_252 VDD VSS sg13g2_decap_8
XFILLER_67_583 VDD VSS sg13g2_decap_8
XFILLER_82_553 VDD VSS sg13g2_decap_8
XFILLER_55_756 VDD VSS sg13g2_fill_1
XFILLER_36_49 VDD VSS sg13g2_decap_8
XFILLER_27_469 VDD VSS sg13g2_decap_8
XFILLER_15_609 VDD VSS sg13g2_decap_8
XFILLER_70_715 VDD VSS sg13g2_decap_8
XFILLER_14_119 VDD VSS sg13g2_decap_8
XFILLER_42_406 VDD VSS sg13g2_decap_8
XFILLER_54_266 VDD VSS sg13g2_decap_8
XFILLER_50_483 VDD VSS sg13g2_decap_8
XFILLER_23_686 VDD VSS sg13g2_decap_8
XFILLER_10_336 VDD VSS sg13g2_decap_8
XFILLER_22_196 VDD VSS sg13g2_decap_8
XFILLER_6_329 VDD VSS sg13g2_decap_8
XFILLER_2_546 VDD VSS sg13g2_decap_8
XFILLER_89_196 VDD VSS sg13g2_decap_8
XFILLER_77_56 VDD VSS sg13g2_decap_8
XFILLER_77_358 VDD VSS sg13g2_decap_8
XFILLER_73_520 VDD VSS sg13g2_decap_8
XFILLER_46_756 VDD VSS sg13g2_fill_1
XFILLER_18_469 VDD VSS sg13g2_decap_8
XFILLER_93_77 VDD VSS sg13g2_decap_8
XFILLER_33_406 VDD VSS sg13g2_decap_8
XFILLER_45_266 VDD VSS sg13g2_decap_8
XFILLER_60_203 VDD VSS sg13g2_decap_8
XFILLER_73_597 VDD VSS sg13g2_decap_8
XFILLER_9_112 VDD VSS sg13g2_decap_8
XFILLER_14_686 VDD VSS sg13g2_decap_8
XFILLER_41_483 VDD VSS sg13g2_decap_8
XFILLER_13_196 VDD VSS sg13g2_decap_8
XFILLER_42_70 VDD VSS sg13g2_decap_8
XFILLER_9_189 VDD VSS sg13g2_decap_8
XFILLER_61_7 VDD VSS sg13g2_decap_8
XFILLER_68_314 VDD VSS sg13g2_decap_8
XFILLER_3_42 VDD VSS sg13g2_decap_8
XFILLER_95_133 VDD VSS sg13g2_decap_8
XFILLER_64_553 VDD VSS sg13g2_decap_8
XFILLER_37_756 VDD VSS sg13g2_fill_1
XFILLER_91_350 VDD VSS sg13g2_decap_8
XFILLER_24_406 VDD VSS sg13g2_decap_8
XFILLER_36_266 VDD VSS sg13g2_decap_8
XFILLER_51_203 VDD VSS sg13g2_decap_8
XFILLER_20_623 VDD VSS sg13g2_decap_8
XFILLER_32_483 VDD VSS sg13g2_decap_8
Xiovss_pads\[0\].iovss_pad IOVDD IOVSS VDD VSS sg13g2_IOPadIOVss
XFILLER_87_623 VDD VSS sg13g2_decap_8
XFILLER_59_336 VDD VSS sg13g2_decap_8
XFILLER_86_133 VDD VSS sg13g2_decap_8
XFILLER_67_380 VDD VSS sg13g2_decap_8
XFILLER_55_553 VDD VSS sg13g2_decap_8
XFILLER_28_756 VDD VSS sg13g2_fill_1
XFILLER_70_512 VDD VSS sg13g2_decap_8
XFILLER_82_350 VDD VSS sg13g2_decap_8
XFILLER_63_14 VDD VSS sg13g2_decap_8
XFILLER_15_406 VDD VSS sg13g2_decap_8
XFILLER_27_266 VDD VSS sg13g2_decap_8
XFILLER_42_203 VDD VSS sg13g2_decap_8
XFILLER_70_589 VDD VSS sg13g2_decap_8
XFILLER_11_623 VDD VSS sg13g2_decap_8
XFILLER_23_483 VDD VSS sg13g2_decap_8
XFILLER_7_616 VDD VSS sg13g2_decap_8
XFILLER_10_133 VDD VSS sg13g2_decap_8
XFILLER_50_280 VDD VSS sg13g2_decap_8
XFILLER_6_126 VDD VSS sg13g2_decap_8
XFILLER_12_84 VDD VSS sg13g2_decap_8
XFILLER_88_77 VDD VSS sg13g2_decap_8
XFILLER_2_343 VDD VSS sg13g2_decap_8
XFILLER_78_623 VDD VSS sg13g2_decap_8
XFILLER_77_133 VDD VSS sg13g2_decap_8
XFILLER_93_637 VDD VSS sg13g2_decap_8
XFILLER_92_147 VDD VSS sg13g2_decap_8
XFILLER_19_756 VDD VSS sg13g2_fill_1
XFILLER_46_553 VDD VSS sg13g2_decap_8
XFILLER_37_70 VDD VSS sg13g2_decap_8
XFILLER_18_266 VDD VSS sg13g2_decap_8
XFILLER_33_203 VDD VSS sg13g2_decap_8
XFILLER_73_394 VDD VSS sg13g2_decap_8
XFILLER_61_567 VDD VSS sg13g2_decap_8
XFILLER_14_483 VDD VSS sg13g2_decap_8
XFILLER_53_91 VDD VSS sg13g2_decap_8
XFILLER_41_280 VDD VSS sg13g2_decap_8
XFILLER_6_693 VDD VSS sg13g2_decap_8
XFILLER_69_601 VDD VSS sg13g2_decap_8
XFILLER_69_678 VDD VSS sg13g2_decap_8
XFILLER_68_133 VDD VSS sg13g2_decap_8
XFILLER_84_637 VDD VSS sg13g2_decap_8
Xclkbuf_0_clk_PAD2CORE clkbuf_0_clk_PAD2CORE/X clk_pad/p2c VDD VSS sg13g2_buf_16
XFILLER_83_147 VDD VSS sg13g2_decap_8
X_69_ _69_/Y _75_/A _69_/B VDD VSS sg13g2_nand2_1
XFILLER_64_350 VDD VSS sg13g2_decap_8
XFILLER_37_553 VDD VSS sg13g2_decap_8
XFILLER_24_203 VDD VSS sg13g2_decap_8
XFILLER_52_567 VDD VSS sg13g2_decap_8
XFILLER_40_707 VDD VSS sg13g2_decap_8
XFILLER_33_28 VDD VSS sg13g2_decap_8
XFILLER_20_420 VDD VSS sg13g2_decap_8
XFILLER_32_280 VDD VSS sg13g2_decap_8
XFILLER_20_497 VDD VSS sg13g2_decap_8
XFILLER_87_420 VDD VSS sg13g2_decap_8
XFILLER_58_14 VDD VSS sg13g2_decap_8
XFILLER_59_133 VDD VSS sg13g2_decap_8
XFILLER_87_497 VDD VSS sg13g2_decap_8
XFILLER_75_648 VDD VSS sg13g2_decap_8
XFILLER_74_147 VDD VSS sg13g2_decap_8
XFILLER_74_35 VDD VSS sg13g2_decap_8
XFILLER_55_350 VDD VSS sg13g2_decap_8
XFILLER_28_553 VDD VSS sg13g2_decap_8
XFILLER_70_320 VDD VSS sg13g2_decap_8
XFILLER_15_203 VDD VSS sg13g2_decap_8
XFILLER_31_707 VDD VSS sg13g2_decap_8
XFILLER_43_567 VDD VSS sg13g2_decap_8
XFILLER_70_397 VDD VSS sg13g2_decap_8
XFILLER_30_217 VDD VSS sg13g2_decap_8
XFILLER_90_56 VDD VSS sg13g2_decap_8
XFILLER_11_420 VDD VSS sg13g2_decap_8
XFILLER_23_280 VDD VSS sg13g2_decap_8
XFILLER_7_413 VDD VSS sg13g2_decap_8
XFILLER_11_497 VDD VSS sg13g2_decap_8
XFILLER_3_630 VDD VSS sg13g2_decap_8
XFILLER_2_140 VDD VSS sg13g2_decap_8
XFILLER_78_420 VDD VSS sg13g2_decap_8
XFILLER_66_604 VDD VSS sg13g2_decap_8
XFILLER_24_7 VDD VSS sg13g2_decap_8
XFILLER_78_497 VDD VSS sg13g2_decap_8
XFILLER_93_434 VDD VSS sg13g2_decap_8
XFILLER_65_147 VDD VSS sg13g2_decap_8
XFILLER_48_91 VDD VSS sg13g2_decap_8
XFILLER_0_21 VDD VSS sg13g2_decap_8
XFILLER_46_350 VDD VSS sg13g2_decap_8
XFILLER_19_553 VDD VSS sg13g2_decap_8
XFILLER_0_98 VDD VSS sg13g2_decap_8
XFILLER_22_707 VDD VSS sg13g2_decap_8
XFILLER_34_567 VDD VSS sg13g2_decap_8
XFILLER_21_217 VDD VSS sg13g2_decap_8
XFILLER_61_364 VDD VSS sg13g2_decap_8
XFILLER_9_63 VDD VSS sg13g2_decap_8
XFILLER_14_280 VDD VSS sg13g2_decap_8
XFILLER_6_490 VDD VSS sg13g2_decap_8
XFILLER_50_0 VDD VSS sg13g2_decap_8
XFILLER_89_707 VDD VSS sg13g2_decap_8
XFILLER_88_217 VDD VSS sg13g2_decap_8
XFILLER_57_637 VDD VSS sg13g2_decap_8
XFILLER_28_28 VDD VSS sg13g2_decap_8
XFILLER_84_434 VDD VSS sg13g2_decap_8
XFILLER_56_147 VDD VSS sg13g2_decap_8
XFILLER_72_607 VDD VSS sg13g2_decap_8
XFILLER_37_350 VDD VSS sg13g2_decap_8
XFILLER_80_651 VDD VSS sg13g2_decap_8
XFILLER_13_707 VDD VSS sg13g2_decap_8
XFILLER_44_49 VDD VSS sg13g2_decap_8
XFILLER_25_567 VDD VSS sg13g2_decap_8
XFILLER_12_217 VDD VSS sg13g2_decap_8
XFILLER_52_364 VDD VSS sg13g2_decap_8
XFILLER_40_504 VDD VSS sg13g2_decap_8
XFILLER_20_294 VDD VSS sg13g2_decap_8
XFILLER_4_427 VDD VSS sg13g2_decap_8
XFILLER_69_35 VDD VSS sg13g2_decap_8
XFILLER_79_217 VDD VSS sg13g2_decap_8
XFILLER_0_644 VDD VSS sg13g2_decap_8
XFILLER_87_294 VDD VSS sg13g2_decap_8
XFILLER_75_423 VDD VSS sg13g2_decap_8
XFILLER_85_56 VDD VSS sg13g2_decap_8
XFILLER_48_637 VDD VSS sg13g2_decap_8
XFILLER_28_350 VDD VSS sg13g2_decap_8
XFILLER_47_147 VDD VSS sg13g2_decap_8
XFILLER_90_448 VDD VSS sg13g2_decap_8
XFILLER_16_567 VDD VSS sg13g2_decap_8
XFILLER_71_695 VDD VSS sg13g2_decap_8
XFILLER_70_161 VDD VSS sg13g2_decap_8
XFILLER_43_364 VDD VSS sg13g2_decap_8
XFILLER_31_504 VDD VSS sg13g2_decap_8
XFILLER_8_700 VDD VSS sg13g2_decap_8
XFILLER_7_210 VDD VSS sg13g2_decap_8
XFILLER_11_294 VDD VSS sg13g2_decap_8
XFILLER_7_287 VDD VSS sg13g2_decap_8
XFILLER_50_70 VDD VSS sg13g2_decap_8
XFILLER_94_721 VDD VSS sg13g2_decap_8
XFILLER_93_231 VDD VSS sg13g2_decap_8
XFILLER_78_294 VDD VSS sg13g2_decap_8
XFILLER_66_434 VDD VSS sg13g2_decap_8
XFILLER_39_637 VDD VSS sg13g2_decap_8
XFILLER_66_478 VDD VSS sg13g2_decap_8
XFILLER_19_350 VDD VSS sg13g2_decap_8
XFILLER_38_147 VDD VSS sg13g2_decap_8
XFILLER_81_448 VDD VSS sg13g2_decap_8
XFILLER_62_651 VDD VSS sg13g2_decap_8
XFILLER_34_364 VDD VSS sg13g2_decap_8
XFILLER_61_161 VDD VSS sg13g2_decap_8
XFILLER_22_504 VDD VSS sg13g2_decap_8
XFILLER_30_581 VDD VSS sg13g2_decap_8
XFILLER_89_504 VDD VSS sg13g2_decap_8
XFILLER_85_721 VDD VSS sg13g2_decap_8
XFILLER_69_261 VDD VSS sg13g2_decap_8
XFILLER_39_49 VDD VSS sg13g2_decap_8
XFILLER_57_434 VDD VSS sg13g2_decap_8
XFILLER_84_231 VDD VSS sg13g2_decap_8
XFILLER_29_147 VDD VSS sg13g2_decap_8
XFILLER_53_651 VDD VSS sg13g2_decap_8
XFILLER_13_504 VDD VSS sg13g2_decap_8
XFILLER_25_364 VDD VSS sg13g2_decap_8
XFILLER_40_301 VDD VSS sg13g2_decap_8
XFILLER_52_161 VDD VSS sg13g2_decap_8
XFILLER_71_14 VDD VSS sg13g2_decap_8
XFILLER_40_378 VDD VSS sg13g2_decap_8
XFILLER_21_581 VDD VSS sg13g2_decap_8
XFILLER_5_714 VDD VSS sg13g2_decap_8
XFILLER_4_224 VDD VSS sg13g2_decap_8
XFILLER_20_84 VDD VSS sg13g2_decap_8
XFILLER_95_518 VDD VSS sg13g2_decap_8
XFILLER_0_441 VDD VSS sg13g2_decap_8
XFILLER_88_581 VDD VSS sg13g2_decap_8
XFILLER_48_434 VDD VSS sg13g2_decap_8
XFILLER_75_264 VDD VSS sg13g2_decap_8
XFILLER_91_735 VDD VSS sg13g2_decap_8
XFILLER_90_245 VDD VSS sg13g2_decap_8
XFILLER_63_448 VDD VSS sg13g2_decap_4
XFILLER_44_651 VDD VSS sg13g2_decap_8
XFILLER_45_70 VDD VSS sg13g2_decap_8
XFILLER_16_364 VDD VSS sg13g2_decap_8
XFILLER_31_301 VDD VSS sg13g2_decap_8
XFILLER_43_161 VDD VSS sg13g2_decap_8
XFILLER_71_492 VDD VSS sg13g2_decap_8
XFILLER_91_7 VDD VSS sg13g2_decap_8
XFILLER_31_378 VDD VSS sg13g2_decap_8
XFILLER_12_581 VDD VSS sg13g2_decap_8
XFILLER_8_574 VDD VSS sg13g2_decap_8
XFILLER_61_91 VDD VSS sg13g2_decap_8
XFILLER_6_42 VDD VSS sg13g2_decap_8
XFILLER_86_518 VDD VSS sg13g2_decap_8
XFILLER_79_581 VDD VSS sg13g2_decap_8
XFILLER_39_434 VDD VSS sg13g2_decap_8
XFILLER_66_231 VDD VSS sg13g2_decap_8
XFILLER_13_0 VDD VSS sg13g2_decap_8
XFILLER_94_595 VDD VSS sg13g2_decap_8
XFILLER_82_735 VDD VSS sg13g2_decap_8
XFILLER_81_245 VDD VSS sg13g2_decap_8
XFILLER_54_448 VDD VSS sg13g2_decap_8
XFILLER_35_651 VDD VSS sg13g2_decap_8
XFILLER_22_301 VDD VSS sg13g2_decap_8
XFILLER_34_161 VDD VSS sg13g2_decap_8
XFILLER_50_665 VDD VSS sg13g2_decap_8
XFILLER_10_518 VDD VSS sg13g2_decap_8
XFILLER_41_28 VDD VSS sg13g2_decap_8
XFILLER_22_378 VDD VSS sg13g2_decap_8
XFILLER_89_301 VDD VSS sg13g2_decap_8
XFILLER_2_728 VDD VSS sg13g2_decap_8
XFILLER_1_238 VDD VSS sg13g2_decap_8
XFILLER_89_378 VDD VSS sg13g2_decap_8
XFILLER_66_14 VDD VSS sg13g2_decap_8
XFILLER_58_721 VDD VSS sg13g2_decap_8
XFILLER_73_702 VDD VSS sg13g2_decap_8
XFILLER_57_231 VDD VSS sg13g2_decap_8
XFILLER_85_595 VDD VSS sg13g2_decap_8
XFILLER_45_448 VDD VSS sg13g2_decap_8
XFILLER_72_256 VDD VSS sg13g2_decap_8
XFILLER_82_35 VDD VSS sg13g2_decap_8
XFILLER_13_301 VDD VSS sg13g2_decap_8
XFILLER_25_161 VDD VSS sg13g2_decap_8
XFILLER_15_84 VDD VSS sg13g2_decap_8
XFILLER_41_665 VDD VSS sg13g2_decap_8
XFILLER_13_378 VDD VSS sg13g2_decap_8
XFILLER_40_175 VDD VSS sg13g2_decap_8
XFILLER_5_511 VDD VSS sg13g2_decap_8
Xiovdd_pads\[0\].iovdd_pad IOVDD IOVSS VDD VSS sg13g2_IOPadIOVdd
XFILLER_5_588 VDD VSS sg13g2_decap_8
XFILLER_95_315 VDD VSS sg13g2_decap_8
XFILLER_49_721 VDD VSS sg13g2_decap_8
XFILLER_48_231 VDD VSS sg13g2_decap_8
XFILLER_76_573 VDD VSS sg13g2_decap_8
XFILLER_64_735 VDD VSS sg13g2_decap_8
XFILLER_91_532 VDD VSS sg13g2_decap_8
XFILLER_63_245 VDD VSS sg13g2_decap_8
XFILLER_56_91 VDD VSS sg13g2_decap_8
XFILLER_36_448 VDD VSS sg13g2_decap_8
XFILLER_17_651 VDD VSS sg13g2_decap_8
XFILLER_16_161 VDD VSS sg13g2_decap_8
XFILLER_32_665 VDD VSS sg13g2_decap_8
XFILLER_31_175 VDD VSS sg13g2_decap_8
XFILLER_8_371 VDD VSS sg13g2_decap_8
XFILLER_59_518 VDD VSS sg13g2_decap_8
XFILLER_86_315 VDD VSS sg13g2_decap_8
XFILLER_67_562 VDD VSS sg13g2_decap_8
XFILLER_39_231 VDD VSS sg13g2_decap_8
XFILLER_55_735 VDD VSS sg13g2_decap_8
XFILLER_36_28 VDD VSS sg13g2_decap_8
XFILLER_82_532 VDD VSS sg13g2_decap_8
XFILLER_94_392 VDD VSS sg13g2_decap_8
XFILLER_27_448 VDD VSS sg13g2_decap_8
XFILLER_54_245 VDD VSS sg13g2_decap_8
XFILLER_23_665 VDD VSS sg13g2_decap_8
XFILLER_10_315 VDD VSS sg13g2_decap_8
XFILLER_52_49 VDD VSS sg13g2_decap_8
XFILLER_22_175 VDD VSS sg13g2_decap_8
XFILLER_50_462 VDD VSS sg13g2_decap_8
XFILLER_6_308 VDD VSS sg13g2_decap_8
XFILLER_2_525 VDD VSS sg13g2_decap_8
XFILLER_77_35 VDD VSS sg13g2_decap_8
XFILLER_89_175 VDD VSS sg13g2_decap_8
XFILLER_77_337 VDD VSS sg13g2_decap_8
XFILLER_92_329 VDD VSS sg13g2_decap_8
XFILLER_58_595 VDD VSS sg13g2_decap_8
XFILLER_46_735 VDD VSS sg13g2_decap_8
XFILLER_85_392 VDD VSS sg13g2_decap_8
XFILLER_93_56 VDD VSS sg13g2_decap_8
XFILLER_18_448 VDD VSS sg13g2_decap_8
XFILLER_45_245 VDD VSS sg13g2_decap_8
XFILLER_73_576 VDD VSS sg13g2_decap_8
XFILLER_61_749 VDD VSS sg13g2_decap_8
XFILLER_60_259 VDD VSS sg13g2_decap_8
XFILLER_14_665 VDD VSS sg13g2_decap_8
XFILLER_13_175 VDD VSS sg13g2_decap_8
XFILLER_41_462 VDD VSS sg13g2_decap_8
XFILLER_9_168 VDD VSS sg13g2_decap_8
XFILLER_54_7 VDD VSS sg13g2_decap_8
XFILLER_5_385 VDD VSS sg13g2_decap_8
XFILLER_3_21 VDD VSS sg13g2_decap_8
Xvdd_pads\[0\].vdd_pad IOVDD IOVSS VDD VSS sg13g2_IOPadVdd
XFILLER_95_112 VDD VSS sg13g2_decap_8
XFILLER_3_98 VDD VSS sg13g2_decap_8
XFILLER_95_189 VDD VSS sg13g2_decap_8
XFILLER_83_329 VDD VSS sg13g2_decap_8
XFILLER_64_532 VDD VSS sg13g2_decap_8
XFILLER_49_595 VDD VSS sg13g2_decap_8
XFILLER_37_735 VDD VSS sg13g2_decap_8
XFILLER_36_245 VDD VSS sg13g2_decap_8
XFILLER_52_749 VDD VSS sg13g2_decap_8
XFILLER_51_259 VDD VSS sg13g2_decap_8
XFILLER_32_462 VDD VSS sg13g2_decap_8
XFILLER_20_602 VDD VSS sg13g2_decap_8
XFILLER_80_0 VDD VSS sg13g2_decap_8
XFILLER_20_679 VDD VSS sg13g2_decap_8
XFILLER_87_602 VDD VSS sg13g2_decap_8
XFILLER_86_112 VDD VSS sg13g2_decap_8
XFILLER_59_315 VDD VSS sg13g2_decap_8
XFILLER_87_679 VDD VSS sg13g2_decap_8
XFILLER_86_189 VDD VSS sg13g2_decap_8
XFILLER_47_49 VDD VSS sg13g2_decap_8
XFILLER_55_532 VDD VSS sg13g2_decap_8
XFILLER_28_735 VDD VSS sg13g2_decap_8
XFILLER_27_245 VDD VSS sg13g2_decap_8
XFILLER_43_749 VDD VSS sg13g2_decap_8
XFILLER_70_568 VDD VSS sg13g2_decap_8
XFILLER_42_259 VDD VSS sg13g2_decap_8
XFILLER_11_602 VDD VSS sg13g2_decap_8
XFILLER_23_462 VDD VSS sg13g2_decap_8
XFILLER_10_112 VDD VSS sg13g2_decap_8
XFILLER_11_679 VDD VSS sg13g2_decap_8
XFILLER_6_105 VDD VSS sg13g2_decap_8
XFILLER_10_189 VDD VSS sg13g2_decap_8
XFILLER_12_63 VDD VSS sg13g2_decap_8
XFILLER_2_322 VDD VSS sg13g2_decap_8
XFILLER_78_602 VDD VSS sg13g2_decap_8
XFILLER_88_56 VDD VSS sg13g2_decap_8
XFILLER_77_112 VDD VSS sg13g2_decap_8
XFILLER_2_399 VDD VSS sg13g2_decap_8
XFILLER_78_679 VDD VSS sg13g2_decap_8
XFILLER_93_616 VDD VSS sg13g2_decap_8
XFILLER_77_189 VDD VSS sg13g2_decap_8
XFILLER_65_329 VDD VSS sg13g2_decap_8
XFILLER_92_126 VDD VSS sg13g2_decap_8
XFILLER_46_532 VDD VSS sg13g2_decap_8
XFILLER_58_392 VDD VSS sg13g2_decap_8
XFILLER_19_735 VDD VSS sg13g2_decap_8
XFILLER_18_245 VDD VSS sg13g2_decap_8
XFILLER_34_749 VDD VSS sg13g2_decap_8
XFILLER_61_546 VDD VSS sg13g2_decap_8
XFILLER_33_259 VDD VSS sg13g2_decap_8
XFILLER_53_70 VDD VSS sg13g2_decap_8
XFILLER_14_462 VDD VSS sg13g2_decap_8
XFILLER_6_672 VDD VSS sg13g2_decap_8
XFILLER_5_182 VDD VSS sg13g2_decap_8
XFILLER_68_112 VDD VSS sg13g2_decap_8
XFILLER_69_657 VDD VSS sg13g2_decap_8
XFILLER_84_616 VDD VSS sg13g2_decap_8
XFILLER_68_189 VDD VSS sg13g2_decap_8
XFILLER_56_329 VDD VSS sg13g2_decap_8
XFILLER_83_126 VDD VSS sg13g2_decap_8
XFILLER_49_392 VDD VSS sg13g2_decap_8
XFILLER_37_532 VDD VSS sg13g2_decap_8
X_68_ _80_/Q _79_/Q _81_/Q _69_/B VDD VSS _68_/D sg13g2_nand4_1
XFILLER_92_693 VDD VSS sg13g2_decap_8
XFILLER_25_749 VDD VSS sg13g2_decap_8
XFILLER_52_546 VDD VSS sg13g2_decap_8
XFILLER_24_259 VDD VSS sg13g2_decap_8
XFILLER_20_476 VDD VSS sg13g2_decap_8
XFILLER_4_609 VDD VSS sg13g2_decap_8
XFILLER_3_119 VDD VSS sg13g2_decap_8
XFILLER_59_112 VDD VSS sg13g2_decap_8
XFILLER_75_627 VDD VSS sg13g2_decap_8
XFILLER_87_476 VDD VSS sg13g2_decap_8
XFILLER_47_329 VDD VSS sg13g2_decap_8
XFILLER_74_126 VDD VSS sg13g2_decap_8
XFILLER_74_14 VDD VSS sg13g2_decap_8
XFILLER_59_189 VDD VSS sg13g2_decap_8
XFILLER_28_532 VDD VSS sg13g2_decap_8
XFILLER_83_693 VDD VSS sg13g2_decap_8
XFILLER_16_749 VDD VSS sg13g2_decap_4
XFILLER_15_259 VDD VSS sg13g2_decap_8
XFILLER_43_546 VDD VSS sg13g2_decap_8
XFILLER_70_376 VDD VSS sg13g2_decap_8
XFILLER_90_35 VDD VSS sg13g2_decap_8
XFILLER_11_476 VDD VSS sg13g2_decap_8
XFILLER_23_84 VDD VSS sg13g2_decap_8
XFILLER_7_469 VDD VSS sg13g2_decap_8
XFILLER_3_686 VDD VSS sg13g2_decap_8
XFILLER_2_196 VDD VSS sg13g2_decap_8
XFILLER_93_413 VDD VSS sg13g2_decap_8
XFILLER_78_476 VDD VSS sg13g2_decap_8
XFILLER_48_70 VDD VSS sg13g2_decap_8
Xoutputs\[1\].output_pad _77_/Q IOVDD IOVSS output_PAD[1] VDD VSS sg13g2_IOPadOut30mA
XFILLER_65_126 VDD VSS sg13g2_decap_8
XFILLER_17_7 VDD VSS sg13g2_decap_8
XFILLER_38_329 VDD VSS sg13g2_decap_8
XFILLER_19_532 VDD VSS sg13g2_decap_8
XFILLER_74_693 VDD VSS sg13g2_decap_8
XFILLER_0_77 VDD VSS sg13g2_decap_8
XFILLER_64_91 VDD VSS sg13g2_decap_8
XFILLER_61_343 VDD VSS sg13g2_decap_8
XFILLER_34_546 VDD VSS sg13g2_decap_8
XFILLER_9_42 VDD VSS sg13g2_decap_8
XFILLER_43_0 VDD VSS sg13g2_decap_8
XFILLER_84_413 VDD VSS sg13g2_decap_8
XFILLER_57_616 VDD VSS sg13g2_decap_8
XFILLER_29_329 VDD VSS sg13g2_decap_8
XFILLER_56_126 VDD VSS sg13g2_decap_8
XFILLER_65_682 VDD VSS sg13g2_decap_8
XFILLER_92_490 VDD VSS sg13g2_decap_8
XFILLER_80_630 VDD VSS sg13g2_decap_8
XFILLER_44_28 VDD VSS sg13g2_decap_8
XFILLER_52_343 VDD VSS sg13g2_decap_8
XFILLER_25_546 VDD VSS sg13g2_decap_8
XFILLER_60_49 VDD VSS sg13g2_decap_8
XFILLER_20_273 VDD VSS sg13g2_decap_8
XFILLER_4_406 VDD VSS sg13g2_decap_8
XFILLER_69_14 VDD VSS sg13g2_decap_8
XFILLER_0_623 VDD VSS sg13g2_decap_8
XFILLER_75_402 VDD VSS sg13g2_decap_8
XFILLER_85_35 VDD VSS sg13g2_decap_8
XFILLER_48_616 VDD VSS sg13g2_decap_8
XFILLER_87_273 VDD VSS sg13g2_decap_8
XFILLER_47_126 VDD VSS sg13g2_decap_8
XFILLER_90_427 VDD VSS sg13g2_decap_8
XFILLER_56_693 VDD VSS sg13g2_decap_8
XFILLER_18_84 VDD VSS sg13g2_decap_8
XFILLER_83_490 VDD VSS sg13g2_decap_8
XFILLER_43_343 VDD VSS sg13g2_decap_8
XFILLER_16_546 VDD VSS sg13g2_decap_8
XFILLER_71_674 VDD VSS sg13g2_decap_8
XFILLER_70_140 VDD VSS sg13g2_decap_8
XFILLER_70_195 VDD VSS sg13g2_decap_8
XFILLER_8_756 VDD VSS sg13g2_fill_1
XFILLER_11_273 VDD VSS sg13g2_decap_8
XFILLER_7_266 VDD VSS sg13g2_decap_8
XFILLER_3_483 VDD VSS sg13g2_decap_8
XFILLER_94_700 VDD VSS sg13g2_decap_8
XFILLER_59_91 VDD VSS sg13g2_decap_8
XFILLER_39_616 VDD VSS sg13g2_decap_8
XFILLER_93_210 VDD VSS sg13g2_decap_8
XFILLER_78_273 VDD VSS sg13g2_decap_8
XFILLER_66_413 VDD VSS sg13g2_decap_8
XFILLER_38_126 VDD VSS sg13g2_decap_8
XFILLER_66_457 VDD VSS sg13g2_decap_8
XFILLER_93_287 VDD VSS sg13g2_decap_8
XFILLER_81_427 VDD VSS sg13g2_decap_8
XFILLER_47_693 VDD VSS sg13g2_decap_8
XFILLER_74_490 VDD VSS sg13g2_decap_8
XFILLER_62_630 VDD VSS sg13g2_decap_8
XFILLER_34_343 VDD VSS sg13g2_decap_8
XFILLER_61_140 VDD VSS sg13g2_decap_8
XFILLER_30_560 VDD VSS sg13g2_decap_8
XFILLER_39_28 VDD VSS sg13g2_decap_8
XFILLER_85_700 VDD VSS sg13g2_decap_8
XFILLER_69_240 VDD VSS sg13g2_fill_1
XFILLER_84_210 VDD VSS sg13g2_decap_8
XFILLER_29_126 VDD VSS sg13g2_decap_8
XFILLER_57_413 VDD VSS sg13g2_decap_8
XFILLER_84_287 VDD VSS sg13g2_decap_8
XFILLER_72_416 VDD VSS sg13g2_decap_8
XFILLER_55_49 VDD VSS sg13g2_decap_8
XFILLER_53_630 VDD VSS sg13g2_decap_8
XFILLER_25_343 VDD VSS sg13g2_decap_8
XFILLER_38_693 VDD VSS sg13g2_decap_8
XFILLER_52_140 VDD VSS sg13g2_decap_8
XFILLER_40_357 VDD VSS sg13g2_decap_8
XFILLER_21_560 VDD VSS sg13g2_decap_8
XFILLER_4_203 VDD VSS sg13g2_decap_8
XFILLER_20_63 VDD VSS sg13g2_decap_8
XFILLER_0_420 VDD VSS sg13g2_decap_8
XFILLER_88_560 VDD VSS sg13g2_decap_8
XFILLER_75_221 VDD VSS sg13g2_decap_8
XFILLER_0_497 VDD VSS sg13g2_decap_8
XFILLER_48_413 VDD VSS sg13g2_decap_8
XFILLER_76_755 VDD VSS sg13g2_fill_2
XFILLER_75_243 VDD VSS sg13g2_decap_8
XFILLER_91_714 VDD VSS sg13g2_decap_8
XFILLER_63_427 VDD VSS sg13g2_decap_8
XFILLER_90_224 VDD VSS sg13g2_decap_8
XFILLER_56_490 VDD VSS sg13g2_decap_8
XFILLER_29_693 VDD VSS sg13g2_decap_8
XFILLER_44_630 VDD VSS sg13g2_decap_8
XFILLER_16_343 VDD VSS sg13g2_decap_8
XFILLER_43_140 VDD VSS sg13g2_decap_8
XFILLER_71_471 VDD VSS sg13g2_decap_8
XFILLER_31_357 VDD VSS sg13g2_decap_8
XFILLER_84_7 VDD VSS sg13g2_decap_8
XFILLER_12_560 VDD VSS sg13g2_decap_8
XFILLER_61_70 VDD VSS sg13g2_decap_8
XFILLER_8_553 VDD VSS sg13g2_decap_8
XFILLER_6_21 VDD VSS sg13g2_decap_8
XFILLER_6_98 VDD VSS sg13g2_decap_8
XFILLER_3_280 VDD VSS sg13g2_decap_8
XFILLER_79_560 VDD VSS sg13g2_decap_8
XFILLER_67_744 VDD VSS sg13g2_decap_8
XFILLER_66_210 VDD VSS sg13g2_decap_8
XFILLER_39_413 VDD VSS sg13g2_decap_8
XFILLER_67_755 VDD VSS sg13g2_fill_2
XFILLER_94_574 VDD VSS sg13g2_decap_8
XFILLER_82_714 VDD VSS sg13g2_decap_8
XFILLER_66_287 VDD VSS sg13g2_decap_8
XFILLER_54_427 VDD VSS sg13g2_decap_8
XFILLER_81_224 VDD VSS sg13g2_decap_8
XFILLER_47_490 VDD VSS sg13g2_decap_8
XFILLER_35_630 VDD VSS sg13g2_decap_8
XFILLER_34_140 VDD VSS sg13g2_decap_8
XFILLER_50_644 VDD VSS sg13g2_decap_8
XFILLER_22_357 VDD VSS sg13g2_decap_8
XFILLER_2_707 VDD VSS sg13g2_decap_8
XFILLER_1_217 VDD VSS sg13g2_decap_8
XFILLER_89_357 VDD VSS sg13g2_decap_8
XFILLER_58_700 VDD VSS sg13g2_decap_8
XFILLER_57_210 VDD VSS sg13g2_decap_8
XFILLER_85_574 VDD VSS sg13g2_decap_8
XFILLER_45_427 VDD VSS sg13g2_decap_8
XFILLER_57_287 VDD VSS sg13g2_decap_8
XFILLER_72_224 VDD VSS sg13g2_decap_8
XFILLER_72_235 VDD VSS sg13g2_decap_8
XFILLER_82_14 VDD VSS sg13g2_decap_8
XFILLER_38_490 VDD VSS sg13g2_decap_8
XFILLER_25_140 VDD VSS sg13g2_decap_8
XFILLER_26_685 VDD VSS sg13g2_decap_8
XFILLER_13_357 VDD VSS sg13g2_decap_8
XFILLER_15_63 VDD VSS sg13g2_decap_8
XFILLER_41_644 VDD VSS sg13g2_decap_8
XFILLER_40_154 VDD VSS sg13g2_decap_8
XFILLER_31_84 VDD VSS sg13g2_decap_8
XFILLER_5_567 VDD VSS sg13g2_decap_8
XFILLER_49_700 VDD VSS sg13g2_decap_8
XFILLER_48_210 VDD VSS sg13g2_decap_8
XFILLER_76_552 VDD VSS sg13g2_decap_8
XFILLER_0_294 VDD VSS sg13g2_decap_8
XFILLER_91_511 VDD VSS sg13g2_decap_8
XFILLER_64_714 VDD VSS sg13g2_decap_8
XFILLER_36_427 VDD VSS sg13g2_decap_8
XFILLER_48_287 VDD VSS sg13g2_decap_8
XFILLER_63_224 VDD VSS sg13g2_decap_8
XFILLER_56_70 VDD VSS sg13g2_decap_8
XFILLER_17_630 VDD VSS sg13g2_decap_8
XFILLER_29_490 VDD VSS sg13g2_decap_8
XFILLER_91_588 VDD VSS sg13g2_decap_8
XFILLER_16_140 VDD VSS sg13g2_decap_8
XFILLER_32_644 VDD VSS sg13g2_decap_8
XFILLER_72_91 VDD VSS sg13g2_decap_8
XFILLER_31_154 VDD VSS sg13g2_decap_8
XFILLER_8_350 VDD VSS sg13g2_decap_8
XFILLER_39_210 VDD VSS sg13g2_decap_8
XFILLER_67_541 VDD VSS sg13g2_decap_8
XFILLER_82_511 VDD VSS sg13g2_decap_8
XFILLER_94_371 VDD VSS sg13g2_decap_8
XFILLER_55_714 VDD VSS sg13g2_decap_8
XFILLER_27_427 VDD VSS sg13g2_decap_8
XFILLER_39_287 VDD VSS sg13g2_decap_8
XFILLER_54_224 VDD VSS sg13g2_decap_8
XFILLER_82_588 VDD VSS sg13g2_decap_8
XFILLER_52_28 VDD VSS sg13g2_decap_8
XFILLER_50_441 VDD VSS sg13g2_decap_8
XFILLER_23_644 VDD VSS sg13g2_decap_8
XFILLER_22_154 VDD VSS sg13g2_decap_8
XFILLER_2_504 VDD VSS sg13g2_decap_8
XFILLER_89_154 VDD VSS sg13g2_decap_8
XFILLER_77_14 VDD VSS sg13g2_decap_8
XFILLER_77_316 VDD VSS sg13g2_decap_8
XFILLER_92_308 VDD VSS sg13g2_decap_8
XFILLER_85_371 VDD VSS sg13g2_decap_8
XFILLER_58_574 VDD VSS sg13g2_decap_8
XFILLER_46_714 VDD VSS sg13g2_decap_8
XFILLER_93_35 VDD VSS sg13g2_decap_8
Xoutputs\[6\].output_pad _82_/Q IOVDD IOVSS output_PAD[6] VDD VSS sg13g2_IOPadOut30mA
XFILLER_18_427 VDD VSS sg13g2_decap_8
XFILLER_45_224 VDD VSS sg13g2_decap_8
XFILLER_73_555 VDD VSS sg13g2_decap_8
XFILLER_61_728 VDD VSS sg13g2_decap_8
XFILLER_26_84 VDD VSS sg13g2_decap_8
XFILLER_26_482 VDD VSS sg13g2_decap_8
XFILLER_60_238 VDD VSS sg13g2_decap_8
XFILLER_41_441 VDD VSS sg13g2_decap_8
XFILLER_14_644 VDD VSS sg13g2_decap_8
XFILLER_13_154 VDD VSS sg13g2_decap_8
XFILLER_9_147 VDD VSS sg13g2_decap_8
XFILLER_5_364 VDD VSS sg13g2_decap_8
XFILLER_47_7 VDD VSS sg13g2_decap_8
XFILLER_68_349 VDD VSS sg13g2_decap_8
XFILLER_1_581 VDD VSS sg13g2_decap_8
XFILLER_3_77 VDD VSS sg13g2_decap_8
XFILLER_64_511 VDD VSS sg13g2_decap_8
XFILLER_95_168 VDD VSS sg13g2_decap_8
XFILLER_83_308 VDD VSS sg13g2_decap_8
XFILLER_67_91 VDD VSS sg13g2_decap_8
XFILLER_49_574 VDD VSS sg13g2_decap_8
XFILLER_37_714 VDD VSS sg13g2_decap_8
XFILLER_36_224 VDD VSS sg13g2_decap_8
XFILLER_64_588 VDD VSS sg13g2_decap_8
XFILLER_91_385 VDD VSS sg13g2_decap_8
XFILLER_52_728 VDD VSS sg13g2_decap_8
XFILLER_32_441 VDD VSS sg13g2_decap_8
XFILLER_51_238 VDD VSS sg13g2_decap_8
XFILLER_20_658 VDD VSS sg13g2_decap_8
XFILLER_73_0 VDD VSS sg13g2_decap_8
XFILLER_87_658 VDD VSS sg13g2_decap_8
XFILLER_47_28 VDD VSS sg13g2_decap_8
XFILLER_86_168 VDD VSS sg13g2_decap_8
XFILLER_28_714 VDD VSS sg13g2_decap_8
XFILLER_55_511 VDD VSS sg13g2_decap_8
XFILLER_27_224 VDD VSS sg13g2_decap_8
XFILLER_82_385 VDD VSS sg13g2_decap_8
XFILLER_63_49 VDD VSS sg13g2_decap_8
XFILLER_55_588 VDD VSS sg13g2_decap_8
XFILLER_43_728 VDD VSS sg13g2_decap_8
XFILLER_70_547 VDD VSS sg13g2_decap_8
XFILLER_23_441 VDD VSS sg13g2_decap_8
XFILLER_42_238 VDD VSS sg13g2_decap_8
XFILLER_11_658 VDD VSS sg13g2_decap_8
XFILLER_10_168 VDD VSS sg13g2_decap_8
XFILLER_12_42 VDD VSS sg13g2_decap_8
XFILLER_88_35 VDD VSS sg13g2_decap_8
XFILLER_2_301 VDD VSS sg13g2_decap_8
XFILLER_2_378 VDD VSS sg13g2_decap_8
XFILLER_78_658 VDD VSS sg13g2_decap_8
XFILLER_77_168 VDD VSS sg13g2_decap_8
XFILLER_65_308 VDD VSS sg13g2_decap_8
XFILLER_92_105 VDD VSS sg13g2_decap_8
XFILLER_19_714 VDD VSS sg13g2_decap_8
XFILLER_46_511 VDD VSS sg13g2_decap_8
XFILLER_18_224 VDD VSS sg13g2_decap_8
XFILLER_58_371 VDD VSS sg13g2_decap_8
XFILLER_73_374 VDD VSS sg13g2_decap_8
XFILLER_61_525 VDD VSS sg13g2_decap_8
XFILLER_46_588 VDD VSS sg13g2_decap_8
XFILLER_34_728 VDD VSS sg13g2_decap_8
XFILLER_14_441 VDD VSS sg13g2_decap_8
XFILLER_33_238 VDD VSS sg13g2_decap_8
XFILLER_6_651 VDD VSS sg13g2_decap_8
XFILLER_5_161 VDD VSS sg13g2_decap_8
XFILLER_69_636 VDD VSS sg13g2_decap_8
XFILLER_68_168 VDD VSS sg13g2_decap_8
XFILLER_83_105 VDD VSS sg13g2_decap_8
XFILLER_56_308 VDD VSS sg13g2_decap_8
XFILLER_49_371 VDD VSS sg13g2_decap_8
XFILLER_37_511 VDD VSS sg13g2_decap_8
X_67_ _80_/D _75_/A _67_/B _74_/D VDD VSS sg13g2_and3_1
XFILLER_92_672 VDD VSS sg13g2_decap_8
XFILLER_64_385 VDD VSS sg13g2_decap_8
XFILLER_52_525 VDD VSS sg13g2_decap_8
XFILLER_25_728 VDD VSS sg13g2_decap_8
XFILLER_37_588 VDD VSS sg13g2_decap_8
XFILLER_91_182 VDD VSS sg13g2_decap_8
XFILLER_24_238 VDD VSS sg13g2_decap_8
XFILLER_20_455 VDD VSS sg13g2_decap_8
XFILLER_87_455 VDD VSS sg13g2_decap_8
XFILLER_58_49 VDD VSS sg13g2_decap_8
XFILLER_75_606 VDD VSS sg13g2_decap_8
XFILLER_74_105 VDD VSS sg13g2_decap_8
XFILLER_47_308 VDD VSS sg13g2_decap_8
XFILLER_59_168 VDD VSS sg13g2_decap_8
XFILLER_28_511 VDD VSS sg13g2_decap_8
XFILLER_90_609 VDD VSS sg13g2_decap_8
XFILLER_83_672 VDD VSS sg13g2_decap_8
XFILLER_55_385 VDD VSS sg13g2_decap_8
XFILLER_16_728 VDD VSS sg13g2_decap_8
XFILLER_28_588 VDD VSS sg13g2_decap_8
XFILLER_43_525 VDD VSS sg13g2_decap_8
XFILLER_82_182 VDD VSS sg13g2_decap_8
XFILLER_15_238 VDD VSS sg13g2_decap_8
XFILLER_70_355 VDD VSS sg13g2_decap_8
XFILLER_90_14 VDD VSS sg13g2_decap_8
XFILLER_11_455 VDD VSS sg13g2_decap_8
XFILLER_23_63 VDD VSS sg13g2_decap_8
XFILLER_7_448 VDD VSS sg13g2_decap_8
XFILLER_3_0 VDD VSS sg13g2_decap_8
XFILLER_3_665 VDD VSS sg13g2_decap_8
XFILLER_2_175 VDD VSS sg13g2_decap_8
XFILLER_78_455 VDD VSS sg13g2_decap_8
XFILLER_65_105 VDD VSS sg13g2_decap_8
XFILLER_38_308 VDD VSS sg13g2_decap_8
XFILLER_66_639 VDD VSS sg13g2_decap_8
XFILLER_19_511 VDD VSS sg13g2_decap_8
XFILLER_81_609 VDD VSS sg13g2_decap_8
XFILLER_93_469 VDD VSS sg13g2_decap_8
XFILLER_74_672 VDD VSS sg13g2_decap_8
XFILLER_80_119 VDD VSS sg13g2_decap_8
XFILLER_0_56 VDD VSS sg13g2_decap_8
XFILLER_46_385 VDD VSS sg13g2_decap_8
XFILLER_19_588 VDD VSS sg13g2_decap_8
XFILLER_34_525 VDD VSS sg13g2_decap_8
XFILLER_73_182 VDD VSS sg13g2_decap_8
XFILLER_64_70 VDD VSS sg13g2_decap_8
XFILLER_61_322 VDD VSS sg13g2_decap_8
XFILLER_9_21 VDD VSS sg13g2_decap_8
XFILLER_61_399 VDD VSS sg13g2_decap_8
XFILLER_30_742 VDD VSS sg13g2_decap_8
XFILLER_80_91 VDD VSS sg13g2_decap_8
XFILLER_9_98 VDD VSS sg13g2_decap_8
XFILLER_69_422 VDD VSS sg13g2_decap_8
XFILLER_36_0 VDD VSS sg13g2_decap_8
XFILLER_29_308 VDD VSS sg13g2_decap_8
XFILLER_56_105 VDD VSS sg13g2_decap_8
XFILLER_84_469 VDD VSS sg13g2_decap_8
XFILLER_65_661 VDD VSS sg13g2_decap_8
XFILLER_71_119 VDD VSS sg13g2_decap_8
XFILLER_37_385 VDD VSS sg13g2_decap_8
XFILLER_25_525 VDD VSS sg13g2_decap_8
XFILLER_64_182 VDD VSS sg13g2_decap_8
XFILLER_52_322 VDD VSS sg13g2_decap_8
XFILLER_80_686 VDD VSS sg13g2_decap_8
XFILLER_52_399 VDD VSS sg13g2_decap_8
XFILLER_40_539 VDD VSS sg13g2_decap_8
XIO_BOND_rst_n_pad rst_n_PAD bondpad_70x70_novias
XFILLER_60_28 VDD VSS sg13g2_decap_8
XFILLER_21_742 VDD VSS sg13g2_decap_8
XFILLER_20_252 VDD VSS sg13g2_decap_8
XFILLER_0_602 VDD VSS sg13g2_decap_8
XFILLER_88_742 VDD VSS sg13g2_decap_8
XFILLER_87_252 VDD VSS sg13g2_decap_8
XFILLER_85_14 VDD VSS sg13g2_decap_8
XFILLER_0_679 VDD VSS sg13g2_decap_8
XFILLER_47_105 VDD VSS sg13g2_decap_8
XFILLER_90_406 VDD VSS sg13g2_decap_8
XFILLER_62_119 VDD VSS sg13g2_decap_8
XFILLER_56_672 VDD VSS sg13g2_decap_8
XFILLER_18_63 VDD VSS sg13g2_decap_8
XFILLER_16_525 VDD VSS sg13g2_decap_8
XFILLER_71_653 VDD VSS sg13g2_decap_8
XFILLER_28_385 VDD VSS sg13g2_decap_8
XFILLER_43_322 VDD VSS sg13g2_decap_8
XFILLER_55_182 VDD VSS sg13g2_decap_8
XFILLER_43_399 VDD VSS sg13g2_decap_8
XFILLER_31_539 VDD VSS sg13g2_decap_8
XFILLER_12_742 VDD VSS sg13g2_decap_8
XFILLER_34_84 VDD VSS sg13g2_decap_8
XFILLER_8_735 VDD VSS sg13g2_decap_8
XFILLER_11_252 VDD VSS sg13g2_decap_8
XFILLER_7_245 VDD VSS sg13g2_decap_8
Xclkbuf_1_1__f_clk_PAD2CORE _83_/CLK clkbuf_0_clk_PAD2CORE/X VDD VSS sg13g2_buf_16
XFILLER_3_462 VDD VSS sg13g2_decap_8
XFILLER_79_742 VDD VSS sg13g2_decap_8
XFILLER_59_70 VDD VSS sg13g2_decap_8
XFILLER_78_252 VDD VSS sg13g2_decap_8
XFILLER_38_105 VDD VSS sg13g2_decap_8
XFILLER_94_756 VDD VSS sg13g2_fill_1
XFILLER_54_609 VDD VSS sg13g2_decap_8
XFILLER_93_266 VDD VSS sg13g2_decap_8
XFILLER_81_406 VDD VSS sg13g2_decap_8
XFILLER_47_672 VDD VSS sg13g2_decap_8
XFILLER_53_119 VDD VSS sg13g2_decap_8
XFILLER_19_385 VDD VSS sg13g2_decap_8
XFILLER_34_322 VDD VSS sg13g2_decap_8
XFILLER_46_182 VDD VSS sg13g2_decap_8
XFILLER_62_686 VDD VSS sg13g2_decap_8
XFILLER_34_399 VDD VSS sg13g2_decap_8
XFILLER_61_196 VDD VSS sg13g2_decap_8
XFILLER_22_539 VDD VSS sg13g2_decap_8
XFILLER_89_539 VDD VSS sg13g2_decap_8
XFILLER_69_296 VDD VSS sg13g2_decap_8
XFILLER_29_105 VDD VSS sg13g2_decap_8
XFILLER_85_756 VDD VSS sg13g2_fill_1
XFILLER_57_469 VDD VSS sg13g2_decap_8
XFILLER_45_609 VDD VSS sg13g2_decap_8
XFILLER_84_266 VDD VSS sg13g2_decap_8
XFILLER_55_28 VDD VSS sg13g2_decap_8
XFILLER_44_119 VDD VSS sg13g2_decap_8
XFILLER_38_672 VDD VSS sg13g2_decap_8
XFILLER_72_439 VDD VSS sg13g2_decap_8
XFILLER_25_322 VDD VSS sg13g2_decap_8
XFILLER_37_182 VDD VSS sg13g2_decap_8
XFILLER_80_483 VDD VSS sg13g2_decap_8
XFILLER_53_686 VDD VSS sg13g2_decap_8
XFILLER_13_539 VDD VSS sg13g2_decap_8
XFILLER_25_399 VDD VSS sg13g2_decap_8
XFILLER_71_49 VDD VSS sg13g2_decap_8
XFILLER_40_336 VDD VSS sg13g2_decap_8
XFILLER_52_196 VDD VSS sg13g2_decap_8
XFILLER_5_749 VDD VSS sg13g2_decap_8
XFILLER_20_42 VDD VSS sg13g2_decap_8
XFILLER_4_259 VDD VSS sg13g2_decap_8
XFILLER_76_734 VDD VSS sg13g2_decap_8
XFILLER_75_200 VDD VSS sg13g2_decap_8
XFILLER_0_476 VDD VSS sg13g2_decap_8
XFILLER_29_84 VDD VSS sg13g2_decap_8
XFILLER_48_469 VDD VSS sg13g2_decap_8
XFILLER_36_609 VDD VSS sg13g2_decap_8
XFILLER_90_203 VDD VSS sg13g2_decap_8
XFILLER_63_406 VDD VSS sg13g2_decap_8
XFILLER_35_119 VDD VSS sg13g2_decap_8
XFILLER_29_672 VDD VSS sg13g2_decap_8
XFILLER_16_322 VDD VSS sg13g2_decap_8
XFILLER_28_182 VDD VSS sg13g2_decap_8
XFILLER_71_450 VDD VSS sg13g2_decap_8
XFILLER_16_399 VDD VSS sg13g2_decap_8
XFILLER_44_686 VDD VSS sg13g2_decap_8
XFILLER_31_336 VDD VSS sg13g2_decap_8
XFILLER_43_196 VDD VSS sg13g2_decap_8
XFILLER_77_7 VDD VSS sg13g2_decap_8
XFILLER_8_532 VDD VSS sg13g2_decap_8
XFILLER_6_77 VDD VSS sg13g2_decap_8
XFILLER_67_723 VDD VSS sg13g2_decap_8
XFILLER_94_553 VDD VSS sg13g2_decap_8
XFILLER_39_469 VDD VSS sg13g2_decap_8
XFILLER_27_609 VDD VSS sg13g2_decap_8
XFILLER_81_203 VDD VSS sg13g2_decap_8
XFILLER_66_266 VDD VSS sg13g2_decap_8
XFILLER_26_119 VDD VSS sg13g2_decap_8
XFILLER_54_406 VDD VSS sg13g2_decap_8
XFILLER_19_182 VDD VSS sg13g2_decap_8
XFILLER_62_483 VDD VSS sg13g2_decap_8
XFILLER_50_623 VDD VSS sg13g2_decap_8
XFILLER_35_686 VDD VSS sg13g2_decap_8
XFILLER_22_336 VDD VSS sg13g2_decap_8
XFILLER_34_196 VDD VSS sg13g2_decap_8
XFILLER_89_336 VDD VSS sg13g2_decap_8
XFILLER_85_553 VDD VSS sg13g2_decap_8
XFILLER_66_49 VDD VSS sg13g2_decap_8
XFILLER_58_756 VDD VSS sg13g2_fill_1
XFILLER_18_609 VDD VSS sg13g2_decap_8
XFILLER_72_203 VDD VSS sg13g2_decap_8
XFILLER_45_406 VDD VSS sg13g2_decap_8
XFILLER_57_266 VDD VSS sg13g2_decap_8
XFILLER_73_737 VDD VSS sg13g2_decap_8
XFILLER_17_119 VDD VSS sg13g2_decap_8
XFILLER_26_664 VDD VSS sg13g2_decap_8
XFILLER_53_483 VDD VSS sg13g2_decap_8
XFILLER_41_623 VDD VSS sg13g2_decap_8
XFILLER_80_280 VDD VSS sg13g2_decap_8
XFILLER_13_336 VDD VSS sg13g2_decap_8
XFILLER_15_42 VDD VSS sg13g2_decap_8
XFILLER_25_196 VDD VSS sg13g2_decap_8
XFILLER_40_133 VDD VSS sg13g2_decap_8
XFILLER_9_329 VDD VSS sg13g2_decap_8
XFILLER_5_546 VDD VSS sg13g2_decap_8
XFILLER_31_63 VDD VSS sg13g2_decap_8
XFILLER_0_273 VDD VSS sg13g2_decap_8
XFILLER_76_531 VDD VSS sg13g2_decap_8
XFILLER_49_756 VDD VSS sg13g2_fill_1
XFILLER_63_203 VDD VSS sg13g2_decap_8
XFILLER_36_406 VDD VSS sg13g2_decap_8
XFILLER_48_266 VDD VSS sg13g2_decap_8
XFILLER_91_567 VDD VSS sg13g2_decap_8
XFILLER_17_686 VDD VSS sg13g2_decap_8
XFILLER_32_623 VDD VSS sg13g2_decap_8
XFILLER_44_483 VDD VSS sg13g2_decap_8
XFILLER_72_70 VDD VSS sg13g2_decap_8
XFILLER_16_196 VDD VSS sg13g2_decap_8
XFILLER_31_133 VDD VSS sg13g2_decap_8
.ends

