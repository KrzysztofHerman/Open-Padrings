module FMD_QNC_Padframe24 (clk_PAD,
    rst_n_PAD,
    VDD,
    VSS,
    IOVSS,
    IOVDD,
    input_PAD,
    output_PAD);
 inout clk_PAD;
 inout rst_n_PAD;
 inout VDD;
 inout VSS;
 inout IOVSS;
 inout IOVDD;
 inout [7:0] input_PAD;
 inout [9:0] output_PAD;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_0_clk_PAD2CORE;
 wire net1;
 wire net2;
 wire clk_PAD2CORE;
 wire \i_chip_core.count[0] ;
 wire \i_chip_core.count[1] ;
 wire \i_chip_core.count[2] ;
 wire \i_chip_core.count[3] ;
 wire \i_chip_core.count[4] ;
 wire \i_chip_core.count[5] ;
 wire \i_chip_core.count[6] ;
 wire \i_chip_core.count[7] ;
 wire \i_chip_core.input_in[0] ;
 wire \i_chip_core.input_in[1] ;
 wire \i_chip_core.input_in[2] ;
 wire \i_chip_core.input_in[3] ;
 wire \i_chip_core.input_in[4] ;
 wire \i_chip_core.input_in[5] ;
 wire \i_chip_core.input_in[6] ;
 wire \i_chip_core.input_in[7] ;
 wire \i_chip_core.rst_n ;
 wire net;
 wire clknet_1_0__leaf_clk_PAD2CORE;
 wire clknet_1_1__leaf_clk_PAD2CORE;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;

 sg13g2_inv_1 _43_ (.VDD(VDD),
    .Y(_08_),
    .A(net21),
    .VSS(VSS));
 sg13g2_inv_1 _44_ (.VDD(VDD),
    .Y(_09_),
    .A(\i_chip_core.count[6] ),
    .VSS(VSS));
 sg13g2_inv_1 _45_ (.VDD(VDD),
    .Y(_10_),
    .A(net19),
    .VSS(VSS));
 sg13g2_inv_1 _46_ (.VDD(VDD),
    .Y(_11_),
    .A(\i_chip_core.count[2] ),
    .VSS(VSS));
 sg13g2_inv_1 _47_ (.VDD(VDD),
    .Y(_12_),
    .A(net10),
    .VSS(VSS));
 sg13g2_nand4_1 _48_ (.B(\i_chip_core.input_in[4] ),
    .C(\i_chip_core.input_in[7] ),
    .A(\i_chip_core.input_in[5] ),
    .Y(_13_),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_chip_core.input_in[6] ));
 sg13g2_nand4_1 _49_ (.B(\i_chip_core.input_in[0] ),
    .C(\i_chip_core.input_in[3] ),
    .A(net13),
    .Y(_14_),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_chip_core.input_in[2] ));
 sg13g2_nor2_1 _50_ (.A(_13_),
    .B(net14),
    .Y(_15_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _51_ (.B(\i_chip_core.input_in[3] ),
    .C(\i_chip_core.input_in[5] ),
    .A(\i_chip_core.input_in[0] ),
    .Y(_16_),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_chip_core.input_in[6] ));
 sg13g2_nand4_1 _52_ (.B(net27),
    .C(\i_chip_core.input_in[4] ),
    .A(net13),
    .Y(_17_),
    .VDD(VDD),
    .VSS(VSS),
    .D(\i_chip_core.input_in[7] ));
 sg13g2_o21ai_1 _53_ (.B1(net10),
    .VDD(VDD),
    .Y(_18_),
    .VSS(VSS),
    .A1(\i_chip_core.count[0] ),
    .A2(net15));
 sg13g2_a21oi_1 _54_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_chip_core.count[0] ),
    .A2(net15),
    .Y(_00_),
    .B1(_18_));
 sg13g2_a21oi_1 _55_ (.VSS(VSS),
    .VDD(VDD),
    .A1(\i_chip_core.count[0] ),
    .A2(net15),
    .Y(_19_),
    .B1(\i_chip_core.count[1] ));
 sg13g2_nand2_1 _56_ (.Y(_20_),
    .A(\i_chip_core.count[1] ),
    .B(\i_chip_core.count[0] ),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _57_ (.A(_16_),
    .B(net28),
    .C(_20_),
    .Y(_21_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _58_ (.A(_12_),
    .B(_19_),
    .C(net29),
    .Y(_01_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor2_1 _59_ (.A(net24),
    .B(_21_),
    .Y(_22_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor4_1 _60_ (.A(_11_),
    .B(_13_),
    .C(net14),
    .D(_20_),
    .Y(_23_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nor3_1 _61_ (.A(_12_),
    .B(net25),
    .C(_23_),
    .Y(_02_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand3_1 _62_ (.B(\i_chip_core.count[2] ),
    .C(_21_),
    .A(net17),
    .Y(_24_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_o21ai_1 _63_ (.B1(net10),
    .VDD(VDD),
    .Y(_25_),
    .VSS(VSS),
    .A1(net17),
    .A2(_23_));
 sg13g2_nor2b_1 _64_ (.A(_25_),
    .B_N(_24_),
    .Y(_03_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand2b_1 _65_ (.Y(_26_),
    .B(_24_),
    .A_N(net22),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _66_ (.B(net17),
    .C(\i_chip_core.count[2] ),
    .A(\i_chip_core.count[4] ),
    .Y(_27_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_21_));
 sg13g2_and3_1 _67_ (.X(_04_),
    .A(net10),
    .B(net23),
    .C(_27_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_nand4_1 _68_ (.B(\i_chip_core.count[4] ),
    .C(\i_chip_core.count[3] ),
    .A(\i_chip_core.count[5] ),
    .Y(_28_),
    .VDD(VDD),
    .VSS(VSS),
    .D(_23_));
 sg13g2_nand2_1 _69_ (.Y(_29_),
    .A(net10),
    .B(_28_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_a21oi_1 _70_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_10_),
    .A2(_27_),
    .Y(_05_),
    .B1(_29_));
 sg13g2_o21ai_1 _71_ (.B1(net10),
    .VDD(VDD),
    .Y(_30_),
    .VSS(VSS),
    .A1(_09_),
    .A2(_28_));
 sg13g2_a21oi_1 _72_ (.VSS(VSS),
    .VDD(VDD),
    .A1(_09_),
    .A2(_28_),
    .Y(_06_),
    .B1(net11));
 sg13g2_o21ai_1 _73_ (.B1(_08_),
    .VDD(VDD),
    .Y(_31_),
    .VSS(VSS),
    .A1(_09_),
    .A2(_28_));
 sg13g2_or4_1 _74_ (.A(_08_),
    .B(_09_),
    .C(_10_),
    .D(_27_),
    .X(_32_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_and3_1 _75_ (.X(_07_),
    .A(net10),
    .B(_31_),
    .C(_32_),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dfrbpq_1 _76_ (.RESET_B(net2),
    .VSS(VSS),
    .VDD(VDD),
    .D(net16),
    .Q(\i_chip_core.count[0] ),
    .CLK(clknet_1_0__leaf_clk_PAD2CORE));
 sg13g2_dfrbpq_1 _77_ (.RESET_B(net9),
    .VSS(VSS),
    .VDD(VDD),
    .D(net30),
    .Q(\i_chip_core.count[1] ),
    .CLK(clknet_1_0__leaf_clk_PAD2CORE));
 sg13g2_dfrbpq_1 _78_ (.RESET_B(net7),
    .VSS(VSS),
    .VDD(VDD),
    .D(net26),
    .Q(\i_chip_core.count[2] ),
    .CLK(clknet_1_0__leaf_clk_PAD2CORE));
 sg13g2_dfrbpq_1 _79_ (.RESET_B(net5),
    .VSS(VSS),
    .VDD(VDD),
    .D(net18),
    .Q(\i_chip_core.count[3] ),
    .CLK(clknet_1_0__leaf_clk_PAD2CORE));
 sg13g2_dfrbpq_1 _80_ (.RESET_B(net3),
    .VSS(VSS),
    .VDD(VDD),
    .D(_04_),
    .Q(\i_chip_core.count[4] ),
    .CLK(clknet_1_1__leaf_clk_PAD2CORE));
 sg13g2_dfrbpq_1 _81_ (.RESET_B(net8),
    .VSS(VSS),
    .VDD(VDD),
    .D(net20),
    .Q(\i_chip_core.count[5] ),
    .CLK(clknet_1_1__leaf_clk_PAD2CORE));
 sg13g2_dfrbpq_1 _82_ (.RESET_B(net4),
    .VSS(VSS),
    .VDD(VDD),
    .D(net12),
    .Q(\i_chip_core.count[6] ),
    .CLK(clknet_1_1__leaf_clk_PAD2CORE));
 sg13g2_dfrbpq_1 _83_ (.RESET_B(net6),
    .VSS(VSS),
    .VDD(VDD),
    .D(_07_),
    .Q(\i_chip_core.count[7] ),
    .CLK(clknet_1_1__leaf_clk_PAD2CORE));
 sg13g2_tiehi _80__4 (.VDD(VDD),
    .VSS(VSS),
    .L_HI(net3));
 sg13g2_tiehi _82__5 (.VDD(VDD),
    .VSS(VSS),
    .L_HI(net4));
 sg13g2_tiehi _79__6 (.VDD(VDD),
    .VSS(VSS),
    .L_HI(net5));
 sg13g2_tiehi _83__7 (.VDD(VDD),
    .VSS(VSS),
    .L_HI(net6));
 sg13g2_tiehi _78__8 (.VDD(VDD),
    .VSS(VSS),
    .L_HI(net7));
 sg13g2_tiehi _81__9 (.VDD(VDD),
    .VSS(VSS),
    .L_HI(net8));
 sg13g2_tiehi _77__10 (.VDD(VDD),
    .VSS(VSS),
    .L_HI(net9));
 sg13g2_buf_16 clkbuf_0_clk_PAD2CORE (.X(clknet_0_clk_PAD2CORE),
    .A(clk_PAD2CORE),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_tielo \outputs[9].output_pad_2  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net1));
 sg13g2_tiehi _76__3 (.VDD(VDD),
    .VSS(VSS),
    .L_HI(net2));
 sg13g2_IOPadIn clk_pad (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(clk_PAD2CORE),
    .pad(clk_PAD),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \inputs[0].input_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\i_chip_core.input_in[0] ),
    .pad(input_PAD[0]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \inputs[1].input_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\i_chip_core.input_in[1] ),
    .pad(input_PAD[1]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \inputs[2].input_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\i_chip_core.input_in[2] ),
    .pad(input_PAD[2]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \inputs[3].input_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\i_chip_core.input_in[3] ),
    .pad(input_PAD[3]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \inputs[4].input_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\i_chip_core.input_in[4] ),
    .pad(input_PAD[4]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \inputs[5].input_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\i_chip_core.input_in[5] ),
    .pad(input_PAD[5]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \inputs[6].input_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\i_chip_core.input_in[6] ),
    .pad(input_PAD[6]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn \inputs[7].input_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\i_chip_core.input_in[7] ),
    .pad(input_PAD[7]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIOVdd \iovdd_pads[0].iovdd_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIOVss \iovss_pads[0].iovss_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \outputs[0].output_pad  (.c2p(\i_chip_core.count[0] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(output_PAD[0]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \outputs[1].output_pad  (.c2p(\i_chip_core.count[1] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(output_PAD[1]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \outputs[2].output_pad  (.c2p(\i_chip_core.count[2] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(output_PAD[2]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \outputs[3].output_pad  (.c2p(\i_chip_core.count[3] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(output_PAD[3]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \outputs[4].output_pad  (.c2p(\i_chip_core.count[4] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(output_PAD[4]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \outputs[5].output_pad  (.c2p(\i_chip_core.count[5] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(output_PAD[5]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \outputs[6].output_pad  (.c2p(\i_chip_core.count[6] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(output_PAD[6]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \outputs[7].output_pad  (.c2p(\i_chip_core.count[7] ),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(output_PAD[7]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \outputs[8].output_pad  (.c2p(net),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(output_PAD[8]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadOut30mA \outputs[9].output_pad  (.c2p(net1),
    .iovdd(IOVDD),
    .iovss(IOVSS),
    .pad(output_PAD[9]),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadIn rst_n_pad (.iovdd(IOVDD),
    .iovss(IOVSS),
    .p2c(\i_chip_core.rst_n ),
    .pad(rst_n_PAD),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadVdd \vdd_pads[0].vdd_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_IOPadVss \vss_pads[0].vss_pad  (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_Corner IO_CORNER_NORTH_WEST_INST (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_Corner IO_CORNER_NORTH_EAST_INST (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_Corner IO_CORNER_SOUTH_WEST_INST (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 sg13g2_Corner IO_CORNER_SOUTH_EAST_INST (.iovdd(IOVDD),
    .iovss(IOVSS),
    .vdd(VDD),
    .vss(VSS));
 bondpad_70x70_novias IO_BOND_clk_pad (.pad(clk_PAD));
 bondpad_70x70_novias IO_BOND_rst_n_pad (.pad(rst_n_PAD));
 bondpad_70x70_novias \IO_BOND_inputs[7].input_pad  (.pad(input_PAD[7]));
 bondpad_70x70_novias \IO_BOND_inputs[6].input_pad  (.pad(input_PAD[6]));
 bondpad_70x70_novias \IO_BOND_vdd_pads[0].vdd_pad  (.pad(VDD));
 bondpad_70x70_novias \IO_BOND_vss_pads[0].vss_pad  (.pad(VSS));
 bondpad_70x70_novias \IO_BOND_outputs[9].output_pad  (.pad(output_PAD[9]));
 bondpad_70x70_novias \IO_BOND_outputs[8].output_pad  (.pad(output_PAD[8]));
 bondpad_70x70_novias \IO_BOND_outputs[7].output_pad  (.pad(output_PAD[7]));
 bondpad_70x70_novias \IO_BOND_outputs[6].output_pad  (.pad(output_PAD[6]));
 bondpad_70x70_novias \IO_BOND_outputs[5].output_pad  (.pad(output_PAD[5]));
 bondpad_70x70_novias \IO_BOND_outputs[4].output_pad  (.pad(output_PAD[4]));
 bondpad_70x70_novias \IO_BOND_iovss_pads[0].iovss_pad  (.pad(IOVSS));
 bondpad_70x70_novias \IO_BOND_iovdd_pads[0].iovdd_pad  (.pad(IOVDD));
 bondpad_70x70_novias \IO_BOND_outputs[3].output_pad  (.pad(output_PAD[3]));
 bondpad_70x70_novias \IO_BOND_outputs[2].output_pad  (.pad(output_PAD[2]));
 bondpad_70x70_novias \IO_BOND_outputs[1].output_pad  (.pad(output_PAD[1]));
 bondpad_70x70_novias \IO_BOND_outputs[0].output_pad  (.pad(output_PAD[0]));
 bondpad_70x70_novias \IO_BOND_inputs[5].input_pad  (.pad(input_PAD[5]));
 bondpad_70x70_novias \IO_BOND_inputs[4].input_pad  (.pad(input_PAD[4]));
 bondpad_70x70_novias \IO_BOND_inputs[3].input_pad  (.pad(input_PAD[3]));
 bondpad_70x70_novias \IO_BOND_inputs[2].input_pad  (.pad(input_PAD[2]));
 bondpad_70x70_novias \IO_BOND_inputs[1].input_pad  (.pad(input_PAD[1]));
 bondpad_70x70_novias \IO_BOND_inputs[0].input_pad  (.pad(input_PAD[0]));
 sg13g2_tielo \outputs[8].output_pad_1  (.VDD(VDD),
    .VSS(VSS),
    .L_LO(net));
 sg13g2_buf_16 clkbuf_1_0__f_clk_PAD2CORE (.X(clknet_1_0__leaf_clk_PAD2CORE),
    .A(clknet_0_clk_PAD2CORE),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_buf_16 clkbuf_1_1__f_clk_PAD2CORE (.X(clknet_1_1__leaf_clk_PAD2CORE),
    .A(clknet_0_clk_PAD2CORE),
    .VDD(VDD),
    .VSS(VSS));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_chip_core.rst_n ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net10));
 sg13g2_dlygate4sd3_1 hold12 (.A(_30_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net11));
 sg13g2_dlygate4sd3_1 hold13 (.A(_06_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net12));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_chip_core.input_in[1] ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net13));
 sg13g2_dlygate4sd3_1 hold15 (.A(_14_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net14));
 sg13g2_dlygate4sd3_1 hold16 (.A(_15_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net15));
 sg13g2_dlygate4sd3_1 hold17 (.A(_00_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net16));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i_chip_core.count[3] ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net17));
 sg13g2_dlygate4sd3_1 hold19 (.A(_03_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net18));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_chip_core.count[5] ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold21 (.A(_05_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_chip_core.count[7] ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold23 (.A(\i_chip_core.count[4] ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold24 (.A(_26_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_chip_core.count[2] ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold26 (.A(_22_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold27 (.A(_02_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_chip_core.input_in[2] ),
    .VDD(VDD),
    .VSS(VSS),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold29 (.A(_17_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold30 (.A(_21_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold31 (.A(_01_),
    .VDD(VDD),
    .VSS(VSS),
    .X(net30));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_0_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_1_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_1_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_2_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_2_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_3_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_3_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_4_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_4_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_5_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_5_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_6_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_6_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_7_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_7_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_8_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_8_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_9_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_9_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_10_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_10_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_11_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_11_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_12_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_12_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_13_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_13_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_14_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_14_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_15_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_15_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_16_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_16_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_17_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_17_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_18_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_18_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_19_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_19_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_20_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_20_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_21_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_21_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_22_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_22_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_23_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_23_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_24_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_24_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_25_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_25_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_26_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_300 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_307 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_314 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_321 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_328 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_335 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_342 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_349 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_356 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_363 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_370 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_377 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_384 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_391 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_398 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_405 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_412 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_419 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_426 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_433 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_440 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_447 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_454 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_461 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_468 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_475 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_482 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_489 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_496 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_503 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_510 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_517 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_524 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_531 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_538 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_545 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_552 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_559 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_566 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_573 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_580 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_587 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_594 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_601 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_608 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_615 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_622 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_629 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_636 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_643 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_650 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_657 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_664 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_671 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_678 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_685 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_692 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_699 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_706 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_713 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_720 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_727 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_734 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_741 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_26_748 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_26_755 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_27_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_27_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_28_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_28_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_29_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_29_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_30_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_30_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_31_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_31_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_32_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_32_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_33_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_33_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_34_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_34_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_35_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_35_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_36_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_36_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_37_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_37_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_38_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_38_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_39_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_39_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_40_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_40_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_41_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_41_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_42_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_42_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_43_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_43_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_44_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_44_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_45_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_45_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_46_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_46_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_47_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_47_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_48_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_48_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_49_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_49_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_50_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_50_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_51_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_51_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_52_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_52_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_53_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_53_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_54_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_54_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_55_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_55_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_56_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_56_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_57_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_57_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_58_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_58_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_59_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_59_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_60_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_60_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_61_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_61_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_62_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_62_457 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_62_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_62_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_63_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_63_452 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_480 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_487 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_494 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_501 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_508 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_515 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_522 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_529 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_536 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_543 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_550 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_557 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_564 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_571 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_578 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_585 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_592 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_599 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_606 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_613 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_620 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_627 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_634 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_641 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_648 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_655 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_662 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_669 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_676 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_683 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_690 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_697 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_704 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_711 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_718 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_725 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_732 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_739 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_63_746 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_63_753 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_64_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_64_32 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_64_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_64_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_65_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_65_471 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_65_475 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_486 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_493 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_500 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_507 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_514 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_521 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_528 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_535 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_542 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_549 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_556 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_563 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_570 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_577 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_584 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_591 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_598 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_605 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_612 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_619 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_626 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_633 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_640 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_647 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_654 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_661 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_668 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_675 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_682 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_689 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_696 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_703 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_710 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_717 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_724 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_731 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_738 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_65_745 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_65_752 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_65_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_66_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_457 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_464 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_471 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_478 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_485 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_492 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_499 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_506 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_513 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_520 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_527 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_534 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_541 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_548 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_555 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_562 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_569 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_576 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_583 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_590 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_597 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_604 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_611 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_618 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_625 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_632 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_639 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_646 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_653 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_660 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_667 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_674 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_681 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_688 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_695 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_702 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_709 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_716 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_723 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_730 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_737 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_66_744 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_66_751 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_66_755 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_67_202 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_212 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_219 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_226 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_233 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_240 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_247 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_254 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_261 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_268 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_275 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_282 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_289 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_296 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_303 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_310 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_317 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_324 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_331 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_338 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_345 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_352 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_359 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_366 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_373 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_380 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_387 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_394 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_401 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_408 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_415 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_422 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_429 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_436 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_443 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_450 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_457 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_464 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_471 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_478 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_485 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_492 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_499 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_506 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_513 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_520 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_527 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_534 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_541 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_548 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_555 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_562 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_569 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_576 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_583 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_590 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_597 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_604 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_611 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_618 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_625 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_632 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_639 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_646 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_653 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_660 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_667 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_674 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_681 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_688 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_695 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_702 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_709 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_716 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_723 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_730 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_737 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_67_744 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_67_751 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_67_755 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_202 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_209 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_216 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_223 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_230 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_237 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_244 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_251 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_258 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_265 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_272 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_279 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_286 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_293 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_300 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_307 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_314 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_321 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_328 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_335 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_342 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_349 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_356 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_363 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_370 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_377 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_384 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_391 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_398 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_405 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_412 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_419 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_426 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_433 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_440 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_68_447 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_454 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_461 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_468 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_475 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_482 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_489 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_496 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_503 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_510 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_517 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_524 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_531 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_538 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_545 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_552 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_559 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_566 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_573 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_580 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_587 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_594 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_601 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_608 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_615 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_622 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_629 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_636 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_643 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_650 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_657 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_664 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_671 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_678 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_685 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_692 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_699 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_706 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_713 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_720 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_727 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_734 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_741 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_68_748 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_68_755 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_69_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_69_240 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_247 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_254 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_261 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_268 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_275 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_282 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_289 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_296 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_303 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_310 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_317 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_324 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_331 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_338 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_345 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_352 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_359 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_366 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_373 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_380 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_387 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_394 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_401 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_408 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_415 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_422 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_429 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_436 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_69_456 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_496 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_503 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_510 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_517 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_524 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_531 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_538 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_545 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_552 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_559 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_566 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_573 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_580 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_587 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_594 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_601 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_608 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_615 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_622 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_629 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_636 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_643 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_650 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_657 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_664 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_671 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_678 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_685 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_692 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_699 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_706 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_713 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_720 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_727 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_734 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_741 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_69_748 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_69_755 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_195 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_202 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_70_209 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_70_211 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_221 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_228 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_235 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_242 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_249 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_256 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_263 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_270 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_277 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_284 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_70_291 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_299 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_306 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_313 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_320 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_327 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_334 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_341 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_348 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_355 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_362 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_369 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_376 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_383 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_390 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_397 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_404 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_411 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_418 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_425 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_432 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_439 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_446 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_70_453 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_70_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_70_478 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_70_480 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_484 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_491 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_498 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_505 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_512 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_519 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_526 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_533 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_540 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_547 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_554 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_561 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_568 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_575 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_582 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_589 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_596 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_603 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_610 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_617 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_624 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_631 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_638 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_645 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_652 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_659 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_666 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_673 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_680 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_687 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_694 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_701 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_708 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_715 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_722 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_729 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_736 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_743 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_70_750 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_71_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_71_212 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_71_222 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_228 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_235 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_242 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_249 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_256 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_263 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_270 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_277 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_71_284 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_71_289 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_317 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_324 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_331 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_338 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_345 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_352 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_71_359 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_71_361 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_387 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_71_394 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_71_396 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_422 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_429 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_436 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_443 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_450 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_457 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_464 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_471 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_478 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_485 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_492 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_499 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_506 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_513 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_520 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_527 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_534 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_541 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_548 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_555 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_562 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_569 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_576 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_583 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_590 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_597 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_604 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_611 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_618 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_625 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_632 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_639 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_646 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_653 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_660 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_667 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_674 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_681 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_688 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_695 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_702 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_709 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_716 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_723 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_730 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_737 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_71_744 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_71_751 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_71_755 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_235 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_242 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_249 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_256 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_263 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_270 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_72_277 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_72_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_311 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_318 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_325 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_72_332 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_72_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_367 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_374 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_381 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_388 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_395 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_402 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_409 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_416 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_423 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_72_430 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_72_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_439 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_446 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_453 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_460 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_467 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_474 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_481 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_488 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_495 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_502 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_509 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_516 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_523 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_530 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_537 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_544 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_551 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_558 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_565 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_572 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_579 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_586 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_593 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_600 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_607 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_614 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_621 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_628 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_635 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_642 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_649 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_656 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_663 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_670 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_677 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_684 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_691 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_698 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_705 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_712 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_719 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_726 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_733 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_740 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_72_747 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_72_754 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_72_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_261 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_73_268 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_73_272 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_297 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_304 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_311 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_318 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_325 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_332 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_73_339 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_73_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_73_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_374 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_73_386 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_394 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_401 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_414 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_421 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_428 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_435 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_442 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_73_449 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_73_451 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_457 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_464 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_471 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_478 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_485 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_492 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_499 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_506 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_513 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_520 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_527 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_534 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_541 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_548 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_555 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_562 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_569 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_576 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_583 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_590 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_597 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_604 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_611 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_618 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_625 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_632 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_639 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_646 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_653 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_660 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_667 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_674 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_681 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_688 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_695 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_702 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_709 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_716 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_723 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_730 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_737 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_73_744 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_73_751 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_73_755 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_74_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_74_235 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_74_250 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_74_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_257 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_272 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_279 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_286 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_74_293 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_74_297 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_302 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_309 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_316 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_323 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_330 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_337 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_344 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_74_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_395 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_402 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_409 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_416 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_423 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_430 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_437 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_74_444 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_74_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_74_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_75_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_39 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_46 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_53 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_60 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_67 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_74 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_81 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_88 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_95 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_102 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_109 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_116 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_123 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_130 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_137 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_144 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_151 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_158 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_165 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_172 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_179 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_186 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_193 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_200 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_207 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_214 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_221 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_228 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_75_235 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_75_237 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_243 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_250 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_257 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_264 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_271 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_75_278 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_75_282 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_320 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_327 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_334 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_341 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_348 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_75_355 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_360 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_367 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_374 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_381 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_388 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_395 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_402 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_409 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_416 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_423 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_430 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_437 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_444 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_75_451 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_473 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_480 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_487 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_494 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_501 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_508 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_515 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_522 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_529 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_536 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_543 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_550 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_557 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_564 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_571 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_578 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_585 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_592 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_599 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_606 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_613 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_620 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_627 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_634 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_641 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_648 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_655 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_662 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_669 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_676 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_683 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_690 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_697 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_704 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_711 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_718 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_725 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_732 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_739 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_75_746 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_75_753 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_76_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_76_228 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_243 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_250 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_257 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_264 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_271 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_278 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_285 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_292 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_299 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_306 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_313 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_320 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_327 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_334 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_341 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_348 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_355 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_362 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_369 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_376 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_383 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_390 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_76_397 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_412 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_419 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_426 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_433 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_440 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_447 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_76_454 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_482 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_489 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_496 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_503 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_510 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_517 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_524 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_531 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_538 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_545 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_552 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_559 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_566 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_573 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_580 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_587 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_594 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_601 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_608 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_615 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_622 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_629 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_636 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_643 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_650 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_657 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_664 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_671 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_678 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_685 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_692 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_699 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_706 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_713 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_720 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_727 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_734 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_741 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_76_748 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_76_755 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_77_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_253 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_260 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_267 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_274 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_281 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_288 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_295 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_302 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_309 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_316 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_323 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_330 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_337 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_344 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_351 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_358 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_365 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_372 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_379 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_386 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_77_393 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_421 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_428 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_435 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_442 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_449 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_77_456 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_464 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_471 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_478 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_485 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_492 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_499 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_506 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_513 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_520 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_527 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_534 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_541 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_548 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_555 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_562 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_569 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_576 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_583 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_590 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_597 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_604 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_611 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_618 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_625 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_632 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_639 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_646 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_653 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_660 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_667 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_674 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_681 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_688 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_695 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_702 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_709 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_716 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_723 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_730 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_737 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_77_744 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_4 FILLER_77_751 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_2 FILLER_77_755 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_78_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_78_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_79_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_79_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_80_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_80_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_81_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_81_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_82_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_82_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_83_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_83_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_84_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_84_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_85_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_85_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_86_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_86_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_87_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_87_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_88_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_88_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_89_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_89_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_90_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_90_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_91_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_91_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_92_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_92_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_93_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_93_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_94_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_94_756 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_0 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_7 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_14 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_21 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_28 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_35 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_42 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_49 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_56 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_63 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_70 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_77 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_84 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_91 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_98 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_105 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_112 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_119 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_126 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_133 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_140 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_147 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_154 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_161 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_168 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_175 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_182 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_189 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_196 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_203 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_210 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_217 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_224 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_231 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_238 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_245 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_252 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_259 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_266 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_273 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_280 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_287 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_294 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_301 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_308 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_315 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_322 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_329 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_336 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_343 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_350 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_357 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_364 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_371 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_378 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_385 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_392 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_399 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_406 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_413 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_420 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_427 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_434 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_441 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_448 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_455 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_462 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_469 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_476 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_483 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_490 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_497 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_504 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_511 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_518 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_525 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_532 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_539 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_546 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_553 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_560 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_567 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_574 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_581 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_588 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_595 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_602 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_609 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_616 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_623 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_630 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_637 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_644 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_651 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_658 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_665 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_672 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_679 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_686 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_693 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_700 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_707 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_714 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_721 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_728 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_735 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_742 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_decap_8 FILLER_95_749 (.VDD(VDD),
    .VSS(VSS));
 sg13g2_fill_1 FILLER_95_756 (.VDD(VDD),
    .VSS(VSS));
endmodule
